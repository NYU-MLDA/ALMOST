//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n647_, new_n648_,
    new_n649_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n856_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n884_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G64gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n204_));
  XOR2_X1   g003(.A(G71gat), .B(G78gat), .Z(new_n205_));
  OR2_X1    g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n205_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n206_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT67), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n206_), .B(KEYINPUT12), .C1(new_n207_), .C2(new_n208_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT64), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT6), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(KEYINPUT10), .B(G99gat), .Z(new_n216_));
  INV_X1    g015(.A(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G85gat), .ZN(new_n219_));
  INV_X1    g018(.A(G92gat), .ZN(new_n220_));
  NOR3_X1   g019(.A1(new_n219_), .A2(new_n220_), .A3(KEYINPUT9), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G85gat), .B(G92gat), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n221_), .B1(new_n223_), .B2(KEYINPUT9), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n215_), .A2(new_n218_), .A3(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G99gat), .A2(G106gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT7), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n226_), .B1(KEYINPUT65), .B2(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(KEYINPUT65), .B(KEYINPUT7), .Z(new_n229_));
  AOI21_X1  g028(.A(new_n228_), .B1(new_n229_), .B2(new_n226_), .ZN(new_n230_));
  AOI211_X1 g029(.A(KEYINPUT8), .B(new_n222_), .C1(new_n215_), .C2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT8), .ZN(new_n232_));
  XOR2_X1   g031(.A(KEYINPUT66), .B(KEYINPUT6), .Z(new_n233_));
  OR2_X1    g032(.A1(new_n213_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n213_), .A2(new_n233_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(new_n235_), .A3(new_n230_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n232_), .B1(new_n236_), .B2(new_n223_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n225_), .B1(new_n231_), .B2(new_n237_), .ZN(new_n238_));
  MUX2_X1   g037(.A(new_n210_), .B(new_n211_), .S(new_n238_), .Z(new_n239_));
  NAND2_X1  g038(.A1(G230gat), .A2(G233gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n210_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n242_));
  AOI21_X1  g041(.A(KEYINPUT70), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n241_), .A2(KEYINPUT70), .A3(new_n242_), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n239_), .B(new_n240_), .C1(new_n243_), .C2(new_n244_), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n238_), .A2(new_n210_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n246_), .A2(KEYINPUT68), .A3(new_n241_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n240_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n247_), .B(new_n248_), .C1(KEYINPUT68), .C2(new_n241_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G120gat), .B(G148gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT5), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G176gat), .B(G204gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n251_), .B(new_n252_), .Z(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n245_), .A2(new_n249_), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT71), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT71), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n245_), .A2(new_n249_), .A3(new_n257_), .A4(new_n254_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n245_), .A2(new_n249_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(new_n253_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n259_), .A2(KEYINPUT13), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(KEYINPUT13), .B1(new_n259_), .B2(new_n261_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n202_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n264_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n266_), .A2(KEYINPUT72), .A3(new_n262_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G229gat), .A2(G233gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G29gat), .B(G36gat), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n270_), .A2(KEYINPUT73), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(KEYINPUT73), .ZN(new_n272_));
  XOR2_X1   g071(.A(G43gat), .B(G50gat), .Z(new_n273_));
  OR3_X1    g072(.A1(new_n271_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n273_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G1gat), .B(G8gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G15gat), .B(G22gat), .ZN(new_n278_));
  INV_X1    g077(.A(G1gat), .ZN(new_n279_));
  INV_X1    g078(.A(G8gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT14), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT75), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n278_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n281_), .A2(new_n282_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n277_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  OR3_X1    g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n277_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n276_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT77), .ZN(new_n288_));
  INV_X1    g087(.A(new_n276_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n286_), .A2(new_n285_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n269_), .B1(new_n288_), .B2(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(new_n269_), .B(KEYINPUT78), .Z(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n276_), .B(KEYINPUT15), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n294_), .B1(new_n295_), .B2(new_n290_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n292_), .B1(new_n288_), .B2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G113gat), .B(G141gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G169gat), .B(G197gat), .ZN(new_n299_));
  XOR2_X1   g098(.A(new_n298_), .B(new_n299_), .Z(new_n300_));
  XNOR2_X1  g099(.A(new_n297_), .B(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n268_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  XOR2_X1   g103(.A(G8gat), .B(G36gat), .Z(new_n305_));
  XNOR2_X1  g104(.A(G64gat), .B(G92gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT101), .B(KEYINPUT18), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  NOR3_X1   g108(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n311_), .A2(KEYINPUT24), .ZN(new_n312_));
  INV_X1    g111(.A(G169gat), .ZN(new_n313_));
  INV_X1    g112(.A(G176gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n310_), .B1(new_n312_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G183gat), .A2(G190gat), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT82), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n317_), .A2(new_n318_), .A3(KEYINPUT23), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(KEYINPUT23), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT23), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n321_), .A2(G183gat), .A3(G190gat), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(new_n322_), .A3(KEYINPUT82), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT26), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(G190gat), .ZN(new_n325_));
  INV_X1    g124(.A(G190gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT26), .ZN(new_n327_));
  INV_X1    g126(.A(G183gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT25), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT25), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(G183gat), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n325_), .A2(new_n327_), .A3(new_n329_), .A4(new_n331_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n316_), .A2(new_n319_), .A3(new_n323_), .A4(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n320_), .A2(new_n322_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n328_), .A2(new_n326_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT22), .B(G169gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n314_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n311_), .B(KEYINPUT98), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n336_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT107), .ZN(new_n341_));
  AND3_X1   g140(.A1(new_n333_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n341_), .B1(new_n333_), .B2(new_n340_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(G204gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT92), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT92), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(G204gat), .ZN(new_n348_));
  INV_X1    g147(.A(G197gat), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n346_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT93), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT21), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n352_), .B1(G197gat), .B2(G204gat), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n350_), .A2(new_n351_), .A3(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n351_), .B1(new_n350_), .B2(new_n353_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G211gat), .B(G218gat), .ZN(new_n357_));
  NOR2_X1   g156(.A1(G197gat), .A2(G204gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n346_), .A2(new_n348_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n358_), .B1(new_n359_), .B2(G197gat), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n357_), .B1(new_n360_), .B2(KEYINPUT21), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT94), .B1(new_n356_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n350_), .A2(new_n353_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT93), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n350_), .A2(new_n351_), .A3(new_n353_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT94), .ZN(new_n367_));
  INV_X1    g166(.A(new_n357_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n358_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT92), .B(G204gat), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n369_), .B1(new_n370_), .B2(new_n349_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n368_), .B1(new_n371_), .B2(new_n352_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n366_), .A2(new_n367_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n362_), .A2(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n357_), .A2(new_n352_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n360_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT95), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n360_), .A2(KEYINPUT95), .A3(new_n375_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n344_), .A2(new_n374_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT22), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT80), .B1(new_n382_), .B2(G169gat), .ZN(new_n383_));
  AOI21_X1  g182(.A(G176gat), .B1(new_n382_), .B2(G169gat), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT80), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(new_n313_), .A3(KEYINPUT22), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n383_), .A2(new_n384_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT81), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT81), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n383_), .A2(new_n384_), .A3(new_n386_), .A4(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n323_), .A2(new_n335_), .A3(new_n319_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n392_), .A3(new_n311_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT83), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n329_), .A2(new_n331_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n325_), .A2(KEYINPUT79), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n325_), .A2(new_n327_), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n395_), .B(new_n396_), .C1(new_n397_), .C2(KEYINPUT79), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(new_n316_), .A3(new_n334_), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n393_), .A2(new_n394_), .A3(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n394_), .B1(new_n393_), .B2(new_n399_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  AOI22_X1  g201(.A1(new_n362_), .A2(new_n373_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n381_), .B(KEYINPUT20), .C1(new_n402_), .C2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT108), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G226gat), .A2(G233gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n404_), .A2(new_n405_), .A3(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT20), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n410_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n408_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n333_), .A2(new_n340_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT99), .B1(new_n403_), .B2(new_n414_), .ZN(new_n415_));
  NOR3_X1   g214(.A1(new_n356_), .A2(new_n361_), .A3(KEYINPUT94), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n367_), .B1(new_n366_), .B2(new_n372_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n380_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT99), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n419_), .A3(new_n413_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n411_), .A2(new_n412_), .A3(new_n415_), .A4(new_n420_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n409_), .A2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n405_), .B1(new_n404_), .B2(new_n408_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n309_), .B1(new_n422_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n393_), .A2(new_n399_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT83), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n393_), .A2(new_n394_), .A3(new_n399_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n403_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n415_), .A2(new_n420_), .A3(new_n429_), .A4(KEYINPUT20), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n408_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n427_), .A2(new_n428_), .ZN(new_n432_));
  AOI211_X1 g231(.A(new_n410_), .B(new_n408_), .C1(new_n432_), .C2(new_n418_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT100), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n434_), .B1(new_n418_), .B2(new_n413_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n403_), .A2(KEYINPUT100), .A3(new_n414_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n433_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n431_), .A2(new_n438_), .A3(new_n309_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT27), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT109), .B1(new_n425_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT27), .ZN(new_n442_));
  AOI22_X1  g241(.A1(new_n408_), .A2(new_n430_), .B1(new_n433_), .B2(new_n437_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n442_), .B1(new_n443_), .B2(new_n309_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT109), .ZN(new_n445_));
  INV_X1    g244(.A(new_n309_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n409_), .A2(new_n421_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n446_), .B1(new_n447_), .B2(new_n423_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n444_), .A2(new_n445_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n441_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n431_), .A2(new_n438_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n446_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n439_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n442_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT91), .ZN(new_n455_));
  OAI21_X1  g254(.A(G228gat), .B1(new_n455_), .B2(G233gat), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n456_), .B1(new_n455_), .B2(G233gat), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n457_), .B1(new_n418_), .B2(KEYINPUT90), .ZN(new_n458_));
  NOR2_X1   g257(.A1(G155gat), .A2(G162gat), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT86), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G155gat), .A2(G162gat), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT87), .ZN(new_n463_));
  OR3_X1    g262(.A1(new_n462_), .A2(new_n463_), .A3(KEYINPUT1), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n463_), .B1(new_n462_), .B2(KEYINPUT1), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n461_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  XOR2_X1   g265(.A(G141gat), .B(G148gat), .Z(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n462_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT3), .ZN(new_n470_));
  INV_X1    g269(.A(G141gat), .ZN(new_n471_));
  INV_X1    g270(.A(G148gat), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n470_), .A2(new_n471_), .A3(new_n472_), .A4(KEYINPUT88), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT2), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n474_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT88), .ZN(new_n476_));
  OAI22_X1  g275(.A1(new_n476_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n477_));
  NAND3_X1  g276(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n473_), .A2(new_n475_), .A3(new_n477_), .A4(new_n478_), .ZN(new_n479_));
  AOI22_X1  g278(.A1(new_n479_), .A2(new_n461_), .B1(KEYINPUT1), .B2(new_n467_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n468_), .B1(new_n469_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT29), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n418_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n458_), .A2(new_n483_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n418_), .B(new_n482_), .C1(KEYINPUT90), .C2(new_n457_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G78gat), .B(G106gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n484_), .A2(new_n485_), .A3(new_n487_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G22gat), .B(G50gat), .ZN(new_n492_));
  OR3_X1    g291(.A1(new_n481_), .A2(KEYINPUT29), .A3(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n492_), .B1(new_n481_), .B2(KEYINPUT29), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(KEYINPUT89), .B(KEYINPUT28), .Z(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n487_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n497_), .B1(new_n498_), .B2(KEYINPUT96), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n491_), .A2(new_n499_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n489_), .A2(KEYINPUT96), .A3(new_n490_), .A4(new_n497_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n450_), .A2(new_n454_), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G227gat), .A2(G233gat), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n505_), .B(G15gat), .Z(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT30), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n432_), .B(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT84), .B(G43gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G127gat), .B(G134gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G113gat), .B(G120gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT85), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT85), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n515_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT31), .ZN(new_n518_));
  XOR2_X1   g317(.A(G71gat), .B(G99gat), .Z(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n510_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n510_), .A2(new_n520_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n479_), .A2(new_n461_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n467_), .A2(KEYINPUT1), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  AOI22_X1  g326(.A1(new_n527_), .A2(new_n462_), .B1(new_n467_), .B2(new_n466_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT102), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n528_), .A2(new_n529_), .A3(new_n513_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n528_), .A2(new_n517_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n468_), .B(new_n513_), .C1(new_n469_), .C2(new_n480_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT102), .ZN(new_n533_));
  OAI211_X1 g332(.A(KEYINPUT4), .B(new_n530_), .C1(new_n531_), .C2(new_n533_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n531_), .A2(KEYINPUT4), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G225gat), .A2(G233gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT103), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  OR2_X1    g338(.A1(new_n531_), .A2(new_n533_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n530_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n538_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(G1gat), .B(G29gat), .Z(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT104), .B(KEYINPUT0), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G57gat), .B(G85gat), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n546_), .B(new_n547_), .Z(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n539_), .A2(new_n543_), .A3(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n542_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n538_), .B1(new_n540_), .B2(new_n530_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n548_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n550_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n524_), .A2(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n504_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT110), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n444_), .A2(new_n445_), .A3(new_n448_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n445_), .B1(new_n444_), .B2(new_n448_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n554_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n454_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n558_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n450_), .A2(KEYINPUT110), .A3(new_n454_), .A4(new_n562_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n539_), .A2(new_n543_), .A3(KEYINPUT33), .A4(new_n549_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT105), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT33), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n550_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n536_), .A2(new_n542_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n541_), .A2(new_n538_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n571_), .A2(new_n548_), .A3(new_n572_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n452_), .A2(new_n570_), .A3(new_n439_), .A4(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n309_), .A2(KEYINPUT32), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n575_), .B1(new_n422_), .B2(new_n424_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(KEYINPUT106), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n554_), .B1(new_n451_), .B2(new_n577_), .ZN(new_n578_));
  OAI22_X1  g377(.A1(new_n568_), .A2(new_n574_), .B1(new_n576_), .B2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(new_n503_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n564_), .A2(new_n565_), .A3(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n557_), .B1(new_n581_), .B2(new_n523_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n304_), .A2(new_n582_), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n238_), .A2(new_n289_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n295_), .A2(new_n238_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G232gat), .A2(G233gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT34), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n587_), .A2(KEYINPUT35), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n584_), .A2(new_n585_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(KEYINPUT35), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G190gat), .B(G218gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G134gat), .B(G162gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT36), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n591_), .A2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n594_), .A2(KEYINPUT36), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n591_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(KEYINPUT74), .B(KEYINPUT37), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n290_), .B(new_n602_), .Z(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n604_), .A2(new_n209_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT17), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G127gat), .B(G155gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G183gat), .B(G211gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n605_), .A2(new_n606_), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n604_), .A2(new_n209_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n604_), .A2(new_n210_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n604_), .A2(new_n210_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n611_), .B(KEYINPUT17), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n615_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n614_), .A2(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n601_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n583_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n622_), .A2(new_n279_), .A3(new_n554_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT38), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n599_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n582_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n619_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(new_n303_), .A3(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(G1gat), .B1(new_n629_), .B2(new_n555_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n623_), .A2(new_n624_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n625_), .A2(new_n630_), .A3(new_n631_), .ZN(G1324gat));
  NAND2_X1  g431(.A1(new_n450_), .A2(new_n454_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(G8gat), .B1(new_n629_), .B2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT39), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n622_), .A2(new_n280_), .A3(new_n633_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT40), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(G1325gat));
  OAI21_X1  g439(.A(G15gat), .B1(new_n629_), .B2(new_n523_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(KEYINPUT111), .B(KEYINPUT41), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n642_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n523_), .A2(G15gat), .ZN(new_n645_));
  OAI211_X1 g444(.A(new_n643_), .B(new_n644_), .C1(new_n621_), .C2(new_n645_), .ZN(G1326gat));
  OAI21_X1  g445(.A(G22gat), .B1(new_n629_), .B2(new_n503_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT42), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n503_), .A2(G22gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n648_), .B1(new_n621_), .B2(new_n649_), .ZN(G1327gat));
  NOR2_X1   g449(.A1(new_n599_), .A2(new_n628_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n583_), .A2(new_n651_), .ZN(new_n652_));
  OR3_X1    g451(.A1(new_n652_), .A2(G29gat), .A3(new_n555_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n601_), .ZN(new_n654_));
  OAI21_X1  g453(.A(KEYINPUT43), .B1(new_n582_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT43), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n454_), .B(new_n562_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n657_));
  AOI22_X1  g456(.A1(new_n657_), .A2(new_n558_), .B1(new_n579_), .B2(new_n503_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n524_), .B1(new_n658_), .B2(new_n565_), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n656_), .B(new_n601_), .C1(new_n659_), .C2(new_n557_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n655_), .A2(new_n660_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n265_), .A2(new_n267_), .A3(new_n619_), .A4(new_n301_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT112), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n661_), .A2(KEYINPUT44), .A3(new_n663_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n666_), .A2(new_n667_), .A3(new_n668_), .A4(new_n554_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(G29gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT44), .B1(new_n661_), .B2(new_n663_), .ZN(new_n671_));
  AOI211_X1 g470(.A(new_n665_), .B(new_n662_), .C1(new_n655_), .C2(new_n660_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n667_), .B1(new_n673_), .B2(new_n554_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n653_), .B1(new_n670_), .B2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT113), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT113), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n677_), .B(new_n653_), .C1(new_n670_), .C2(new_n674_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(G1328gat));
  NOR2_X1   g478(.A1(new_n634_), .A2(G36gat), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  OR3_X1    g480(.A1(new_n652_), .A2(KEYINPUT45), .A3(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(KEYINPUT45), .B1(new_n652_), .B2(new_n681_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n671_), .A2(new_n672_), .A3(new_n634_), .ZN(new_n685_));
  INV_X1    g484(.A(G36gat), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n685_), .A2(KEYINPUT114), .A3(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT114), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n666_), .A2(new_n633_), .A3(new_n668_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(G36gat), .ZN(new_n690_));
  OAI211_X1 g489(.A(KEYINPUT46), .B(new_n684_), .C1(new_n687_), .C2(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(KEYINPUT114), .B1(new_n685_), .B2(new_n686_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n689_), .A2(new_n688_), .A3(G36gat), .ZN(new_n693_));
  AOI22_X1  g492(.A1(new_n692_), .A2(new_n693_), .B1(new_n683_), .B2(new_n682_), .ZN(new_n694_));
  XOR2_X1   g493(.A(KEYINPUT115), .B(KEYINPUT46), .Z(new_n695_));
  OAI21_X1  g494(.A(new_n691_), .B1(new_n694_), .B2(new_n695_), .ZN(G1329gat));
  INV_X1    g495(.A(new_n652_), .ZN(new_n697_));
  INV_X1    g496(.A(G43gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n697_), .A2(new_n698_), .A3(new_n524_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n671_), .A2(new_n672_), .A3(new_n523_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n699_), .B1(new_n700_), .B2(new_n698_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g501(.A(G50gat), .B1(new_n697_), .B2(new_n502_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n502_), .A2(G50gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n673_), .B2(new_n704_), .ZN(G1331gat));
  INV_X1    g504(.A(new_n268_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n706_), .A2(new_n301_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n707_), .A2(new_n628_), .A3(new_n627_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT116), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(new_n554_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(G57gat), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n706_), .A2(new_n582_), .A3(new_n301_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n620_), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n555_), .A2(G57gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n711_), .B1(new_n713_), .B2(new_n714_), .ZN(G1332gat));
  INV_X1    g514(.A(new_n713_), .ZN(new_n716_));
  INV_X1    g515(.A(G64gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n716_), .A2(new_n717_), .A3(new_n633_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT48), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n709_), .A2(new_n633_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n720_), .B2(G64gat), .ZN(new_n721_));
  AOI211_X1 g520(.A(KEYINPUT48), .B(new_n717_), .C1(new_n709_), .C2(new_n633_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n718_), .B1(new_n721_), .B2(new_n722_), .ZN(G1333gat));
  INV_X1    g522(.A(G71gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n716_), .A2(new_n724_), .A3(new_n524_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT49), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n709_), .A2(new_n524_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n727_), .B2(G71gat), .ZN(new_n728_));
  AOI211_X1 g527(.A(KEYINPUT49), .B(new_n724_), .C1(new_n709_), .C2(new_n524_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(G1334gat));
  INV_X1    g529(.A(KEYINPUT50), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n709_), .A2(new_n502_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n732_), .B2(G78gat), .ZN(new_n733_));
  INV_X1    g532(.A(G78gat), .ZN(new_n734_));
  AOI211_X1 g533(.A(KEYINPUT50), .B(new_n734_), .C1(new_n709_), .C2(new_n502_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n502_), .A2(new_n734_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT117), .Z(new_n737_));
  OAI22_X1  g536(.A1(new_n733_), .A2(new_n735_), .B1(new_n713_), .B2(new_n737_), .ZN(G1335gat));
  NAND2_X1  g537(.A1(new_n712_), .A2(new_n651_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n740_), .A2(new_n219_), .A3(new_n554_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n661_), .A2(new_n619_), .A3(new_n707_), .ZN(new_n742_));
  OAI21_X1  g541(.A(G85gat), .B1(new_n742_), .B2(new_n555_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1336gat));
  NAND3_X1  g543(.A1(new_n740_), .A2(new_n220_), .A3(new_n633_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G92gat), .B1(new_n742_), .B2(new_n634_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1337gat));
  INV_X1    g546(.A(new_n742_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(new_n524_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n524_), .A2(new_n216_), .ZN(new_n750_));
  AOI22_X1  g549(.A1(new_n749_), .A2(G99gat), .B1(new_n740_), .B2(new_n750_), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g551(.A1(new_n740_), .A2(new_n217_), .A3(new_n502_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n748_), .A2(new_n502_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n755_), .B2(G106gat), .ZN(new_n756_));
  AOI211_X1 g555(.A(KEYINPUT52), .B(new_n217_), .C1(new_n748_), .C2(new_n502_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT53), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT53), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n760_), .B(new_n753_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1339gat));
  NOR2_X1   g561(.A1(new_n263_), .A2(new_n264_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n764_));
  AND4_X1   g563(.A1(new_n620_), .A2(new_n763_), .A3(new_n302_), .A4(new_n764_), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n601_), .A2(new_n619_), .A3(new_n301_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n764_), .B1(new_n766_), .B2(new_n763_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n765_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n245_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT119), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n245_), .A2(new_n769_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT119), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n245_), .A2(new_n773_), .A3(new_n769_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n239_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n248_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n771_), .A2(new_n772_), .A3(new_n774_), .A4(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n253_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT56), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT120), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n777_), .A2(KEYINPUT120), .A3(new_n779_), .A4(new_n253_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n259_), .A2(new_n301_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n781_), .A2(new_n782_), .A3(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n259_), .A2(new_n261_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n288_), .A2(new_n291_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n293_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n293_), .B1(new_n295_), .B2(new_n290_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n300_), .B1(new_n789_), .B2(new_n288_), .ZN(new_n790_));
  AOI22_X1  g589(.A1(new_n297_), .A2(new_n300_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n786_), .A2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n626_), .B1(new_n785_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n778_), .A2(KEYINPUT56), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT58), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT121), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n777_), .A2(new_n779_), .A3(new_n253_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n259_), .A2(new_n791_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n794_), .A2(new_n796_), .A3(new_n797_), .A4(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n601_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n798_), .B1(new_n778_), .B2(KEYINPUT56), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n796_), .B1(new_n802_), .B2(new_n797_), .ZN(new_n803_));
  OAI22_X1  g602(.A1(new_n793_), .A2(KEYINPUT57), .B1(new_n801_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT122), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n803_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n807_), .A2(new_n601_), .A3(new_n800_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT57), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n783_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n810_));
  AOI22_X1  g609(.A1(new_n810_), .A2(new_n782_), .B1(new_n786_), .B2(new_n791_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n809_), .B1(new_n811_), .B2(new_n626_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n808_), .A2(new_n812_), .A3(KEYINPUT122), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n793_), .A2(KEYINPUT57), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n806_), .A2(new_n813_), .A3(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n768_), .B1(new_n815_), .B2(new_n619_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n504_), .A2(new_n555_), .A3(new_n523_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT59), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(KEYINPUT123), .B1(new_n816_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT123), .ZN(new_n821_));
  INV_X1    g620(.A(new_n819_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n811_), .A2(new_n809_), .A3(new_n626_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n823_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n628_), .B1(new_n824_), .B2(new_n813_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n821_), .B(new_n822_), .C1(new_n825_), .C2(new_n768_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n619_), .B1(new_n804_), .B2(new_n823_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n765_), .B2(new_n767_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n817_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT59), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n820_), .A2(new_n301_), .A3(new_n826_), .A4(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(G113gat), .ZN(new_n832_));
  OR3_X1    g631(.A1(new_n829_), .A2(G113gat), .A3(new_n302_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(G1340gat));
  NAND4_X1  g633(.A1(new_n820_), .A2(new_n268_), .A3(new_n826_), .A4(new_n830_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(G120gat), .ZN(new_n836_));
  INV_X1    g635(.A(new_n829_), .ZN(new_n837_));
  INV_X1    g636(.A(G120gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n706_), .B2(KEYINPUT60), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n837_), .B(new_n839_), .C1(KEYINPUT60), .C2(new_n838_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n836_), .A2(new_n840_), .ZN(G1341gat));
  NAND4_X1  g640(.A1(new_n820_), .A2(new_n628_), .A3(new_n826_), .A4(new_n830_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(G127gat), .ZN(new_n843_));
  OR3_X1    g642(.A1(new_n829_), .A2(G127gat), .A3(new_n619_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(G1342gat));
  NAND4_X1  g644(.A1(new_n820_), .A2(new_n601_), .A3(new_n826_), .A4(new_n830_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(G134gat), .ZN(new_n847_));
  OR3_X1    g646(.A1(new_n829_), .A2(G134gat), .A3(new_n599_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1343gat));
  NAND3_X1  g648(.A1(new_n808_), .A2(new_n814_), .A3(new_n812_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n768_), .B1(new_n850_), .B2(new_n619_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n523_), .A2(new_n502_), .A3(new_n554_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n851_), .A2(new_n633_), .A3(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n301_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g654(.A1(new_n853_), .A2(new_n268_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g656(.A1(new_n853_), .A2(new_n628_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(KEYINPUT61), .B(G155gat), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1346gat));
  AOI21_X1  g659(.A(G162gat), .B1(new_n853_), .B2(new_n626_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n601_), .A2(G162gat), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT124), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n861_), .B1(new_n853_), .B2(new_n863_), .ZN(G1347gat));
  NOR3_X1   g663(.A1(new_n634_), .A2(new_n502_), .A3(new_n556_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n301_), .B(new_n865_), .C1(new_n825_), .C2(new_n768_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(G169gat), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT62), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n866_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n870_));
  INV_X1    g669(.A(new_n337_), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n869_), .B(new_n870_), .C1(new_n871_), .C2(new_n866_), .ZN(G1348gat));
  INV_X1    g671(.A(new_n816_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n873_), .A2(new_n865_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n268_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n828_), .A2(new_n865_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n706_), .A2(new_n314_), .ZN(new_n877_));
  AOI22_X1  g676(.A1(new_n875_), .A2(new_n314_), .B1(new_n876_), .B2(new_n877_), .ZN(G1349gat));
  AOI21_X1  g677(.A(G183gat), .B1(new_n876_), .B2(new_n628_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n619_), .A2(new_n395_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n874_), .B2(new_n880_), .ZN(G1350gat));
  NAND3_X1  g680(.A1(new_n874_), .A2(new_n626_), .A3(new_n397_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n873_), .A2(new_n865_), .ZN(new_n883_));
  OAI21_X1  g682(.A(G190gat), .B1(new_n883_), .B2(new_n654_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n882_), .A2(new_n884_), .ZN(G1351gat));
  INV_X1    g684(.A(KEYINPUT125), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n633_), .A2(new_n523_), .A3(new_n562_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n828_), .A2(new_n886_), .A3(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(KEYINPUT125), .B1(new_n851_), .B2(new_n887_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n301_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g692(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n894_));
  AND4_X1   g693(.A1(new_n359_), .A2(new_n891_), .A3(new_n268_), .A4(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n345_), .A2(KEYINPUT126), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n896_), .B1(new_n891_), .B2(new_n268_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n895_), .A2(new_n897_), .ZN(G1353gat));
  OR2_X1    g697(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n899_));
  NAND2_X1  g698(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n900_));
  AND4_X1   g699(.A1(new_n628_), .A2(new_n891_), .A3(new_n899_), .A4(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n899_), .B1(new_n891_), .B2(new_n628_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1354gat));
  AND3_X1   g702(.A1(new_n891_), .A2(G218gat), .A3(new_n601_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n599_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT127), .ZN(new_n906_));
  AOI21_X1  g705(.A(G218gat), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n891_), .A2(new_n626_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(KEYINPUT127), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n904_), .B1(new_n907_), .B2(new_n909_), .ZN(G1355gat));
endmodule


