//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 0 0 0 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n808_, new_n809_, new_n811_,
    new_n812_, new_n814_, new_n815_, new_n816_, new_n817_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G50gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT74), .B(G43gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT15), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT66), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n207_), .B1(new_n208_), .B2(KEYINPUT67), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT7), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT6), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT7), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n213_), .B1(new_n208_), .B2(new_n207_), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n210_), .B(new_n212_), .C1(new_n209_), .C2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT68), .ZN(new_n216_));
  XOR2_X1   g015(.A(G85gat), .B(G92gat), .Z(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT8), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(G85gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n222_), .A2(KEYINPUT9), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n221_), .A2(G85gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(G92gat), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(KEYINPUT10), .B(G99gat), .Z(new_n226_));
  INV_X1    g025(.A(G106gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n217_), .A2(KEYINPUT9), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n225_), .A2(new_n228_), .A3(new_n229_), .A4(new_n212_), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n215_), .A2(new_n216_), .A3(KEYINPUT8), .A4(new_n217_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n220_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n206_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n205_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G232gat), .A2(G233gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT34), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT35), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n233_), .A2(new_n235_), .A3(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n238_), .A2(new_n239_), .ZN(new_n242_));
  OR2_X1    g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT76), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n241_), .A2(new_n242_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(G134gat), .B(G162gat), .Z(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(G218gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT75), .B(G190gat), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n248_), .B(new_n249_), .Z(new_n250_));
  NOR2_X1   g049(.A1(new_n250_), .A2(KEYINPUT36), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n246_), .A2(new_n252_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .A4(new_n251_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT37), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n243_), .A2(new_n245_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(KEYINPUT36), .A3(new_n250_), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n255_), .A2(new_n256_), .A3(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n256_), .B1(new_n255_), .B2(new_n258_), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT69), .B(G71gat), .ZN(new_n262_));
  INV_X1    g061(.A(G78gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT11), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n262_), .B(G78gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT11), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT70), .B(G57gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(G64gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n271_), .B1(KEYINPUT11), .B2(new_n264_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G15gat), .B(G22gat), .ZN(new_n276_));
  INV_X1    g075(.A(G1gat), .ZN(new_n277_));
  INV_X1    g076(.A(G8gat), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT14), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n276_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G1gat), .B(G8gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G231gat), .A2(G233gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT77), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n282_), .B(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n275_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G127gat), .B(G155gat), .ZN(new_n287_));
  INV_X1    g086(.A(G211gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT16), .B(G183gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT17), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n286_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT78), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n291_), .A2(new_n292_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n286_), .A2(new_n294_), .A3(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n261_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT13), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G120gat), .B(G148gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(G204gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT5), .B(G176gat), .ZN(new_n304_));
  XOR2_X1   g103(.A(new_n303_), .B(new_n304_), .Z(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT71), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n307_), .A2(KEYINPUT12), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n308_), .B1(new_n275_), .B2(new_n232_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n275_), .A2(new_n232_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n273_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n311_), .A2(new_n230_), .A3(new_n220_), .A4(new_n231_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n307_), .A2(KEYINPUT12), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n310_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n309_), .B1(new_n314_), .B2(new_n308_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G230gat), .A2(G233gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT64), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n315_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT72), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n315_), .A2(KEYINPUT72), .A3(new_n318_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n318_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n306_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  AOI211_X1 g125(.A(new_n324_), .B(new_n305_), .C1(new_n321_), .C2(new_n322_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n301_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n322_), .ZN(new_n329_));
  AOI21_X1  g128(.A(KEYINPUT72), .B1(new_n315_), .B2(new_n318_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n325_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(new_n305_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n323_), .A2(new_n325_), .A3(new_n306_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(KEYINPUT13), .A3(new_n333_), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n328_), .A2(new_n334_), .A3(KEYINPUT73), .ZN(new_n335_));
  AOI21_X1  g134(.A(KEYINPUT73), .B1(new_n328_), .B2(new_n334_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n300_), .A2(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n338_), .B(KEYINPUT79), .Z(new_n339_));
  INV_X1    g138(.A(KEYINPUT80), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n234_), .A2(new_n282_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n341_), .B1(new_n206_), .B2(new_n282_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G229gat), .A2(G233gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n205_), .B(new_n282_), .Z(new_n345_));
  INV_X1    g144(.A(new_n343_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n340_), .B1(new_n344_), .B2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n348_), .B1(new_n340_), .B2(new_n347_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G113gat), .B(G141gat), .ZN(new_n350_));
  INV_X1    g149(.A(G197gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT81), .B(G169gat), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n352_), .B(new_n353_), .Z(new_n354_));
  XNOR2_X1  g153(.A(new_n349_), .B(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT86), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G155gat), .A2(G162gat), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n357_), .B1(new_n358_), .B2(KEYINPUT1), .ZN(new_n359_));
  OR2_X1    g158(.A1(G155gat), .A2(G162gat), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT1), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n361_), .A2(KEYINPUT86), .A3(G155gat), .A4(G162gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n358_), .A2(KEYINPUT1), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n359_), .A2(new_n360_), .A3(new_n362_), .A4(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G141gat), .A2(G148gat), .ZN(new_n365_));
  OR2_X1    g164(.A1(G141gat), .A2(G148gat), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n364_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT87), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n366_), .A2(KEYINPUT3), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT2), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n365_), .A2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n366_), .A2(KEYINPUT3), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n370_), .A2(new_n372_), .A3(new_n373_), .A4(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(new_n360_), .A3(new_n358_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n369_), .A2(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G127gat), .B(G134gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G113gat), .B(G120gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT97), .B(KEYINPUT4), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n377_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  OR2_X1    g182(.A1(new_n383_), .A2(KEYINPUT98), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n369_), .A2(new_n376_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n380_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n377_), .A2(new_n381_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(KEYINPUT4), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G225gat), .A2(G233gat), .ZN(new_n389_));
  XOR2_X1   g188(.A(new_n389_), .B(KEYINPUT96), .Z(new_n390_));
  NAND2_X1  g189(.A1(new_n383_), .A2(KEYINPUT98), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n384_), .A2(new_n388_), .A3(new_n390_), .A4(new_n391_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n386_), .A2(new_n387_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n390_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n392_), .A2(new_n395_), .ZN(new_n396_));
  XOR2_X1   g195(.A(G1gat), .B(G29gat), .Z(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(G85gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT0), .B(G57gat), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n398_), .B(new_n399_), .Z(new_n400_));
  NAND2_X1  g199(.A1(new_n396_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n400_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n392_), .A2(new_n395_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT90), .ZN(new_n405_));
  INV_X1    g204(.A(G204gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(KEYINPUT90), .A2(G204gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n351_), .A3(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT91), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  OR2_X1    g210(.A1(KEYINPUT89), .A2(G197gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(KEYINPUT89), .A2(G197gat), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n412_), .A2(new_n406_), .A3(new_n413_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n407_), .A2(KEYINPUT91), .A3(new_n351_), .A4(new_n408_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n411_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT21), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT92), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  XOR2_X1   g218(.A(G211gat), .B(G218gat), .Z(new_n420_));
  AOI21_X1  g219(.A(new_n406_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n407_), .A2(new_n408_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n421_), .B1(G197gat), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT21), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n420_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n416_), .A2(KEYINPUT92), .A3(KEYINPUT21), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n419_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n420_), .ZN(new_n428_));
  OR3_X1    g227(.A1(new_n423_), .A2(new_n424_), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G183gat), .A2(G190gat), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT23), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(KEYINPUT84), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT84), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n435_), .A2(G183gat), .A3(G190gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n433_), .B1(new_n437_), .B2(new_n432_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G169gat), .A2(G176gat), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n438_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n442_));
  NOR3_X1   g241(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT25), .B(G183gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT26), .B(G190gat), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n443_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n431_), .A2(new_n432_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n447_), .B1(new_n437_), .B2(new_n432_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n448_), .B1(G183gat), .B2(G190gat), .ZN(new_n449_));
  XOR2_X1   g248(.A(new_n439_), .B(KEYINPUT83), .Z(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT22), .B(G169gat), .ZN(new_n451_));
  INV_X1    g250(.A(G176gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n450_), .A2(new_n453_), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n442_), .A2(new_n446_), .B1(new_n449_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n430_), .A2(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(G183gat), .A2(G190gat), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n454_), .B1(new_n438_), .B2(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n443_), .B1(new_n450_), .B2(new_n441_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT82), .ZN(new_n461_));
  INV_X1    g260(.A(G190gat), .ZN(new_n462_));
  OR3_X1    g261(.A1(new_n461_), .A2(new_n462_), .A3(KEYINPUT26), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT26), .B1(new_n461_), .B2(new_n462_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n463_), .A2(new_n464_), .A3(new_n444_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n460_), .A2(new_n448_), .A3(new_n465_), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n459_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n467_), .A2(new_n427_), .A3(new_n429_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n457_), .A2(KEYINPUT20), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G226gat), .A2(G233gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT19), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT95), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n427_), .A2(new_n429_), .A3(new_n455_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n474_), .A2(KEYINPUT20), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n459_), .A2(new_n466_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n471_), .B1(new_n430_), .B2(new_n476_), .ZN(new_n477_));
  AOI22_X1  g276(.A1(new_n469_), .A2(new_n473_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G8gat), .B(G36gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(G92gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT18), .B(G64gat), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n480_), .B(new_n481_), .Z(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT32), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n478_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT100), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n474_), .A2(KEYINPUT20), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT99), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n467_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n474_), .A2(KEYINPUT99), .A3(KEYINPUT20), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n488_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(new_n471_), .ZN(new_n493_));
  AND4_X1   g292(.A1(KEYINPUT20), .A2(new_n457_), .A3(new_n472_), .A4(new_n468_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n483_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n485_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n494_), .B1(new_n492_), .B2(new_n471_), .ZN(new_n499_));
  NOR3_X1   g298(.A1(new_n499_), .A2(KEYINPUT100), .A3(new_n483_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n404_), .B(new_n484_), .C1(new_n498_), .C2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT101), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n478_), .A2(new_n482_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n384_), .A2(new_n388_), .A3(new_n394_), .A4(new_n391_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n393_), .A2(new_n390_), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n506_), .A2(new_n400_), .A3(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n478_), .A2(new_n482_), .ZN(new_n509_));
  NOR3_X1   g308(.A1(new_n505_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n403_), .B(KEYINPUT33), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT88), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT29), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n512_), .B1(new_n385_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G228gat), .A2(G233gat), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n377_), .A2(KEYINPUT88), .A3(KEYINPUT29), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n514_), .A2(new_n515_), .A3(new_n430_), .A4(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n430_), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n513_), .A2(KEYINPUT93), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n513_), .A2(KEYINPUT93), .ZN(new_n520_));
  AOI211_X1 g319(.A(new_n519_), .B(new_n520_), .C1(new_n369_), .C2(new_n376_), .ZN(new_n521_));
  OAI211_X1 g320(.A(G228gat), .B(G233gat), .C1(new_n518_), .C2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n517_), .A2(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(G78gat), .B(G106gat), .Z(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n517_), .A2(new_n522_), .A3(new_n524_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n377_), .A2(KEYINPUT29), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT28), .B(G22gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(G50gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n528_), .B(new_n530_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n526_), .B(new_n527_), .C1(KEYINPUT94), .C2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n526_), .A2(new_n527_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n531_), .B1(new_n527_), .B2(KEYINPUT94), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  AOI22_X1  g334(.A1(new_n510_), .A2(new_n511_), .B1(new_n532_), .B2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n496_), .A2(new_n485_), .A3(new_n497_), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT100), .B1(new_n499_), .B2(new_n483_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n539_), .A2(KEYINPUT101), .A3(new_n404_), .A4(new_n484_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n503_), .A2(new_n536_), .A3(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(KEYINPUT85), .B(KEYINPUT31), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT30), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n476_), .B(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G15gat), .B(G43gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G227gat), .A2(G233gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n544_), .B(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G71gat), .B(G99gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n380_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n548_), .B(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n404_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT27), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n553_), .B1(new_n505_), .B2(new_n509_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n482_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n471_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n489_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n556_), .B1(new_n557_), .B2(new_n491_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n555_), .B1(new_n558_), .B2(new_n494_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT102), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n553_), .B1(new_n478_), .B2(new_n482_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n559_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n560_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n552_), .B(new_n554_), .C1(new_n562_), .C2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n535_), .A2(new_n532_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n551_), .B1(new_n564_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n541_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT103), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n565_), .A2(new_n551_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n569_), .B1(new_n564_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n509_), .ZN(new_n572_));
  AOI21_X1  g371(.A(KEYINPUT27), .B1(new_n572_), .B2(new_n504_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n482_), .B1(new_n493_), .B2(new_n495_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n504_), .A2(KEYINPUT27), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT102), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n559_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n573_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n551_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n579_), .B1(new_n535_), .B2(new_n532_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n578_), .A2(KEYINPUT103), .A3(new_n580_), .A4(new_n552_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n571_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n568_), .A2(new_n582_), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n339_), .A2(new_n356_), .A3(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n584_), .A2(new_n277_), .A3(new_n404_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT38), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n335_), .A2(new_n336_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n587_), .A2(new_n355_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n588_), .A2(new_n583_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n255_), .A2(new_n258_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n590_), .A2(new_n299_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(G1gat), .B1(new_n592_), .B2(new_n552_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n586_), .A2(new_n593_), .ZN(G1324gat));
  OAI21_X1  g393(.A(G8gat), .B1(new_n592_), .B2(new_n578_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT104), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  OAI211_X1 g396(.A(KEYINPUT104), .B(G8gat), .C1(new_n592_), .C2(new_n578_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n597_), .A2(KEYINPUT39), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n578_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n584_), .A2(new_n278_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT39), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n595_), .A2(new_n596_), .A3(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n599_), .A2(new_n601_), .A3(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n599_), .A2(new_n601_), .A3(new_n603_), .A4(new_n605_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(G1325gat));
  OAI21_X1  g408(.A(G15gat), .B1(new_n592_), .B2(new_n579_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT41), .Z(new_n611_));
  INV_X1    g410(.A(G15gat), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n584_), .A2(new_n612_), .A3(new_n551_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(G1326gat));
  XNOR2_X1  g413(.A(new_n565_), .B(KEYINPUT106), .ZN(new_n615_));
  OAI21_X1  g414(.A(G22gat), .B1(new_n592_), .B2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT42), .ZN(new_n617_));
  INV_X1    g416(.A(G22gat), .ZN(new_n618_));
  INV_X1    g417(.A(new_n615_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n584_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(new_n620_), .ZN(G1327gat));
  INV_X1    g420(.A(new_n590_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n299_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n589_), .A2(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(G29gat), .B1(new_n625_), .B2(new_n404_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n583_), .A2(new_n261_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT43), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT43), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n583_), .A2(new_n629_), .A3(new_n261_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n631_), .A2(new_n588_), .A3(new_n299_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT44), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n634_), .A2(G29gat), .A3(new_n404_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n632_), .A2(new_n633_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n626_), .B1(new_n635_), .B2(new_n636_), .ZN(G1328gat));
  INV_X1    g436(.A(G36gat), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n625_), .A2(new_n638_), .A3(new_n600_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT45), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n636_), .A2(new_n600_), .A3(new_n634_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(G36gat), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT46), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n640_), .A2(KEYINPUT46), .A3(new_n642_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(G1329gat));
  NAND4_X1  g446(.A1(new_n636_), .A2(G43gat), .A3(new_n551_), .A4(new_n634_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n625_), .A2(new_n551_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n648_), .B1(G43gat), .B2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g450(.A(G50gat), .B1(new_n625_), .B2(new_n619_), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n636_), .A2(G50gat), .A3(new_n634_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n652_), .B1(new_n653_), .B2(new_n566_), .ZN(G1331gat));
  AND4_X1   g453(.A1(new_n355_), .A2(new_n587_), .A3(new_n583_), .A4(new_n591_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(KEYINPUT108), .B(G57gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(new_n404_), .A3(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT109), .ZN(new_n658_));
  INV_X1    g457(.A(G57gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n356_), .B1(new_n568_), .B2(new_n582_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT107), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n661_), .A2(new_n587_), .A3(new_n300_), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n662_), .A2(new_n552_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n658_), .B1(new_n659_), .B2(new_n663_), .ZN(G1332gat));
  INV_X1    g463(.A(G64gat), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n665_), .B1(new_n655_), .B2(new_n600_), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n666_), .B(KEYINPUT48), .Z(new_n667_));
  NAND2_X1  g466(.A1(new_n600_), .A2(new_n665_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n667_), .B1(new_n662_), .B2(new_n668_), .ZN(G1333gat));
  INV_X1    g468(.A(G71gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n670_), .B1(new_n655_), .B2(new_n551_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT49), .Z(new_n672_));
  NAND2_X1  g471(.A1(new_n551_), .A2(new_n670_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n672_), .B1(new_n662_), .B2(new_n673_), .ZN(G1334gat));
  AOI21_X1  g473(.A(new_n263_), .B1(new_n655_), .B2(new_n619_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT50), .Z(new_n676_));
  NAND2_X1  g475(.A1(new_n619_), .A2(new_n263_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n676_), .B1(new_n662_), .B2(new_n677_), .ZN(G1335gat));
  NAND3_X1  g477(.A1(new_n661_), .A2(new_n587_), .A3(new_n624_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT110), .ZN(new_n680_));
  AOI21_X1  g479(.A(G85gat), .B1(new_n680_), .B2(new_n404_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n631_), .A2(KEYINPUT111), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n355_), .B(new_n299_), .C1(new_n335_), .C2(new_n336_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT111), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n628_), .A2(new_n685_), .A3(new_n630_), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n682_), .A2(new_n684_), .A3(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n224_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n552_), .B1(new_n688_), .B2(new_n222_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n681_), .B1(new_n687_), .B2(new_n689_), .ZN(G1336gat));
  AND3_X1   g489(.A1(new_n687_), .A2(G92gat), .A3(new_n600_), .ZN(new_n691_));
  AOI21_X1  g490(.A(G92gat), .B1(new_n680_), .B2(new_n600_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT112), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n693_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n691_), .B1(new_n694_), .B2(new_n695_), .ZN(G1337gat));
  NAND4_X1  g495(.A1(new_n682_), .A2(new_n551_), .A3(new_n684_), .A4(new_n686_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT113), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n697_), .A2(new_n698_), .A3(G99gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n697_), .B2(G99gat), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT110), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n679_), .B(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n551_), .A2(new_n226_), .ZN(new_n703_));
  OAI22_X1  g502(.A1(new_n699_), .A2(new_n700_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g504(.A1(new_n680_), .A2(new_n227_), .A3(new_n566_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n683_), .A2(new_n565_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n629_), .B1(new_n583_), .B2(new_n261_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n259_), .A2(new_n260_), .ZN(new_n709_));
  AOI211_X1 g508(.A(KEYINPUT43), .B(new_n709_), .C1(new_n568_), .C2(new_n582_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n707_), .B1(new_n708_), .B2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT114), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT114), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n713_), .B(new_n707_), .C1(new_n708_), .C2(new_n710_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n712_), .A2(G106gat), .A3(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT115), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT52), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT115), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n712_), .A2(new_n718_), .A3(G106gat), .A4(new_n714_), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n716_), .A2(new_n717_), .A3(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n717_), .B1(new_n716_), .B2(new_n719_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n706_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n723_), .B(new_n706_), .C1(new_n720_), .C2(new_n721_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1339gat));
  INV_X1    g526(.A(G113gat), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n328_), .A2(new_n334_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n300_), .A2(new_n355_), .A3(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n731_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n300_), .A2(new_n355_), .A3(new_n729_), .A4(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n354_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n345_), .A2(new_n343_), .ZN(new_n738_));
  AOI211_X1 g537(.A(new_n737_), .B(new_n738_), .C1(new_n346_), .C2(new_n342_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n349_), .B2(new_n737_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n315_), .A2(KEYINPUT55), .A3(new_n318_), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n315_), .A2(new_n318_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n329_), .A2(new_n330_), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n741_), .B(new_n742_), .C1(new_n743_), .C2(KEYINPUT55), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n744_), .A2(KEYINPUT56), .A3(new_n305_), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT56), .B1(new_n744_), .B2(new_n305_), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n333_), .B(new_n740_), .C1(new_n745_), .C2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT58), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n744_), .A2(new_n305_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT56), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n744_), .A2(KEYINPUT56), .A3(new_n305_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n754_), .A2(KEYINPUT58), .A3(new_n333_), .A4(new_n740_), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n749_), .A2(new_n755_), .A3(new_n261_), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n356_), .B(new_n333_), .C1(new_n745_), .C2(new_n746_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n740_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(KEYINPUT57), .B1(new_n759_), .B2(new_n622_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT57), .ZN(new_n761_));
  AOI211_X1 g560(.A(new_n761_), .B(new_n590_), .C1(new_n757_), .C2(new_n758_), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n756_), .A2(new_n760_), .A3(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n736_), .B1(new_n763_), .B2(new_n623_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n764_), .A2(new_n404_), .A3(new_n578_), .A4(new_n580_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n728_), .B1(new_n765_), .B2(new_n355_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT118), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT118), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n768_), .B(new_n728_), .C1(new_n765_), .C2(new_n355_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT59), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n765_), .A2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n759_), .A2(new_n622_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n761_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n749_), .A2(new_n755_), .A3(new_n261_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n759_), .A2(KEYINPUT57), .A3(new_n622_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n774_), .A2(new_n775_), .A3(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n299_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n600_), .B1(new_n778_), .B2(new_n736_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n779_), .A2(KEYINPUT59), .A3(new_n404_), .A4(new_n580_), .ZN(new_n780_));
  AOI211_X1 g579(.A(new_n728_), .B(new_n355_), .C1(new_n772_), .C2(new_n780_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n770_), .A2(new_n781_), .ZN(G1340gat));
  INV_X1    g581(.A(new_n765_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT60), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n784_), .B1(new_n337_), .B2(G120gat), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n783_), .B(new_n785_), .C1(new_n784_), .C2(G120gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n337_), .B1(new_n772_), .B2(new_n780_), .ZN(new_n787_));
  INV_X1    g586(.A(G120gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n786_), .B1(new_n787_), .B2(new_n788_), .ZN(G1341gat));
  INV_X1    g588(.A(G127gat), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n790_), .B1(new_n765_), .B2(new_n299_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT119), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  OAI211_X1 g592(.A(KEYINPUT119), .B(new_n790_), .C1(new_n765_), .C2(new_n299_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  AOI211_X1 g594(.A(new_n790_), .B(new_n299_), .C1(new_n772_), .C2(new_n780_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n795_), .A2(new_n796_), .ZN(G1342gat));
  AOI21_X1  g596(.A(G134gat), .B1(new_n783_), .B2(new_n590_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n709_), .B1(new_n772_), .B2(new_n780_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(G134gat), .ZN(G1343gat));
  AOI21_X1  g599(.A(new_n735_), .B1(new_n777_), .B2(new_n299_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n801_), .A2(new_n552_), .A3(new_n600_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n565_), .A2(new_n551_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n804_), .A2(new_n355_), .ZN(new_n805_));
  INV_X1    g604(.A(G141gat), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n805_), .B(new_n806_), .ZN(G1344gat));
  NOR2_X1   g606(.A1(new_n804_), .A2(new_n337_), .ZN(new_n808_));
  XOR2_X1   g607(.A(KEYINPUT120), .B(G148gat), .Z(new_n809_));
  XNOR2_X1  g608(.A(new_n808_), .B(new_n809_), .ZN(G1345gat));
  NOR2_X1   g609(.A1(new_n804_), .A2(new_n299_), .ZN(new_n811_));
  XOR2_X1   g610(.A(KEYINPUT61), .B(G155gat), .Z(new_n812_));
  XNOR2_X1  g611(.A(new_n811_), .B(new_n812_), .ZN(G1346gat));
  INV_X1    g612(.A(G162gat), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n804_), .A2(new_n814_), .A3(new_n709_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n804_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n590_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n815_), .B1(new_n814_), .B2(new_n817_), .ZN(G1347gat));
  NOR2_X1   g617(.A1(new_n578_), .A2(new_n404_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n551_), .ZN(new_n820_));
  XOR2_X1   g619(.A(new_n820_), .B(KEYINPUT121), .Z(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n801_), .A2(new_n619_), .A3(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n823_), .A2(new_n356_), .A3(new_n451_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n801_), .A2(new_n619_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n821_), .A2(new_n356_), .ZN(new_n826_));
  XOR2_X1   g625(.A(new_n826_), .B(KEYINPUT122), .Z(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(G169gat), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n829_), .A2(KEYINPUT62), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n829_), .A2(KEYINPUT62), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n824_), .B1(new_n830_), .B2(new_n831_), .ZN(G1348gat));
  AOI21_X1  g631(.A(G176gat), .B1(new_n823_), .B2(new_n587_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n801_), .A2(new_n566_), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n822_), .A2(new_n452_), .A3(new_n337_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n833_), .B1(new_n834_), .B2(new_n835_), .ZN(G1349gat));
  INV_X1    g635(.A(new_n823_), .ZN(new_n837_));
  OR2_X1    g636(.A1(new_n299_), .A2(new_n444_), .ZN(new_n838_));
  NOR4_X1   g637(.A1(new_n801_), .A2(new_n566_), .A3(new_n299_), .A4(new_n822_), .ZN(new_n839_));
  OAI22_X1  g638(.A1(new_n837_), .A2(new_n838_), .B1(new_n839_), .B2(G183gat), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT123), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n840_), .B(new_n841_), .ZN(G1350gat));
  INV_X1    g641(.A(KEYINPUT124), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n823_), .A2(new_n261_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(G190gat), .ZN(new_n845_));
  AOI211_X1 g644(.A(KEYINPUT124), .B(new_n462_), .C1(new_n823_), .C2(new_n261_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n590_), .A2(new_n445_), .ZN(new_n847_));
  XOR2_X1   g646(.A(new_n847_), .B(KEYINPUT125), .Z(new_n848_));
  OAI22_X1  g647(.A1(new_n845_), .A2(new_n846_), .B1(new_n837_), .B2(new_n848_), .ZN(G1351gat));
  NAND2_X1  g648(.A1(new_n819_), .A2(new_n803_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n764_), .A2(KEYINPUT126), .A3(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT126), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(new_n801_), .B2(new_n850_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n356_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(G197gat), .ZN(G1352gat));
  AOI21_X1  g656(.A(new_n337_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n422_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n406_), .B2(new_n858_), .ZN(G1353gat));
  AOI21_X1  g659(.A(KEYINPUT126), .B1(new_n764_), .B2(new_n851_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n801_), .A2(new_n853_), .A3(new_n850_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n623_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT127), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT63), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n863_), .A2(new_n864_), .A3(new_n865_), .A4(new_n288_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n299_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n288_), .ZN(new_n868_));
  OAI21_X1  g667(.A(KEYINPUT127), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  XOR2_X1   g668(.A(KEYINPUT63), .B(G211gat), .Z(new_n870_));
  AOI22_X1  g669(.A1(new_n866_), .A2(new_n869_), .B1(new_n867_), .B2(new_n870_), .ZN(G1354gat));
  AOI21_X1  g670(.A(G218gat), .B1(new_n855_), .B2(new_n590_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n709_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n872_), .B1(G218gat), .B2(new_n873_), .ZN(G1355gat));
endmodule


