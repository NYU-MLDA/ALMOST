//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 0 0 0 0 0 1 0 1 1 1 1 1 1 0 0 0 0 0 1 1 0 0 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 1 0 0 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n635_,
    new_n636_, new_n637_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n706_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n866_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_;
  XNOR2_X1  g000(.A(KEYINPUT18), .B(G64gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G92gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G8gat), .B(G36gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  XOR2_X1   g004(.A(G211gat), .B(G218gat), .Z(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G197gat), .B(G204gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT21), .ZN(new_n209_));
  NOR3_X1   g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(KEYINPUT21), .B1(new_n208_), .B2(KEYINPUT85), .ZN(new_n211_));
  INV_X1    g010(.A(G204gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(G197gat), .ZN(new_n213_));
  INV_X1    g012(.A(G197gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(G204gat), .ZN(new_n215_));
  AND4_X1   g014(.A1(KEYINPUT85), .A2(new_n213_), .A3(new_n215_), .A4(KEYINPUT21), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n207_), .B1(new_n211_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT86), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n213_), .A2(new_n215_), .A3(KEYINPUT85), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n209_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n208_), .A2(KEYINPUT85), .A3(KEYINPUT21), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(KEYINPUT86), .A3(new_n207_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n210_), .B1(new_n219_), .B2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT91), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n226_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT22), .B(G169gat), .ZN(new_n230_));
  INV_X1    g029(.A(G176gat), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n229_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n228_), .B1(new_n232_), .B2(new_n227_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT92), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT92), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n235_), .B(new_n228_), .C1(new_n232_), .C2(new_n227_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G183gat), .A2(G190gat), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n237_), .B(KEYINPUT23), .Z(new_n238_));
  NOR2_X1   g037(.A1(G183gat), .A2(G190gat), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n234_), .B(new_n236_), .C1(new_n238_), .C2(new_n239_), .ZN(new_n240_));
  OR2_X1    g039(.A1(G169gat), .A2(G176gat), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n241_), .A2(KEYINPUT24), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n241_), .A2(KEYINPUT24), .A3(new_n226_), .ZN(new_n243_));
  NOR3_X1   g042(.A1(new_n238_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT26), .B(G190gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT25), .B(G183gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n244_), .A2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n225_), .B1(new_n240_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n210_), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT86), .B1(new_n223_), .B2(new_n207_), .ZN(new_n251_));
  AOI211_X1 g050(.A(new_n218_), .B(new_n206_), .C1(new_n221_), .C2(new_n222_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n250_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT25), .ZN(new_n254_));
  NOR2_X1   g053(.A1(KEYINPUT79), .A2(G183gat), .ZN(new_n255_));
  AND2_X1   g054(.A1(KEYINPUT79), .A2(G183gat), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT80), .ZN(new_n257_));
  AOI211_X1 g056(.A(new_n254_), .B(new_n255_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(new_n254_), .A3(G183gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n245_), .A2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT81), .B1(new_n258_), .B2(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n255_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT25), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT81), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n263_), .A2(new_n264_), .A3(new_n259_), .A4(new_n245_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n244_), .A2(new_n261_), .A3(new_n265_), .ZN(new_n266_));
  NOR3_X1   g065(.A1(new_n256_), .A2(new_n255_), .A3(G190gat), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n232_), .B1(new_n238_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT20), .B1(new_n253_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G226gat), .A2(G233gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT19), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NOR3_X1   g072(.A1(new_n249_), .A2(new_n270_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT20), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n275_), .B1(new_n253_), .B2(new_n269_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n240_), .A2(new_n225_), .A3(new_n248_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n272_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n205_), .B1(new_n274_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n278_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n240_), .A2(new_n248_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n253_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n225_), .A2(new_n268_), .A3(new_n266_), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n282_), .A2(new_n283_), .A3(KEYINPUT20), .A4(new_n272_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n205_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n280_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT93), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n279_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n280_), .A2(KEYINPUT93), .A3(new_n284_), .A4(new_n285_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n290_), .A2(KEYINPUT27), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G225gat), .A2(G233gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT94), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT4), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G141gat), .A2(G148gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(G141gat), .A2(G148gat), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(G155gat), .ZN(new_n299_));
  INV_X1    g098(.A(G162gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n299_), .A2(new_n300_), .A3(KEYINPUT83), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT83), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n302_), .B1(G155gat), .B2(G162gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT1), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT84), .B1(new_n305_), .B2(KEYINPUT1), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT84), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT1), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n309_), .A2(new_n310_), .A3(G155gat), .A4(G162gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n298_), .B1(new_n307_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT3), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n297_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT2), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n295_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n315_), .A2(new_n317_), .A3(new_n318_), .A4(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n320_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n313_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(G120gat), .ZN(new_n323_));
  INV_X1    g122(.A(G127gat), .ZN(new_n324_));
  INV_X1    g123(.A(G134gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(G113gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G127gat), .A2(G134gat), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n327_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n323_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n331_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n333_), .A2(G120gat), .A3(new_n329_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT95), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n322_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n313_), .A2(new_n334_), .A3(new_n332_), .A4(new_n321_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n294_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n313_), .A2(new_n321_), .B1(new_n332_), .B2(new_n334_), .ZN(new_n340_));
  AOI21_X1  g139(.A(KEYINPUT4), .B1(new_n340_), .B2(new_n336_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n293_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n322_), .A2(new_n335_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n343_), .A2(new_n340_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n293_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n342_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT97), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G1gat), .B(G29gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G57gat), .B(G85gat), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n351_), .B(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n347_), .A2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n342_), .A2(new_n346_), .A3(new_n354_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n356_), .A2(KEYINPUT99), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT99), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n347_), .A2(new_n359_), .A3(new_n355_), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n249_), .A2(new_n270_), .A3(new_n272_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n273_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n285_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n279_), .A2(new_n365_), .A3(KEYINPUT27), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n291_), .A2(new_n362_), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT90), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n322_), .A2(KEYINPUT29), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G22gat), .B(G50gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT28), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n370_), .B(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(G228gat), .ZN(new_n375_));
  INV_X1    g174(.A(G233gat), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT87), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n321_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n298_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n308_), .A2(new_n311_), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n301_), .A2(new_n303_), .B1(KEYINPUT1), .B2(new_n305_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n380_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT29), .B1(new_n379_), .B2(new_n383_), .ZN(new_n384_));
  NOR3_X1   g183(.A1(new_n375_), .A2(new_n376_), .A3(KEYINPUT87), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n378_), .B1(new_n387_), .B2(new_n225_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n385_), .B1(new_n322_), .B2(KEYINPUT29), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n253_), .A2(new_n389_), .A3(new_n377_), .ZN(new_n390_));
  XOR2_X1   g189(.A(G78gat), .B(G106gat), .Z(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n388_), .A2(new_n390_), .A3(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n392_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n393_), .B1(new_n394_), .B2(KEYINPUT88), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT88), .ZN(new_n396_));
  AOI211_X1 g195(.A(new_n396_), .B(new_n392_), .C1(new_n388_), .C2(new_n390_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n374_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT89), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT89), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n400_), .B(new_n374_), .C1(new_n395_), .C2(new_n397_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n253_), .A2(new_n389_), .A3(new_n377_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n377_), .B1(new_n253_), .B2(new_n389_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n391_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n405_), .A2(new_n373_), .A3(new_n393_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n369_), .B1(new_n402_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n406_), .ZN(new_n408_));
  AOI211_X1 g207(.A(KEYINPUT90), .B(new_n408_), .C1(new_n399_), .C2(new_n401_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n269_), .B(new_n335_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT82), .B(KEYINPUT30), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G71gat), .B(G99gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT31), .ZN(new_n414_));
  XOR2_X1   g213(.A(G15gat), .B(G43gat), .Z(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G227gat), .A2(G233gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n412_), .B(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NOR3_X1   g219(.A1(new_n407_), .A2(new_n409_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n401_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n405_), .A2(new_n396_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n394_), .A2(KEYINPUT88), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(new_n424_), .A3(new_n393_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n400_), .B1(new_n425_), .B2(new_n374_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n406_), .B1(new_n422_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT90), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n402_), .A2(new_n369_), .A3(new_n406_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n419_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n368_), .B1(new_n421_), .B2(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n407_), .A2(new_n409_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT100), .ZN(new_n433_));
  OAI211_X1 g232(.A(KEYINPUT32), .B(new_n205_), .C1(new_n363_), .C2(new_n364_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n435_), .B1(new_n274_), .B2(new_n278_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n361_), .A2(new_n433_), .A3(new_n434_), .A4(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n345_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n355_), .A2(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n439_), .B1(new_n293_), .B2(new_n344_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT33), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n357_), .A2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n357_), .A2(KEYINPUT98), .A3(new_n441_), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT98), .B1(new_n357_), .B2(new_n441_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n290_), .A2(new_n443_), .A3(new_n446_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n358_), .A2(new_n360_), .A3(new_n434_), .A4(new_n436_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT100), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n437_), .A2(new_n447_), .A3(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n432_), .A2(new_n420_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n431_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(G57gat), .ZN(new_n453_));
  INV_X1    g252(.A(G64gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT11), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G57gat), .A2(G64gat), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G71gat), .A2(G78gat), .ZN(new_n459_));
  INV_X1    g258(.A(G71gat), .ZN(new_n460_));
  INV_X1    g259(.A(G78gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n458_), .A2(new_n459_), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT66), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n456_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT66), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n458_), .A2(new_n466_), .A3(new_n459_), .A4(new_n462_), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n464_), .A2(new_n465_), .A3(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n465_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(G85gat), .ZN(new_n471_));
  INV_X1    g270(.A(G92gat), .ZN(new_n472_));
  NOR3_X1   g271(.A1(new_n471_), .A2(new_n472_), .A3(KEYINPUT9), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G99gat), .A2(G106gat), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT6), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  XOR2_X1   g277(.A(G85gat), .B(G92gat), .Z(new_n479_));
  AOI211_X1 g278(.A(new_n473_), .B(new_n478_), .C1(KEYINPUT9), .C2(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(KEYINPUT10), .B(G99gat), .Z(new_n481_));
  INV_X1    g280(.A(G106gat), .ZN(new_n482_));
  AOI21_X1  g281(.A(KEYINPUT64), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n481_), .A2(KEYINPUT64), .A3(new_n482_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n480_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT7), .ZN(new_n486_));
  INV_X1    g285(.A(G99gat), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n486_), .A2(new_n487_), .A3(new_n482_), .A4(KEYINPUT65), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT65), .ZN(new_n489_));
  OAI22_X1  g288(.A1(new_n489_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(KEYINPUT7), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n476_), .A2(new_n477_), .A3(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n479_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT8), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT8), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n496_), .B(new_n479_), .C1(new_n491_), .C2(new_n493_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n485_), .A2(new_n498_), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n470_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n470_), .A2(new_n499_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G230gat), .A2(G233gat), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n498_), .A2(KEYINPUT67), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT67), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n495_), .A2(new_n507_), .A3(new_n497_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n506_), .A2(new_n485_), .A3(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n509_), .A2(KEYINPUT12), .A3(new_n470_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT12), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n501_), .A2(new_n511_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n510_), .A2(new_n512_), .A3(new_n503_), .A4(new_n500_), .ZN(new_n513_));
  XOR2_X1   g312(.A(G120gat), .B(G148gat), .Z(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G176gat), .B(G204gat), .ZN(new_n517_));
  XOR2_X1   g316(.A(new_n516_), .B(new_n517_), .Z(new_n518_));
  NAND3_X1  g317(.A1(new_n505_), .A2(new_n513_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n518_), .B1(new_n505_), .B2(new_n513_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  AND2_X1   g322(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n523_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G169gat), .B(G197gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(G141gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT77), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(new_n327_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G15gat), .B(G22gat), .ZN(new_n534_));
  INV_X1    g333(.A(G1gat), .ZN(new_n535_));
  INV_X1    g334(.A(G8gat), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT14), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n534_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G1gat), .B(G8gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G29gat), .B(G36gat), .ZN(new_n541_));
  INV_X1    g340(.A(G43gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(G50gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n541_), .B(G43gat), .ZN(new_n545_));
  INV_X1    g344(.A(G50gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n544_), .A2(new_n547_), .A3(KEYINPUT15), .ZN(new_n548_));
  AOI21_X1  g347(.A(KEYINPUT15), .B1(new_n544_), .B2(new_n547_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n540_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT75), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G229gat), .A2(G233gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n544_), .A2(new_n547_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n553_), .A2(new_n540_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT75), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n555_), .B(new_n540_), .C1(new_n548_), .C2(new_n549_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n551_), .A2(new_n552_), .A3(new_n554_), .A4(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n553_), .B(new_n540_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n552_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n557_), .A2(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n533_), .B1(new_n561_), .B2(KEYINPUT76), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n562_), .B1(KEYINPUT76), .B2(new_n561_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n557_), .A2(new_n560_), .A3(new_n533_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT78), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT78), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n557_), .A2(new_n560_), .A3(new_n566_), .A4(new_n533_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n563_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n529_), .A2(new_n570_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n452_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G232gat), .A2(G233gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT70), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT34), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(KEYINPUT35), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n499_), .A2(new_n553_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n509_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n578_), .B1(new_n579_), .B2(KEYINPUT71), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n579_), .A2(KEYINPUT71), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n576_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n575_), .B(KEYINPUT35), .Z(new_n583_));
  NAND3_X1  g382(.A1(new_n579_), .A2(new_n577_), .A3(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n582_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT72), .B(G190gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(G218gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G134gat), .B(G162gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n590_), .A2(KEYINPUT36), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n586_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT73), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT37), .ZN(new_n594_));
  INV_X1    g393(.A(new_n586_), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n590_), .B(KEYINPUT36), .Z(new_n596_));
  AOI21_X1  g395(.A(new_n594_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n593_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n540_), .B(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(new_n470_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(KEYINPUT16), .B(G183gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(G211gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G127gat), .B(G155gat), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n603_), .B(new_n604_), .Z(new_n605_));
  INV_X1    g404(.A(KEYINPUT17), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n605_), .A2(new_n606_), .ZN(new_n608_));
  NOR3_X1   g407(.A1(new_n601_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n609_), .B1(new_n607_), .B2(new_n601_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n586_), .A2(KEYINPUT74), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT74), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n612_), .B1(new_n582_), .B2(new_n585_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n611_), .A2(new_n596_), .A3(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(new_n592_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n594_), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n598_), .A2(new_n610_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n572_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n619_), .A2(new_n535_), .A3(new_n361_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT38), .ZN(new_n621_));
  INV_X1    g420(.A(new_n615_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n610_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n572_), .A2(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(G1gat), .B1(new_n625_), .B2(new_n362_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n621_), .A2(new_n626_), .ZN(G1324gat));
  NAND2_X1  g426(.A1(new_n291_), .A2(new_n366_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(G8gat), .B1(new_n625_), .B2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT39), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n619_), .A2(new_n536_), .A3(new_n628_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g433(.A(G15gat), .B1(new_n625_), .B2(new_n420_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT41), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n618_), .A2(G15gat), .A3(new_n420_), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n636_), .A2(new_n637_), .ZN(G1326gat));
  XOR2_X1   g437(.A(new_n432_), .B(KEYINPUT101), .Z(new_n639_));
  OAI21_X1  g438(.A(G22gat), .B1(new_n625_), .B2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT42), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n639_), .A2(G22gat), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n641_), .B1(new_n618_), .B2(new_n642_), .ZN(G1327gat));
  NAND2_X1  g442(.A1(new_n622_), .A2(new_n623_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT104), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n645_), .A2(new_n452_), .A3(new_n571_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT105), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n572_), .A2(KEYINPUT105), .A3(new_n645_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  OR3_X1    g449(.A1(new_n650_), .A2(G29gat), .A3(new_n362_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT43), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n598_), .A2(new_n616_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n452_), .A2(KEYINPUT102), .A3(new_n652_), .A4(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n420_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n428_), .A2(new_n429_), .A3(new_n419_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n367_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  AND4_X1   g456(.A1(new_n428_), .A2(new_n450_), .A3(new_n429_), .A4(new_n420_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n652_), .B(new_n653_), .C1(new_n657_), .C2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n653_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(KEYINPUT43), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n654_), .A2(new_n661_), .A3(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n664_), .A2(new_n571_), .A3(new_n623_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n664_), .A2(KEYINPUT44), .A3(new_n571_), .A4(new_n623_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(new_n361_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n670_), .A2(new_n671_), .A3(G29gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n670_), .B2(G29gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n651_), .B1(new_n672_), .B2(new_n673_), .ZN(G1328gat));
  INV_X1    g473(.A(G36gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n669_), .B2(new_n628_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n628_), .B(KEYINPUT106), .Z(new_n678_));
  NAND4_X1  g477(.A1(new_n648_), .A2(new_n649_), .A3(new_n675_), .A4(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n679_), .A2(KEYINPUT107), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(KEYINPUT107), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n681_), .A2(new_n682_), .A3(KEYINPUT45), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT45), .ZN(new_n684_));
  INV_X1    g483(.A(new_n682_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n684_), .B1(new_n685_), .B2(new_n680_), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n677_), .A2(KEYINPUT46), .A3(new_n683_), .A4(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT46), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n683_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(new_n676_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n687_), .A2(new_n690_), .ZN(G1329gat));
  NAND4_X1  g490(.A1(new_n667_), .A2(G43gat), .A3(new_n419_), .A4(new_n668_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT108), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n542_), .B1(new_n650_), .B2(new_n420_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n692_), .A2(new_n693_), .A3(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n693_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT47), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n696_), .A2(new_n697_), .A3(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n692_), .A2(new_n694_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT108), .ZN(new_n701_));
  AOI21_X1  g500(.A(KEYINPUT47), .B1(new_n701_), .B2(new_n695_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n699_), .A2(new_n702_), .ZN(G1330gat));
  INV_X1    g502(.A(new_n432_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n669_), .A2(G50gat), .A3(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n546_), .B1(new_n650_), .B2(new_n639_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1331gat));
  AOI211_X1 g506(.A(new_n528_), .B(new_n569_), .C1(new_n431_), .C2(new_n451_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n624_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n709_), .A2(new_n453_), .A3(new_n362_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n617_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n361_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n710_), .B1(new_n453_), .B2(new_n713_), .ZN(G1332gat));
  INV_X1    g513(.A(new_n709_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n454_), .B1(new_n715_), .B2(new_n678_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT48), .Z(new_n717_));
  NAND3_X1  g516(.A1(new_n712_), .A2(new_n454_), .A3(new_n678_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT109), .ZN(G1333gat));
  OAI21_X1  g519(.A(G71gat), .B1(new_n709_), .B2(new_n420_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT49), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n712_), .A2(new_n460_), .A3(new_n419_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT110), .Z(G1334gat));
  OAI21_X1  g524(.A(G78gat), .B1(new_n709_), .B2(new_n639_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT50), .ZN(new_n727_));
  INV_X1    g526(.A(new_n639_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n712_), .A2(new_n461_), .A3(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1335gat));
  NOR3_X1   g529(.A1(new_n528_), .A2(new_n569_), .A3(new_n610_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n664_), .A2(new_n731_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n732_), .A2(new_n471_), .A3(new_n362_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n708_), .A2(new_n645_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT111), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(new_n361_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n733_), .B1(new_n736_), .B2(new_n471_), .ZN(G1336gat));
  AOI21_X1  g536(.A(G92gat), .B1(new_n735_), .B2(new_n628_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n732_), .A2(new_n472_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n678_), .B2(new_n739_), .ZN(G1337gat));
  NAND3_X1  g539(.A1(new_n735_), .A2(new_n481_), .A3(new_n419_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G99gat), .B1(new_n732_), .B2(new_n420_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g543(.A1(new_n664_), .A2(new_n704_), .A3(new_n731_), .ZN(new_n745_));
  XOR2_X1   g544(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n745_), .A2(G106gat), .A3(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT113), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT113), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n745_), .A2(new_n750_), .A3(G106gat), .A4(new_n747_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT114), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n745_), .A2(G106gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n754_), .B2(new_n746_), .ZN(new_n755_));
  AOI211_X1 g554(.A(KEYINPUT114), .B(new_n747_), .C1(new_n745_), .C2(G106gat), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n752_), .A2(new_n755_), .A3(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n735_), .A2(new_n482_), .A3(new_n704_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(KEYINPUT53), .B1(new_n757_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT53), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n755_), .A2(new_n756_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n761_), .B(new_n758_), .C1(new_n762_), .C2(new_n752_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n760_), .A2(new_n763_), .ZN(G1339gat));
  INV_X1    g563(.A(KEYINPUT57), .ZN(new_n765_));
  INV_X1    g564(.A(new_n518_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT55), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n510_), .A2(new_n512_), .A3(new_n500_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(new_n504_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n513_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n768_), .A2(new_n767_), .A3(new_n504_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n766_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT56), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  OAI211_X1 g574(.A(KEYINPUT56), .B(new_n766_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(KEYINPUT116), .A3(new_n776_), .ZN(new_n777_));
  OR2_X1    g576(.A1(new_n776_), .A2(KEYINPUT116), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n777_), .A2(new_n778_), .A3(new_n519_), .A4(new_n569_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT118), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n551_), .A2(new_n554_), .A3(new_n556_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT117), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT117), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n551_), .A2(new_n783_), .A3(new_n554_), .A4(new_n556_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n782_), .A2(new_n559_), .A3(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n533_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n558_), .A2(new_n552_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n785_), .A2(new_n786_), .A3(new_n787_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n788_), .A2(new_n568_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n780_), .B1(new_n789_), .B2(new_n523_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n568_), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n791_), .A2(KEYINPUT118), .A3(new_n522_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  AOI211_X1 g592(.A(new_n765_), .B(new_n622_), .C1(new_n779_), .C2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n775_), .A2(KEYINPUT120), .A3(new_n776_), .ZN(new_n795_));
  OR2_X1    g594(.A1(new_n776_), .A2(KEYINPUT120), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n795_), .A2(new_n796_), .A3(new_n519_), .A4(new_n789_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT58), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(KEYINPUT121), .A3(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n798_), .B1(new_n797_), .B2(KEYINPUT121), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n794_), .B1(new_n802_), .B2(new_n653_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n779_), .A2(new_n793_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n615_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n765_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n803_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n623_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT123), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  AND2_X1   g609(.A1(KEYINPUT115), .A2(KEYINPUT54), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n617_), .A2(new_n528_), .A3(new_n570_), .A4(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(KEYINPUT115), .A2(KEYINPUT54), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n811_), .A2(new_n813_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n598_), .A2(new_n528_), .A3(new_n616_), .A4(new_n610_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n814_), .B1(new_n815_), .B2(new_n569_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n812_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n807_), .A2(KEYINPUT123), .A3(new_n623_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n810_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT59), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n656_), .A2(new_n362_), .A3(new_n628_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n820_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT122), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT119), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n825_), .B1(new_n805_), .B2(new_n765_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n622_), .B1(new_n779_), .B2(new_n793_), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n827_), .A2(KEYINPUT119), .A3(KEYINPUT57), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n610_), .B1(new_n829_), .B2(new_n803_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n824_), .B1(new_n830_), .B2(new_n817_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n801_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(new_n653_), .A3(new_n799_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n805_), .A2(new_n825_), .A3(new_n765_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n794_), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT119), .B1(new_n827_), .B2(KEYINPUT57), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n833_), .A2(new_n834_), .A3(new_n835_), .A4(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n623_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n838_), .A2(KEYINPUT122), .A3(new_n818_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n831_), .A2(new_n839_), .A3(new_n822_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT59), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n823_), .A2(new_n841_), .A3(G113gat), .A4(new_n569_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n327_), .B1(new_n840_), .B2(new_n570_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n842_), .A2(new_n843_), .ZN(G1340gat));
  XOR2_X1   g643(.A(KEYINPUT124), .B(G120gat), .Z(new_n845_));
  INV_X1    g644(.A(KEYINPUT60), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n831_), .A2(new_n839_), .A3(new_n822_), .A4(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n845_), .B1(new_n529_), .B2(new_n846_), .ZN(new_n849_));
  OR3_X1    g648(.A1(new_n848_), .A2(KEYINPUT125), .A3(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(KEYINPUT125), .B1(new_n848_), .B2(new_n849_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n823_), .A2(new_n841_), .A3(new_n529_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n845_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n854_), .ZN(G1341gat));
  NAND4_X1  g654(.A1(new_n823_), .A2(new_n841_), .A3(G127gat), .A4(new_n610_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n324_), .B1(new_n840_), .B2(new_n623_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(G1342gat));
  NAND4_X1  g657(.A1(new_n823_), .A2(new_n841_), .A3(G134gat), .A4(new_n653_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n325_), .B1(new_n840_), .B2(new_n615_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n859_), .A2(new_n860_), .ZN(G1343gat));
  NOR2_X1   g660(.A1(new_n678_), .A2(new_n655_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n831_), .A2(new_n361_), .A3(new_n839_), .A4(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(new_n570_), .ZN(new_n864_));
  XOR2_X1   g663(.A(new_n864_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g664(.A1(new_n863_), .A2(new_n528_), .ZN(new_n866_));
  XOR2_X1   g665(.A(new_n866_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g666(.A1(new_n863_), .A2(new_n623_), .ZN(new_n868_));
  XOR2_X1   g667(.A(KEYINPUT61), .B(G155gat), .Z(new_n869_));
  XNOR2_X1  g668(.A(new_n868_), .B(new_n869_), .ZN(G1346gat));
  AOI21_X1  g669(.A(KEYINPUT122), .B1(new_n838_), .B2(new_n818_), .ZN(new_n871_));
  AOI211_X1 g670(.A(new_n824_), .B(new_n817_), .C1(new_n837_), .C2(new_n623_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n871_), .A2(new_n872_), .A3(new_n362_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n873_), .A2(new_n300_), .A3(new_n622_), .A4(new_n862_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n653_), .ZN(new_n875_));
  OAI21_X1  g674(.A(G162gat), .B1(new_n863_), .B2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT126), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT126), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n874_), .A2(new_n876_), .A3(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n880_), .ZN(G1347gat));
  AND2_X1   g680(.A1(new_n678_), .A2(new_n362_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n419_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(new_n728_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n820_), .A2(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(G169gat), .B1(new_n885_), .B2(new_n570_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n885_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n889_), .A2(new_n569_), .A3(new_n230_), .ZN(new_n890_));
  OAI211_X1 g689(.A(KEYINPUT62), .B(G169gat), .C1(new_n885_), .C2(new_n570_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n888_), .A2(new_n890_), .A3(new_n891_), .ZN(G1348gat));
  AOI21_X1  g691(.A(G176gat), .B1(new_n889_), .B2(new_n529_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n871_), .A2(new_n872_), .A3(new_n704_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n883_), .A2(new_n231_), .A3(new_n528_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n894_), .B2(new_n895_), .ZN(G1349gat));
  NOR3_X1   g695(.A1(new_n885_), .A2(new_n246_), .A3(new_n623_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n256_), .A2(new_n255_), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n894_), .A2(new_n419_), .A3(new_n610_), .A4(new_n882_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n897_), .B1(new_n898_), .B2(new_n899_), .ZN(G1350gat));
  NAND3_X1  g699(.A1(new_n889_), .A2(new_n245_), .A3(new_n622_), .ZN(new_n901_));
  OAI21_X1  g700(.A(G190gat), .B1(new_n885_), .B2(new_n875_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1351gat));
  NAND4_X1  g702(.A1(new_n831_), .A2(new_n430_), .A3(new_n839_), .A4(new_n882_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n570_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(new_n214_), .ZN(G1352gat));
  NOR2_X1   g705(.A1(new_n904_), .A2(new_n528_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(new_n212_), .ZN(G1353gat));
  OR2_X1    g707(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n909_));
  XNOR2_X1  g708(.A(KEYINPUT63), .B(G211gat), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n904_), .A2(new_n623_), .ZN(new_n911_));
  MUX2_X1   g710(.A(new_n909_), .B(new_n910_), .S(new_n911_), .Z(G1354gat));
  INV_X1    g711(.A(G218gat), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n904_), .A2(new_n913_), .A3(new_n875_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n871_), .A2(new_n872_), .A3(new_n655_), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n915_), .A2(KEYINPUT127), .A3(new_n622_), .A4(new_n882_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT127), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n917_), .B1(new_n904_), .B2(new_n615_), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n916_), .A2(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n914_), .B1(new_n919_), .B2(new_n913_), .ZN(G1355gat));
endmodule


