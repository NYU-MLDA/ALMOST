//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 0 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n881_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n913_, new_n915_, new_n916_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT82), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT1), .ZN(new_n207_));
  INV_X1    g006(.A(G155gat), .ZN(new_n208_));
  INV_X1    g007(.A(G162gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n208_), .A2(new_n209_), .A3(KEYINPUT83), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT83), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n211_), .B1(G155gat), .B2(G162gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n204_), .B(new_n205_), .C1(new_n207_), .C2(new_n213_), .ZN(new_n214_));
  AND3_X1   g013(.A1(new_n210_), .A2(new_n212_), .A3(new_n206_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n203_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT2), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n205_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n217_), .A2(new_n219_), .A3(new_n220_), .A4(new_n221_), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n215_), .A2(new_n222_), .A3(KEYINPUT84), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT84), .B1(new_n215_), .B2(new_n222_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n214_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G127gat), .B(G134gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G113gat), .B(G120gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n226_), .B(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n225_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n225_), .A2(KEYINPUT85), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT85), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n233_), .B(new_n214_), .C1(new_n223_), .C2(new_n224_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n228_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT4), .B1(new_n231_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n232_), .A2(new_n234_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(new_n229_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT4), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n202_), .B1(new_n236_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n238_), .A2(new_n230_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n202_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(G57gat), .B(G85gat), .Z(new_n245_));
  XNOR2_X1  g044(.A(G1gat), .B(G29gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NOR3_X1   g049(.A1(new_n241_), .A2(new_n244_), .A3(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT33), .B1(new_n251_), .B2(KEYINPUT95), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G8gat), .B(G36gat), .ZN(new_n253_));
  INV_X1    g052(.A(G92gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT18), .B(G64gat), .ZN(new_n256_));
  XOR2_X1   g055(.A(new_n255_), .B(new_n256_), .Z(new_n257_));
  INV_X1    g056(.A(KEYINPUT20), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT25), .B(G183gat), .ZN(new_n259_));
  INV_X1    g058(.A(G190gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT26), .B1(new_n260_), .B2(KEYINPUT74), .ZN(new_n261_));
  OR2_X1    g060(.A1(new_n260_), .A2(KEYINPUT26), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n259_), .B(new_n261_), .C1(new_n262_), .C2(KEYINPUT74), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT75), .B1(G169gat), .B2(G176gat), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NOR3_X1   g065(.A1(KEYINPUT75), .A2(G169gat), .A3(G176gat), .ZN(new_n267_));
  OAI211_X1 g066(.A(KEYINPUT24), .B(new_n264_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n267_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT24), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n269_), .A2(new_n270_), .A3(new_n265_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT23), .ZN(new_n272_));
  INV_X1    g071(.A(G183gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n272_), .B1(new_n273_), .B2(new_n260_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n263_), .A2(new_n268_), .A3(new_n271_), .A4(new_n276_), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n274_), .B(new_n275_), .C1(G183gat), .C2(G190gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT77), .B(G176gat), .ZN(new_n279_));
  INV_X1    g078(.A(G169gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT22), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n279_), .B1(KEYINPUT76), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(KEYINPUT76), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n280_), .A2(KEYINPUT22), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n264_), .B(new_n278_), .C1(new_n282_), .C2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n277_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT78), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT78), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n277_), .A2(new_n286_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(G211gat), .B(G218gat), .Z(new_n292_));
  INV_X1    g091(.A(G204gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(G197gat), .ZN(new_n294_));
  INV_X1    g093(.A(G197gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G204gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n292_), .A2(KEYINPUT21), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n292_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT87), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n294_), .A2(new_n296_), .A3(new_n301_), .A4(KEYINPUT21), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT87), .B1(new_n295_), .B2(G204gat), .ZN(new_n304_));
  AOI22_X1  g103(.A1(new_n304_), .A2(KEYINPUT21), .B1(new_n294_), .B2(new_n296_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n300_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT88), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT88), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n308_), .B(new_n300_), .C1(new_n303_), .C2(new_n305_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n299_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n258_), .B1(new_n291_), .B2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G226gat), .A2(G233gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n268_), .A2(new_n276_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(G176gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n270_), .A2(new_n280_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n259_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT26), .B(G190gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT92), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n318_), .B(new_n320_), .C1(new_n321_), .C2(new_n323_), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n284_), .A2(new_n281_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(new_n279_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n264_), .B(KEYINPUT93), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n326_), .A2(new_n278_), .A3(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n310_), .A2(new_n324_), .A3(new_n328_), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n312_), .A2(new_n316_), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n324_), .A2(new_n328_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n258_), .B1(new_n311_), .B2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n310_), .A2(new_n288_), .A3(new_n290_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n316_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n257_), .B1(new_n330_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n332_), .A2(new_n333_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n315_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n257_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n312_), .A2(new_n316_), .A3(new_n329_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n335_), .A2(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n243_), .B1(new_n236_), .B2(new_n240_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n242_), .A2(new_n202_), .ZN(new_n343_));
  NOR3_X1   g142(.A1(new_n342_), .A2(new_n343_), .A3(new_n249_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n341_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n236_), .A2(new_n240_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(new_n243_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n244_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n347_), .A2(new_n348_), .A3(new_n249_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT95), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT33), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n349_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n252_), .A2(new_n345_), .A3(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n338_), .A2(KEYINPUT32), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n337_), .A2(new_n354_), .A3(new_n339_), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n332_), .A2(new_n316_), .A3(new_n333_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n316_), .B1(new_n312_), .B2(new_n329_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n249_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n359_));
  OAI221_X1 g158(.A(new_n355_), .B1(new_n354_), .B2(new_n358_), .C1(new_n359_), .C2(new_n251_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n353_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT90), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G22gat), .B(G50gat), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT28), .B1(new_n237_), .B2(KEYINPUT29), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT28), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT29), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n232_), .A2(new_n365_), .A3(new_n366_), .A4(new_n234_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n363_), .B1(new_n364_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n364_), .A2(new_n367_), .A3(new_n363_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n237_), .A2(KEYINPUT29), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT86), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(G228gat), .ZN(new_n375_));
  INV_X1    g174(.A(G233gat), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n366_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n377_), .B1(new_n378_), .B2(KEYINPUT86), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n374_), .A2(new_n379_), .A3(new_n311_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n225_), .A2(KEYINPUT29), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n377_), .B1(new_n381_), .B2(new_n310_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT89), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT89), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n384_), .B(new_n377_), .C1(new_n381_), .C2(new_n310_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G78gat), .B(G106gat), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n380_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n387_), .B1(new_n380_), .B2(new_n386_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n362_), .B(new_n371_), .C1(new_n388_), .C2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n380_), .A2(new_n386_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n387_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n370_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n362_), .B1(new_n394_), .B2(new_n368_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n369_), .A2(KEYINPUT90), .A3(new_n370_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n380_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n393_), .A2(new_n395_), .A3(new_n396_), .A4(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n390_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n361_), .A2(new_n399_), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n390_), .A2(new_n398_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT96), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n359_), .A2(new_n251_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n257_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n404_), .A2(new_n340_), .A3(KEYINPUT27), .ZN(new_n405_));
  AOI21_X1  g204(.A(KEYINPUT27), .B1(new_n335_), .B2(new_n340_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n401_), .A2(new_n402_), .A3(new_n403_), .A4(new_n407_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n407_), .A2(new_n403_), .A3(new_n390_), .A4(new_n398_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT96), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n400_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G227gat), .A2(G233gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(G15gat), .ZN(new_n413_));
  INV_X1    g212(.A(G43gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  XOR2_X1   g214(.A(G71gat), .B(G99gat), .Z(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT30), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n291_), .B(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT79), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n420_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n417_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n423_), .B1(new_n421_), .B2(new_n417_), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n228_), .B(KEYINPUT81), .Z(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT31), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n426_), .A2(KEYINPUT80), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n424_), .B(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n403_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT97), .ZN(new_n431_));
  INV_X1    g230(.A(new_n407_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n431_), .B1(new_n401_), .B2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n399_), .A2(KEYINPUT97), .A3(new_n407_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  AOI22_X1  g234(.A1(new_n411_), .A2(new_n428_), .B1(new_n430_), .B2(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(KEYINPUT71), .B(G8gat), .Z(new_n437_));
  INV_X1    g236(.A(G1gat), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT14), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(G8gat), .ZN(new_n440_));
  XOR2_X1   g239(.A(G15gat), .B(G22gat), .Z(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n439_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT14), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT71), .B(G8gat), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n444_), .B1(new_n445_), .B2(G1gat), .ZN(new_n446_));
  OAI21_X1  g245(.A(G8gat), .B1(new_n446_), .B2(new_n441_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n443_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(KEYINPUT72), .B(G1gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n443_), .A2(new_n447_), .A3(new_n449_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G231gat), .A2(G233gat), .ZN(new_n454_));
  XOR2_X1   g253(.A(new_n453_), .B(new_n454_), .Z(new_n455_));
  OR2_X1    g254(.A1(G57gat), .A2(G64gat), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT11), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G57gat), .A2(G64gat), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  AND2_X1   g258(.A1(G57gat), .A2(G64gat), .ZN(new_n460_));
  NOR2_X1   g259(.A1(G57gat), .A2(G64gat), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT11), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(G78gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(G71gat), .ZN(new_n464_));
  INV_X1    g263(.A(G71gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(G78gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n459_), .A2(new_n462_), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n456_), .A2(new_n458_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n469_), .A2(KEYINPUT11), .A3(new_n464_), .A4(new_n466_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(new_n455_), .B(new_n471_), .Z(new_n472_));
  XOR2_X1   g271(.A(G127gat), .B(G155gat), .Z(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(G211gat), .ZN(new_n474_));
  XOR2_X1   g273(.A(KEYINPUT16), .B(G183gat), .Z(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n472_), .A2(KEYINPUT17), .A3(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n471_), .A2(KEYINPUT65), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT65), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n468_), .A2(new_n470_), .A3(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n455_), .B(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(new_n476_), .B(KEYINPUT17), .Z(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n477_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n436_), .A2(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(KEYINPUT10), .B(G99gat), .Z(new_n488_));
  INV_X1    g287(.A(G106gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G85gat), .A2(G92gat), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n491_), .A2(KEYINPUT9), .ZN(new_n492_));
  INV_X1    g291(.A(G85gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n254_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n494_), .A2(KEYINPUT9), .A3(new_n491_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n490_), .A2(new_n492_), .A3(new_n495_), .A4(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT7), .ZN(new_n501_));
  INV_X1    g300(.A(G99gat), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n501_), .A2(new_n502_), .A3(new_n489_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G99gat), .A2(G106gat), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT6), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n503_), .A2(new_n506_), .A3(new_n496_), .A4(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT8), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n494_), .A2(new_n491_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n509_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n500_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT67), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT67), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n500_), .B(new_n516_), .C1(new_n512_), .C2(new_n513_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G29gat), .B(G36gat), .ZN(new_n519_));
  INV_X1    g318(.A(G50gat), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n520_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(KEYINPUT70), .B(G43gat), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n521_), .A2(new_n522_), .A3(new_n524_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n526_), .A2(KEYINPUT15), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT15), .ZN(new_n529_));
  INV_X1    g328(.A(new_n527_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n524_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n529_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  AND3_X1   g331(.A1(new_n518_), .A2(new_n528_), .A3(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n530_), .A2(new_n531_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G232gat), .A2(G233gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT34), .ZN(new_n536_));
  OAI22_X1  g335(.A1(new_n534_), .A2(new_n514_), .B1(KEYINPUT35), .B2(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n533_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(KEYINPUT35), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  OAI211_X1 g339(.A(KEYINPUT35), .B(new_n536_), .C1(new_n533_), .C2(new_n537_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G190gat), .B(G218gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G134gat), .B(G162gat), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n543_), .B(new_n544_), .Z(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT36), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n542_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT36), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n545_), .A2(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n542_), .A2(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(KEYINPUT37), .B1(new_n548_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT37), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n547_), .B(new_n553_), .C1(new_n550_), .C2(new_n542_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n487_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G113gat), .B(G141gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G169gat), .B(G197gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n534_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n453_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n453_), .A2(new_n560_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G229gat), .A2(G233gat), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n451_), .A2(new_n532_), .A3(new_n452_), .A4(new_n528_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n561_), .A2(new_n567_), .A3(new_n565_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n559_), .B1(new_n566_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT73), .ZN(new_n571_));
  INV_X1    g370(.A(new_n559_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n568_), .B(new_n572_), .C1(new_n564_), .C2(new_n565_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n570_), .A2(new_n571_), .A3(new_n573_), .ZN(new_n574_));
  OAI211_X1 g373(.A(KEYINPUT73), .B(new_n559_), .C1(new_n566_), .C2(new_n569_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G230gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT64), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n468_), .A2(new_n479_), .A3(new_n470_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n479_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n579_), .B1(new_n582_), .B2(new_n514_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT68), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n508_), .A2(new_n510_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT8), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(new_n511_), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n587_), .B(new_n500_), .C1(new_n581_), .C2(new_n580_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT68), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(new_n589_), .A3(new_n579_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n584_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT12), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n471_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n582_), .A2(new_n514_), .ZN(new_n594_));
  AOI22_X1  g393(.A1(new_n518_), .A2(new_n593_), .B1(new_n594_), .B2(new_n592_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n591_), .A2(new_n595_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n499_), .A2(new_n495_), .A3(new_n492_), .ZN(new_n597_));
  AOI22_X1  g396(.A1(new_n586_), .A2(new_n511_), .B1(new_n597_), .B2(new_n490_), .ZN(new_n598_));
  AOI21_X1  g397(.A(KEYINPUT66), .B1(new_n481_), .B2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(new_n594_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n596_), .B1(new_n579_), .B2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(G176gat), .B(G204gat), .Z(new_n602_));
  XNOR2_X1  g401(.A(G120gat), .B(G148gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n601_), .B(new_n607_), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n608_), .A2(KEYINPUT13), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(KEYINPUT13), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n556_), .A2(new_n576_), .A3(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n613_), .A2(new_n438_), .A3(new_n429_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT98), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n613_), .A2(KEYINPUT98), .A3(new_n438_), .A4(new_n429_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT38), .ZN(new_n619_));
  OAI21_X1  g418(.A(KEYINPUT99), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT99), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n616_), .A2(new_n621_), .A3(KEYINPUT38), .A4(new_n617_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n548_), .A2(new_n551_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n436_), .A2(new_n624_), .A3(new_n486_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n612_), .A2(new_n576_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n625_), .A2(KEYINPUT100), .A3(new_n626_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n429_), .B1(new_n630_), .B2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(G1gat), .ZN(new_n634_));
  AOI21_X1  g433(.A(KEYINPUT101), .B1(new_n618_), .B2(new_n619_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n618_), .A2(KEYINPUT101), .A3(new_n619_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n623_), .B(new_n634_), .C1(new_n635_), .C2(new_n636_), .ZN(G1324gat));
  OAI21_X1  g436(.A(G8gat), .B1(new_n627_), .B2(new_n407_), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n638_), .A2(KEYINPUT102), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(KEYINPUT102), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n639_), .A2(KEYINPUT39), .A3(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n613_), .A2(new_n437_), .A3(new_n432_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT39), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n638_), .A2(KEYINPUT102), .A3(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n641_), .A2(new_n642_), .A3(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT40), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(G1325gat));
  INV_X1    g446(.A(G15gat), .ZN(new_n648_));
  INV_X1    g447(.A(new_n428_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n613_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n649_), .B1(new_n630_), .B2(new_n632_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n651_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(KEYINPUT41), .B1(new_n651_), .B2(G15gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n650_), .B1(new_n652_), .B2(new_n653_), .ZN(G1326gat));
  INV_X1    g453(.A(KEYINPUT104), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n399_), .B(KEYINPUT103), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n656_), .B1(new_n629_), .B2(new_n631_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n655_), .B1(new_n658_), .B2(G22gat), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT42), .ZN(new_n660_));
  INV_X1    g459(.A(G22gat), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n657_), .A2(KEYINPUT104), .A3(new_n661_), .ZN(new_n662_));
  OR3_X1    g461(.A1(new_n659_), .A2(new_n660_), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n656_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n613_), .A2(new_n661_), .A3(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n660_), .B1(new_n659_), .B2(new_n662_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n663_), .A2(new_n665_), .A3(new_n666_), .ZN(G1327gat));
  INV_X1    g466(.A(new_n624_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n436_), .A2(new_n668_), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n612_), .A2(new_n576_), .A3(new_n485_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(G29gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(new_n672_), .A3(new_n429_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n411_), .A2(new_n428_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n430_), .A2(new_n435_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n555_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(KEYINPUT43), .B1(new_n676_), .B2(KEYINPUT105), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n678_), .B(new_n679_), .C1(new_n436_), .C2(new_n555_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n677_), .A2(new_n670_), .A3(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT106), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n681_), .A2(KEYINPUT106), .A3(KEYINPUT44), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n403_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n673_), .B1(new_n686_), .B2(new_n672_), .ZN(G1328gat));
  INV_X1    g486(.A(G36gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n671_), .A2(new_n688_), .A3(new_n432_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT45), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n407_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n690_), .B1(new_n691_), .B2(new_n688_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT46), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(G1329gat));
  NAND3_X1  g493(.A1(new_n671_), .A2(new_n414_), .A3(new_n649_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n428_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n696_), .B2(new_n414_), .ZN(new_n697_));
  XOR2_X1   g496(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(G1330gat));
  NAND3_X1  g498(.A1(new_n671_), .A2(new_n520_), .A3(new_n664_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n399_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n700_), .B1(new_n701_), .B2(new_n520_), .ZN(G1331gat));
  INV_X1    g501(.A(new_n576_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n556_), .A2(new_n703_), .A3(new_n611_), .ZN(new_n704_));
  AOI21_X1  g503(.A(G57gat), .B1(new_n704_), .B2(new_n429_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n611_), .A2(new_n703_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n625_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT108), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n707_), .B(new_n708_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n709_), .A2(new_n429_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n705_), .B1(new_n710_), .B2(G57gat), .ZN(G1332gat));
  INV_X1    g510(.A(G64gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n704_), .A2(new_n712_), .A3(new_n432_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT48), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n709_), .A2(new_n432_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n715_), .B2(G64gat), .ZN(new_n716_));
  AOI211_X1 g515(.A(KEYINPUT48), .B(new_n712_), .C1(new_n709_), .C2(new_n432_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n713_), .B1(new_n716_), .B2(new_n717_), .ZN(G1333gat));
  NAND3_X1  g517(.A1(new_n704_), .A2(new_n465_), .A3(new_n649_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT49), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n709_), .A2(new_n649_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n721_), .B2(G71gat), .ZN(new_n722_));
  AOI211_X1 g521(.A(KEYINPUT49), .B(new_n465_), .C1(new_n709_), .C2(new_n649_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n719_), .B1(new_n722_), .B2(new_n723_), .ZN(G1334gat));
  NAND3_X1  g523(.A1(new_n704_), .A2(new_n463_), .A3(new_n664_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT50), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n709_), .A2(new_n664_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n727_), .B2(G78gat), .ZN(new_n728_));
  AOI211_X1 g527(.A(KEYINPUT50), .B(new_n463_), .C1(new_n709_), .C2(new_n664_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(G1335gat));
  NAND2_X1  g529(.A1(new_n706_), .A2(new_n486_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n677_), .A2(new_n680_), .A3(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(G85gat), .B1(new_n733_), .B2(new_n403_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n669_), .A2(new_n732_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n736_), .A2(new_n493_), .A3(new_n429_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n734_), .A2(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT109), .ZN(G1336gat));
  NOR3_X1   g538(.A1(new_n733_), .A2(new_n254_), .A3(new_n407_), .ZN(new_n740_));
  AOI21_X1  g539(.A(G92gat), .B1(new_n736_), .B2(new_n432_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1337gat));
  OAI21_X1  g541(.A(G99gat), .B1(new_n733_), .B2(new_n428_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n736_), .A2(new_n488_), .A3(new_n649_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g545(.A1(new_n736_), .A2(new_n489_), .A3(new_n401_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n677_), .A2(new_n401_), .A3(new_n680_), .A4(new_n732_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n749_), .B(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n748_), .B1(new_n751_), .B2(G106gat), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n749_), .A2(KEYINPUT110), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n749_), .A2(KEYINPUT110), .ZN(new_n754_));
  NOR4_X1   g553(.A1(new_n753_), .A2(new_n754_), .A3(KEYINPUT52), .A4(new_n489_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n747_), .B1(new_n752_), .B2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT53), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT53), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n758_), .B(new_n747_), .C1(new_n752_), .C2(new_n755_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(G1339gat));
  NAND3_X1  g559(.A1(new_n555_), .A2(new_n485_), .A3(new_n576_), .ZN(new_n761_));
  OR3_X1    g560(.A1(new_n761_), .A2(new_n612_), .A3(KEYINPUT54), .ZN(new_n762_));
  OAI21_X1  g561(.A(KEYINPUT54), .B1(new_n761_), .B2(new_n612_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT117), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n561_), .A2(new_n567_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT113), .ZN(new_n767_));
  INV_X1    g566(.A(new_n565_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n561_), .A2(new_n567_), .A3(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n767_), .A2(new_n768_), .A3(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n565_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n559_), .A3(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n573_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT114), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT114), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n773_), .A2(new_n776_), .A3(new_n573_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n601_), .A2(new_n607_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n591_), .A2(new_n595_), .A3(KEYINPUT55), .ZN(new_n781_));
  INV_X1    g580(.A(new_n517_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n516_), .B1(new_n587_), .B2(new_n500_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n593_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n594_), .A2(new_n592_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n784_), .A2(new_n785_), .A3(new_n588_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n578_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n781_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789_));
  AOI211_X1 g588(.A(KEYINPUT68), .B(new_n578_), .C1(new_n481_), .C2(new_n598_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n589_), .B1(new_n588_), .B2(new_n579_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n784_), .A2(new_n785_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n789_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n596_), .A2(KEYINPUT111), .A3(new_n789_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n788_), .A2(new_n796_), .A3(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(KEYINPUT56), .A3(new_n607_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT56), .B1(new_n798_), .B2(new_n607_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n778_), .B(new_n780_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT58), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT116), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n555_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT56), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT111), .B1(new_n596_), .B2(new_n789_), .ZN(new_n807_));
  AOI211_X1 g606(.A(new_n795_), .B(KEYINPUT55), .C1(new_n591_), .C2(new_n595_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n781_), .A2(new_n787_), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n807_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n806_), .B1(new_n810_), .B2(new_n606_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n779_), .B1(new_n811_), .B2(new_n799_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n812_), .A2(new_n813_), .A3(KEYINPUT58), .A4(new_n778_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n804_), .A2(new_n805_), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n811_), .A2(new_n816_), .A3(new_n799_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n779_), .B1(new_n801_), .B2(KEYINPUT112), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n703_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n778_), .A2(new_n608_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n668_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT57), .B1(new_n822_), .B2(KEYINPUT115), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n624_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT115), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n824_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n765_), .B(new_n815_), .C1(new_n823_), .C2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n486_), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n804_), .A2(new_n805_), .A3(new_n814_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n822_), .A2(KEYINPUT115), .A3(KEYINPUT57), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n826_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n830_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n833_), .A2(new_n765_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n764_), .B1(new_n829_), .B2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n435_), .A2(new_n429_), .A3(new_n649_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT59), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n764_), .B1(new_n833_), .B2(new_n485_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n837_), .A3(new_n841_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n839_), .A2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n843_), .A2(G113gat), .A3(new_n703_), .ZN(new_n844_));
  INV_X1    g643(.A(G113gat), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(new_n838_), .B2(new_n576_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n844_), .A2(new_n846_), .ZN(G1340gat));
  NAND3_X1  g646(.A1(new_n839_), .A2(new_n612_), .A3(new_n842_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(KEYINPUT119), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n839_), .A2(new_n850_), .A3(new_n612_), .A4(new_n842_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n849_), .A2(G120gat), .A3(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n838_), .ZN(new_n853_));
  INV_X1    g652(.A(G120gat), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n611_), .B2(KEYINPUT60), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n853_), .B(new_n855_), .C1(KEYINPUT60), .C2(new_n854_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n852_), .A2(new_n856_), .ZN(G1341gat));
  NAND3_X1  g656(.A1(new_n843_), .A2(G127gat), .A3(new_n485_), .ZN(new_n858_));
  INV_X1    g657(.A(G127gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n838_), .B2(new_n486_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n858_), .A2(new_n860_), .ZN(G1342gat));
  AOI21_X1  g660(.A(G134gat), .B1(new_n853_), .B2(new_n624_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT120), .B(G134gat), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n555_), .A2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n862_), .B1(new_n843_), .B2(new_n864_), .ZN(G1343gat));
  INV_X1    g664(.A(new_n764_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n485_), .B1(new_n833_), .B2(new_n765_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n815_), .B1(new_n823_), .B2(new_n827_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(KEYINPUT117), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n866_), .B1(new_n867_), .B2(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n432_), .A2(new_n399_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n428_), .A2(new_n871_), .A3(new_n429_), .ZN(new_n872_));
  OAI21_X1  g671(.A(KEYINPUT121), .B1(new_n870_), .B2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT121), .ZN(new_n874_));
  INV_X1    g673(.A(new_n872_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n835_), .A2(new_n874_), .A3(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n873_), .A2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n703_), .ZN(new_n878_));
  XOR2_X1   g677(.A(KEYINPUT122), .B(G141gat), .Z(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1344gat));
  NAND2_X1  g679(.A1(new_n877_), .A2(new_n612_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g681(.A1(new_n877_), .A2(new_n485_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT61), .B(G155gat), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n883_), .B(new_n884_), .ZN(G1346gat));
  AOI21_X1  g684(.A(G162gat), .B1(new_n877_), .B2(new_n624_), .ZN(new_n886_));
  AOI211_X1 g685(.A(new_n209_), .B(new_n555_), .C1(new_n873_), .C2(new_n876_), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT123), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n555_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n877_), .A2(G162gat), .A3(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT123), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n668_), .B1(new_n873_), .B2(new_n876_), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n890_), .B(new_n891_), .C1(G162gat), .C2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n888_), .A2(new_n893_), .ZN(G1347gat));
  NOR3_X1   g693(.A1(new_n428_), .A2(new_n429_), .A3(new_n407_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n840_), .A2(new_n656_), .A3(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(G169gat), .B1(new_n896_), .B2(new_n576_), .ZN(new_n897_));
  OR2_X1    g696(.A1(new_n897_), .A2(KEYINPUT124), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(KEYINPUT124), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n898_), .A2(KEYINPUT62), .A3(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT125), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n896_), .A2(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n896_), .A2(new_n901_), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n703_), .B(new_n325_), .C1(new_n902_), .C2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT62), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n897_), .A2(KEYINPUT124), .A3(new_n905_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n900_), .A2(new_n904_), .A3(new_n906_), .ZN(G1348gat));
  OAI21_X1  g706(.A(new_n612_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n908_));
  NOR4_X1   g707(.A1(new_n870_), .A2(new_n319_), .A3(new_n611_), .A4(new_n401_), .ZN(new_n909_));
  AOI22_X1  g708(.A1(new_n908_), .A2(new_n279_), .B1(new_n895_), .B2(new_n909_), .ZN(G1349gat));
  NOR2_X1   g709(.A1(new_n902_), .A2(new_n903_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n911_), .A2(new_n486_), .A3(new_n259_), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n835_), .A2(new_n485_), .A3(new_n399_), .A4(new_n895_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(new_n273_), .B2(new_n913_), .ZN(G1350gat));
  OAI21_X1  g713(.A(G190gat), .B1(new_n911_), .B2(new_n555_), .ZN(new_n915_));
  OR2_X1    g714(.A1(new_n668_), .A2(new_n323_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n911_), .B2(new_n916_), .ZN(G1351gat));
  NOR2_X1   g716(.A1(new_n429_), .A2(new_n407_), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n835_), .A2(new_n428_), .A3(new_n401_), .A4(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n919_), .A2(new_n576_), .ZN(new_n920_));
  XOR2_X1   g719(.A(KEYINPUT126), .B(G197gat), .Z(new_n921_));
  XNOR2_X1  g720(.A(new_n920_), .B(new_n921_), .ZN(G1352gat));
  NOR2_X1   g721(.A1(new_n919_), .A2(new_n611_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n923_), .B1(KEYINPUT127), .B2(new_n293_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(KEYINPUT127), .B(G204gat), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n923_), .B2(new_n925_), .ZN(G1353gat));
  NOR2_X1   g725(.A1(new_n919_), .A2(new_n486_), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n927_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n928_));
  XOR2_X1   g727(.A(KEYINPUT63), .B(G211gat), .Z(new_n929_));
  AOI21_X1  g728(.A(new_n928_), .B1(new_n927_), .B2(new_n929_), .ZN(G1354gat));
  INV_X1    g729(.A(G218gat), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n919_), .A2(new_n931_), .A3(new_n555_), .ZN(new_n932_));
  OR2_X1    g731(.A1(new_n919_), .A2(new_n668_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n932_), .B1(new_n931_), .B2(new_n933_), .ZN(G1355gat));
endmodule


