//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n567_, new_n568_, new_n569_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n610_,
    new_n611_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n634_, new_n635_, new_n636_, new_n637_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n791_, new_n792_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n804_, new_n805_, new_n806_, new_n807_, new_n809_,
    new_n810_, new_n811_, new_n813_, new_n814_, new_n815_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(G141gat), .B(G148gat), .Z(new_n203_));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT1), .ZN(new_n205_));
  OR2_X1    g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n204_), .A2(KEYINPUT1), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n203_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT85), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  XOR2_X1   g010(.A(new_n211_), .B(KEYINPUT3), .Z(new_n212_));
  NAND2_X1  g011(.A1(G141gat), .A2(G148gat), .ZN(new_n213_));
  XOR2_X1   g012(.A(new_n213_), .B(KEYINPUT2), .Z(new_n214_));
  OAI211_X1 g013(.A(new_n204_), .B(new_n206_), .C1(new_n212_), .C2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n210_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G127gat), .B(G134gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT84), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G113gat), .B(G120gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n218_), .B(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n216_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT90), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n216_), .A2(new_n220_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT4), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT91), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n221_), .A2(KEYINPUT4), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G225gat), .A2(G233gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n226_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT92), .ZN(new_n231_));
  AOI22_X1  g030(.A1(new_n230_), .A2(new_n231_), .B1(new_n224_), .B2(new_n228_), .ZN(new_n232_));
  XOR2_X1   g031(.A(G57gat), .B(G85gat), .Z(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT94), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(G1gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n236_));
  INV_X1    g035(.A(G29gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(new_n235_), .B(new_n238_), .Z(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n226_), .A2(new_n229_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT92), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n232_), .A2(new_n240_), .A3(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT33), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n232_), .A2(KEYINPUT33), .A3(new_n240_), .A4(new_n242_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n228_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n240_), .B1(new_n224_), .B2(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(new_n248_), .B(KEYINPUT95), .Z(new_n249_));
  NOR2_X1   g048(.A1(new_n227_), .A2(new_n247_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n249_), .B1(new_n226_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT20), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT25), .B(G183gat), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n253_), .B(KEYINPUT87), .Z(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT26), .B(G190gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(G169gat), .ZN(new_n257_));
  INV_X1    g056(.A(G176gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n259_), .A2(KEYINPUT24), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G169gat), .A2(G176gat), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n259_), .A2(KEYINPUT24), .A3(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G183gat), .A2(G190gat), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n264_), .A2(KEYINPUT23), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n263_), .B(KEYINPUT80), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n265_), .B1(new_n266_), .B2(KEYINPUT23), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n256_), .A2(new_n260_), .A3(new_n262_), .A4(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT88), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT22), .B(G169gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n258_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT23), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n264_), .A2(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n274_), .B1(new_n266_), .B2(new_n273_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(G183gat), .A2(G190gat), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n261_), .B(new_n272_), .C1(new_n275_), .C2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n270_), .A2(new_n277_), .ZN(new_n278_));
  XOR2_X1   g077(.A(G197gat), .B(G204gat), .Z(new_n279_));
  OR2_X1    g078(.A1(new_n279_), .A2(KEYINPUT21), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(KEYINPUT21), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G211gat), .B(G218gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n281_), .A2(new_n282_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n252_), .B1(new_n278_), .B2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n267_), .B1(G183gat), .B2(G190gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT81), .ZN(new_n288_));
  AOI22_X1  g087(.A1(new_n272_), .A2(new_n288_), .B1(G169gat), .B2(G176gat), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n287_), .B(new_n289_), .C1(new_n288_), .C2(new_n272_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n275_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(new_n260_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n255_), .A2(new_n253_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n262_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT79), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n290_), .B1(new_n292_), .B2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT82), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n286_), .B1(new_n285_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G226gat), .A2(G233gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT19), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n285_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n285_), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n302_), .A2(new_n277_), .ZN(new_n303_));
  AOI211_X1 g102(.A(new_n252_), .B(new_n300_), .C1(new_n270_), .C2(new_n303_), .ZN(new_n304_));
  AOI22_X1  g103(.A1(new_n298_), .A2(new_n300_), .B1(new_n301_), .B2(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(G8gat), .B(G36gat), .Z(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G64gat), .B(G92gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n305_), .B(new_n310_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n251_), .A2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n245_), .A2(new_n246_), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT96), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n302_), .B1(new_n216_), .B2(KEYINPUT29), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G228gat), .A2(G233gat), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n316_), .B(new_n317_), .Z(new_n318_));
  XOR2_X1   g117(.A(G78gat), .B(G106gat), .Z(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT86), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n216_), .A2(KEYINPUT29), .ZN(new_n322_));
  XOR2_X1   g121(.A(G22gat), .B(G50gat), .Z(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT28), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n322_), .B(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n321_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n318_), .B(new_n319_), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n326_), .B(new_n327_), .Z(new_n328_));
  NAND2_X1  g127(.A1(new_n232_), .A2(new_n242_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n239_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n243_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n310_), .A2(KEYINPUT32), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n305_), .A2(KEYINPUT97), .A3(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n298_), .A2(new_n300_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT98), .B(KEYINPUT20), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n335_), .B1(new_n303_), .B2(new_n268_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n301_), .A2(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n334_), .B1(new_n300_), .B2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT97), .B1(new_n338_), .B2(new_n332_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n305_), .A2(new_n332_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n333_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n328_), .B1(new_n331_), .B2(new_n341_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n245_), .A2(KEYINPUT96), .A3(new_n246_), .A4(new_n312_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n315_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(G71gat), .B(G99gat), .Z(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT83), .B(G43gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n345_), .B(new_n346_), .Z(new_n347_));
  XNOR2_X1  g146(.A(new_n297_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(new_n220_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G227gat), .A2(G233gat), .ZN(new_n350_));
  INV_X1    g149(.A(G15gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT30), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT31), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n349_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n349_), .A2(new_n355_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT27), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n311_), .A2(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n360_), .B1(new_n305_), .B2(new_n310_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n362_), .B1(new_n310_), .B2(new_n338_), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n330_), .A2(new_n243_), .A3(new_n361_), .A4(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n359_), .B1(new_n364_), .B2(new_n328_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n344_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n331_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n361_), .A2(new_n363_), .ZN(new_n368_));
  NOR3_X1   g167(.A1(new_n368_), .A2(new_n328_), .A3(new_n358_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n366_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT66), .ZN(new_n372_));
  INV_X1    g171(.A(G99gat), .ZN(new_n373_));
  INV_X1    g172(.A(G106gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT65), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT7), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT7), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT65), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n375_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  AOI22_X1  g179(.A1(new_n373_), .A2(new_n374_), .B1(new_n378_), .B2(KEYINPUT65), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n372_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G99gat), .A2(G106gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT6), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n375_), .A2(new_n379_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT65), .B(KEYINPUT7), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n385_), .B(KEYINPUT66), .C1(new_n386_), .C2(new_n375_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n382_), .A2(new_n384_), .A3(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(G85gat), .B(G92gat), .Z(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT8), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n388_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n389_), .A2(KEYINPUT9), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT9), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n394_), .A2(G85gat), .A3(G92gat), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n384_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT10), .B(G99gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT64), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n393_), .B(new_n396_), .C1(new_n398_), .C2(G106gat), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n385_), .B1(new_n386_), .B2(new_n375_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT6), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n383_), .B(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n389_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT8), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n392_), .A2(new_n399_), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G29gat), .B(G36gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT71), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G43gat), .B(G50gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT35), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G232gat), .A2(G233gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT34), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  AOI22_X1  g214(.A1(new_n407_), .A2(new_n411_), .B1(new_n412_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT68), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n402_), .B1(new_n400_), .B2(new_n372_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n390_), .B1(new_n418_), .B2(new_n387_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n384_), .B(new_n385_), .C1(new_n375_), .C2(new_n386_), .ZN(new_n420_));
  AOI21_X1  g219(.A(KEYINPUT8), .B1(new_n420_), .B2(new_n389_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n417_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n392_), .A2(KEYINPUT68), .A3(new_n405_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(KEYINPUT69), .B1(new_n424_), .B2(new_n399_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT69), .ZN(new_n426_));
  INV_X1    g225(.A(new_n399_), .ZN(new_n427_));
  AOI211_X1 g226(.A(new_n426_), .B(new_n427_), .C1(new_n422_), .C2(new_n423_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n425_), .A2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n411_), .B(KEYINPUT15), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n416_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n415_), .A2(new_n412_), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n433_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G190gat), .B(G218gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT72), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT73), .ZN(new_n439_));
  XOR2_X1   g238(.A(G134gat), .B(G162gat), .Z(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(new_n441_), .B(KEYINPUT36), .Z(new_n442_));
  AND2_X1   g241(.A1(new_n436_), .A2(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n441_), .A2(KEYINPUT36), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT74), .B1(new_n436_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT74), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n434_), .A2(new_n447_), .A3(new_n444_), .A4(new_n435_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n443_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(KEYINPUT76), .B(G8gat), .Z(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT14), .B1(new_n451_), .B2(new_n202_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G15gat), .B(G22gat), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G1gat), .B(G8gat), .ZN(new_n455_));
  XOR2_X1   g254(.A(new_n454_), .B(new_n455_), .Z(new_n456_));
  NAND2_X1  g255(.A1(G231gat), .A2(G233gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G57gat), .B(G64gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT11), .ZN(new_n460_));
  XOR2_X1   g259(.A(G71gat), .B(G78gat), .Z(new_n461_));
  OR2_X1    g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n459_), .A2(KEYINPUT11), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n460_), .A2(new_n461_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n462_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n458_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT17), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G127gat), .B(G155gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G183gat), .B(G211gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  NOR3_X1   g271(.A1(new_n466_), .A2(new_n467_), .A3(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n473_), .B1(new_n458_), .B2(new_n465_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n472_), .B(new_n467_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n465_), .A2(KEYINPUT67), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT67), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n462_), .B(new_n477_), .C1(new_n463_), .C2(new_n464_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n475_), .B1(new_n458_), .B2(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n480_), .B1(new_n458_), .B2(new_n479_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n474_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n371_), .A2(new_n450_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT12), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n465_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n487_), .B1(new_n425_), .B2(new_n428_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n479_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n485_), .B1(new_n489_), .B2(new_n407_), .ZN(new_n490_));
  INV_X1    g289(.A(G230gat), .ZN(new_n491_));
  INV_X1    g290(.A(G233gat), .ZN(new_n492_));
  OAI22_X1  g291(.A1(new_n479_), .A2(new_n406_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT70), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT70), .ZN(new_n495_));
  OAI221_X1 g294(.A(new_n495_), .B1(new_n491_), .B2(new_n492_), .C1(new_n479_), .C2(new_n406_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n488_), .A2(new_n490_), .A3(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n491_), .A2(new_n492_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n489_), .A2(new_n407_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n489_), .A2(new_n407_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n499_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n498_), .A2(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(G120gat), .B(G148gat), .Z(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT5), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G176gat), .B(G204gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n504_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n504_), .A2(new_n508_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT13), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n509_), .A2(KEYINPUT13), .A3(new_n510_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n430_), .A2(new_n456_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT78), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G229gat), .A2(G233gat), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n456_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n520_), .B1(new_n521_), .B2(new_n411_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n411_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n456_), .B(new_n523_), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n518_), .A2(new_n522_), .B1(new_n524_), .B2(new_n520_), .ZN(new_n525_));
  XOR2_X1   g324(.A(G113gat), .B(G141gat), .Z(new_n526_));
  XNOR2_X1  g325(.A(G169gat), .B(G197gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n525_), .B(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n515_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n484_), .A2(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n202_), .B1(new_n533_), .B2(new_n331_), .ZN(new_n534_));
  AOI22_X1  g333(.A1(new_n344_), .A2(new_n365_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n535_), .A2(new_n530_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n536_), .A2(KEYINPUT99), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n536_), .A2(KEYINPUT99), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  AOI211_X1 g338(.A(KEYINPUT37), .B(new_n443_), .C1(new_n446_), .C2(new_n448_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT37), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n446_), .A2(new_n448_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n442_), .B(KEYINPUT75), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n436_), .A2(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n541_), .B1(new_n542_), .B2(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n540_), .A2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n546_), .A2(new_n482_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n515_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n539_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n551_), .A2(new_n202_), .A3(new_n331_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n534_), .B1(new_n553_), .B2(KEYINPUT38), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT38), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n552_), .A2(KEYINPUT100), .A3(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(KEYINPUT100), .B1(new_n552_), .B2(new_n555_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n554_), .B1(new_n556_), .B2(new_n557_), .ZN(G1324gat));
  NAND2_X1  g357(.A1(new_n533_), .A2(new_n368_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(G8gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT39), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n551_), .A2(new_n451_), .A3(new_n368_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n563_), .B(new_n565_), .ZN(G1325gat));
  NAND3_X1  g365(.A1(new_n551_), .A2(new_n351_), .A3(new_n359_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n351_), .B1(new_n533_), .B2(new_n359_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT41), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(G1326gat));
  INV_X1    g369(.A(G22gat), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n571_), .B1(new_n533_), .B2(new_n328_), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n572_), .B(KEYINPUT42), .Z(new_n573_));
  NAND3_X1  g372(.A1(new_n551_), .A2(new_n571_), .A3(new_n328_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(G1327gat));
  NAND2_X1  g374(.A1(new_n449_), .A2(new_n482_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n576_), .A2(new_n515_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n539_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(G29gat), .B1(new_n579_), .B2(new_n331_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n546_), .ZN(new_n581_));
  OAI21_X1  g380(.A(KEYINPUT43), .B1(new_n581_), .B2(KEYINPUT102), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n371_), .A2(new_n582_), .A3(new_n546_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n582_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n584_), .B1(new_n535_), .B2(new_n581_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n483_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(new_n531_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT44), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n586_), .A2(KEYINPUT44), .A3(new_n531_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n367_), .A2(new_n237_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n580_), .B1(new_n591_), .B2(new_n592_), .ZN(G1328gat));
  NAND3_X1  g392(.A1(new_n589_), .A2(new_n368_), .A3(new_n590_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(G36gat), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n368_), .B(KEYINPUT103), .Z(new_n596_));
  NOR2_X1   g395(.A1(new_n596_), .A2(G36gat), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n577_), .B(new_n597_), .C1(new_n537_), .C2(new_n538_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT45), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n595_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT46), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(G1329gat));
  NAND3_X1  g401(.A1(new_n591_), .A2(G43gat), .A3(new_n359_), .ZN(new_n603_));
  INV_X1    g402(.A(G43gat), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n604_), .B1(new_n578_), .B2(new_n358_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n603_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n606_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(G1330gat));
  AOI21_X1  g408(.A(G50gat), .B1(new_n579_), .B2(new_n328_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n328_), .A2(G50gat), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n610_), .B1(new_n591_), .B2(new_n611_), .ZN(G1331gat));
  AND4_X1   g411(.A1(new_n530_), .A2(new_n371_), .A3(new_n547_), .A4(new_n515_), .ZN(new_n613_));
  INV_X1    g412(.A(G57gat), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n613_), .A2(new_n614_), .A3(new_n331_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n548_), .A2(new_n529_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NOR3_X1   g416(.A1(new_n484_), .A2(new_n367_), .A3(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n615_), .B1(new_n618_), .B2(new_n614_), .ZN(G1332gat));
  NOR2_X1   g418(.A1(new_n484_), .A2(new_n617_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(G64gat), .B1(new_n621_), .B2(new_n596_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT48), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n596_), .A2(G64gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT105), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n613_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n623_), .A2(new_n626_), .ZN(G1333gat));
  INV_X1    g426(.A(G71gat), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n628_), .B1(new_n620_), .B2(new_n359_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(KEYINPUT106), .B(KEYINPUT49), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n613_), .A2(new_n628_), .A3(new_n359_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(G1334gat));
  INV_X1    g432(.A(G78gat), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n634_), .B1(new_n620_), .B2(new_n328_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT50), .Z(new_n636_));
  NAND3_X1  g435(.A1(new_n613_), .A2(new_n634_), .A3(new_n328_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(G1335gat));
  NOR4_X1   g437(.A1(new_n535_), .A2(new_n529_), .A3(new_n548_), .A4(new_n576_), .ZN(new_n639_));
  AOI21_X1  g438(.A(G85gat), .B1(new_n639_), .B2(new_n331_), .ZN(new_n640_));
  AOI211_X1 g439(.A(new_n483_), .B(new_n617_), .C1(new_n583_), .C2(new_n585_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n331_), .A2(G85gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT107), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n640_), .B1(new_n641_), .B2(new_n643_), .ZN(G1336gat));
  INV_X1    g443(.A(new_n641_), .ZN(new_n645_));
  OAI21_X1  g444(.A(G92gat), .B1(new_n645_), .B2(new_n596_), .ZN(new_n646_));
  INV_X1    g445(.A(G92gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n639_), .A2(new_n647_), .A3(new_n368_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(G1337gat));
  OAI21_X1  g448(.A(G99gat), .B1(new_n645_), .B2(new_n358_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n398_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n639_), .A2(new_n359_), .A3(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(KEYINPUT108), .B(KEYINPUT51), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(G1338gat));
  NAND3_X1  g454(.A1(new_n586_), .A2(new_n328_), .A3(new_n616_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT109), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n641_), .A2(KEYINPUT109), .A3(new_n328_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n658_), .A2(new_n659_), .A3(G106gat), .ZN(new_n660_));
  NOR2_X1   g459(.A1(KEYINPUT110), .A2(KEYINPUT52), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  XOR2_X1   g461(.A(KEYINPUT110), .B(KEYINPUT52), .Z(new_n663_));
  NAND4_X1  g462(.A1(new_n658_), .A2(new_n659_), .A3(G106gat), .A4(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n639_), .A2(new_n374_), .A3(new_n328_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n662_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT53), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT53), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n662_), .A2(new_n668_), .A3(new_n664_), .A4(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(G1339gat));
  NAND2_X1  g469(.A1(new_n369_), .A2(new_n331_), .ZN(new_n671_));
  OAI211_X1 g470(.A(new_n518_), .B(new_n520_), .C1(new_n523_), .C2(new_n456_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n528_), .B1(new_n524_), .B2(new_n519_), .ZN(new_n673_));
  AOI22_X1  g472(.A1(new_n672_), .A2(new_n673_), .B1(new_n525_), .B2(new_n528_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n511_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n529_), .A2(new_n509_), .ZN(new_n676_));
  XOR2_X1   g475(.A(KEYINPUT111), .B(KEYINPUT55), .Z(new_n677_));
  NAND2_X1  g476(.A1(new_n498_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT112), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT112), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n498_), .A2(new_n680_), .A3(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n488_), .A2(new_n500_), .A3(new_n490_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(new_n499_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n498_), .ZN(new_n685_));
  AOI22_X1  g484(.A1(new_n684_), .A2(KEYINPUT113), .B1(new_n685_), .B2(KEYINPUT55), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT113), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n683_), .A2(new_n687_), .A3(new_n499_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n682_), .A2(new_n686_), .A3(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT56), .B1(new_n689_), .B2(new_n508_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n676_), .B1(new_n690_), .B2(KEYINPUT114), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n684_), .A2(KEYINPUT113), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n685_), .A2(KEYINPUT55), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(new_n688_), .A3(new_n693_), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n498_), .A2(new_n680_), .A3(new_n677_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n680_), .B1(new_n498_), .B2(new_n677_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n508_), .B1(new_n694_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT56), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT114), .ZN(new_n701_));
  OAI211_X1 g500(.A(KEYINPUT56), .B(new_n508_), .C1(new_n694_), .C2(new_n697_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n700_), .A2(new_n701_), .A3(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n675_), .B1(new_n691_), .B2(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n704_), .A2(new_n449_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT57), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT117), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT58), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n674_), .A2(new_n509_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n700_), .B2(new_n702_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n708_), .B1(new_n710_), .B2(KEYINPUT116), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT116), .ZN(new_n712_));
  AOI211_X1 g511(.A(new_n712_), .B(new_n709_), .C1(new_n700_), .C2(new_n702_), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n707_), .B(new_n546_), .C1(new_n711_), .C2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n710_), .A2(KEYINPUT58), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n709_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n702_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n717_), .B1(new_n718_), .B2(new_n690_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n712_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n710_), .A2(KEYINPUT116), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n720_), .A2(new_n721_), .A3(new_n708_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n707_), .B1(new_n722_), .B2(new_n546_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n706_), .B1(new_n716_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT57), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n725_), .B1(new_n704_), .B2(new_n449_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT115), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT115), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n728_), .B(new_n725_), .C1(new_n704_), .C2(new_n449_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(KEYINPUT118), .B1(new_n724_), .B2(new_n730_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n727_), .A2(new_n729_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n546_), .B1(new_n711_), .B2(new_n713_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT117), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(new_n715_), .A3(new_n714_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT118), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n732_), .A2(new_n735_), .A3(new_n736_), .A4(new_n706_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n731_), .A2(new_n482_), .A3(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n549_), .A2(new_n529_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT54), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n739_), .B(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n671_), .B1(new_n738_), .B2(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(G113gat), .B1(new_n742_), .B2(new_n529_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT119), .ZN(new_n744_));
  INV_X1    g543(.A(new_n742_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n726_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n482_), .B1(new_n724_), .B2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(new_n741_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n671_), .A2(KEYINPUT59), .ZN(new_n749_));
  AOI22_X1  g548(.A1(new_n745_), .A2(KEYINPUT59), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n529_), .A2(G113gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n744_), .B1(new_n750_), .B2(new_n751_), .ZN(G1340gat));
  AOI21_X1  g551(.A(new_n548_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT59), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n753_), .B1(new_n742_), .B2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT120), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT120), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n757_), .B(new_n753_), .C1(new_n742_), .C2(new_n754_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n756_), .A2(G120gat), .A3(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(G120gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n760_), .B1(new_n548_), .B2(KEYINPUT60), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n742_), .B(new_n761_), .C1(KEYINPUT60), .C2(new_n760_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n759_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT121), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n759_), .A2(KEYINPUT121), .A3(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(G1341gat));
  INV_X1    g566(.A(G127gat), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n742_), .A2(new_n768_), .A3(new_n483_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n750_), .A2(new_n483_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n769_), .B1(new_n771_), .B2(new_n768_), .ZN(G1342gat));
  INV_X1    g571(.A(G134gat), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n742_), .A2(new_n773_), .A3(new_n449_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n750_), .A2(new_n546_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n774_), .B1(new_n776_), .B2(new_n773_), .ZN(G1343gat));
  AND2_X1   g576(.A1(new_n358_), .A2(new_n328_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n779_), .B1(new_n738_), .B2(new_n741_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n780_), .A2(new_n331_), .A3(new_n596_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n781_), .A2(new_n530_), .ZN(new_n782_));
  XOR2_X1   g581(.A(KEYINPUT122), .B(G141gat), .Z(new_n783_));
  XNOR2_X1  g582(.A(new_n782_), .B(new_n783_), .ZN(G1344gat));
  NOR2_X1   g583(.A1(new_n781_), .A2(new_n548_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(KEYINPUT123), .B(G148gat), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n785_), .B(new_n786_), .ZN(G1345gat));
  NOR2_X1   g586(.A1(new_n781_), .A2(new_n482_), .ZN(new_n788_));
  XOR2_X1   g587(.A(KEYINPUT61), .B(G155gat), .Z(new_n789_));
  XNOR2_X1  g588(.A(new_n788_), .B(new_n789_), .ZN(G1346gat));
  OAI21_X1  g589(.A(G162gat), .B1(new_n781_), .B2(new_n581_), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n450_), .A2(G162gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n791_), .B1(new_n781_), .B2(new_n792_), .ZN(G1347gat));
  AOI21_X1  g592(.A(new_n328_), .B1(new_n747_), .B2(new_n741_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n596_), .A2(new_n331_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n796_), .A2(new_n358_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n794_), .A2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n257_), .B1(new_n798_), .B2(new_n529_), .ZN(new_n799_));
  OR2_X1    g598(.A1(new_n799_), .A2(KEYINPUT62), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n798_), .A2(new_n529_), .A3(new_n271_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(KEYINPUT62), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n800_), .A2(new_n801_), .A3(new_n802_), .ZN(G1348gat));
  AOI21_X1  g602(.A(G176gat), .B1(new_n798_), .B2(new_n515_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n328_), .B1(new_n738_), .B2(new_n741_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n797_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n806_), .A2(new_n258_), .A3(new_n548_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n804_), .B1(new_n805_), .B2(new_n807_), .ZN(G1349gat));
  NOR2_X1   g607(.A1(new_n806_), .A2(new_n482_), .ZN(new_n809_));
  AOI21_X1  g608(.A(G183gat), .B1(new_n805_), .B2(new_n809_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n806_), .A2(new_n254_), .A3(new_n482_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n810_), .B1(new_n794_), .B2(new_n811_), .ZN(G1350gat));
  NAND3_X1  g611(.A1(new_n798_), .A2(new_n255_), .A3(new_n449_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n798_), .A2(new_n546_), .ZN(new_n814_));
  INV_X1    g613(.A(G190gat), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n813_), .B1(new_n814_), .B2(new_n815_), .ZN(G1351gat));
  NAND2_X1  g615(.A1(new_n780_), .A2(new_n795_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT124), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n780_), .A2(KEYINPUT124), .A3(new_n795_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n530_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT126), .B1(new_n821_), .B2(G197gat), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT126), .ZN(new_n823_));
  INV_X1    g622(.A(G197gat), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n780_), .A2(KEYINPUT124), .A3(new_n795_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT124), .B1(new_n780_), .B2(new_n795_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n823_), .B(new_n824_), .C1(new_n827_), .C2(new_n530_), .ZN(new_n828_));
  OAI211_X1 g627(.A(G197gat), .B(new_n529_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT125), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n819_), .A2(new_n820_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT125), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n831_), .A2(new_n832_), .A3(G197gat), .A4(new_n529_), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n822_), .A2(new_n828_), .B1(new_n830_), .B2(new_n833_), .ZN(G1352gat));
  INV_X1    g633(.A(KEYINPUT127), .ZN(new_n835_));
  AOI211_X1 g634(.A(new_n835_), .B(G204gat), .C1(new_n831_), .C2(new_n515_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n835_), .A2(G204gat), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n835_), .A2(G204gat), .ZN(new_n838_));
  NOR4_X1   g637(.A1(new_n827_), .A2(new_n548_), .A3(new_n837_), .A4(new_n838_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n836_), .A2(new_n839_), .ZN(G1353gat));
  OR2_X1    g639(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n841_));
  NAND2_X1  g640(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n842_));
  AND4_X1   g641(.A1(new_n483_), .A2(new_n831_), .A3(new_n841_), .A4(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n841_), .B1(new_n831_), .B2(new_n483_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(G1354gat));
  OR3_X1    g644(.A1(new_n827_), .A2(G218gat), .A3(new_n450_), .ZN(new_n846_));
  OAI21_X1  g645(.A(G218gat), .B1(new_n827_), .B2(new_n581_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(G1355gat));
endmodule


