//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 0 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n865_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(G190gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT81), .B(G183gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT25), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n207_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT24), .ZN(new_n214_));
  INV_X1    g013(.A(G169gat), .ZN(new_n215_));
  INV_X1    g014(.A(G176gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  MUX2_X1   g016(.A(KEYINPUT24), .B(new_n214_), .S(new_n217_), .Z(new_n218_));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT23), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n212_), .A2(new_n218_), .A3(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G190gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n208_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n219_), .B(KEYINPUT23), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT82), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n226_), .B1(new_n215_), .B2(KEYINPUT22), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT83), .B(G176gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT22), .B(G169gat), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n227_), .B(new_n228_), .C1(new_n229_), .C2(new_n226_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n225_), .A2(new_n230_), .A3(new_n213_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n221_), .A2(new_n231_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n232_), .A2(KEYINPUT84), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n232_), .A2(KEYINPUT84), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(G197gat), .B(G204gat), .Z(new_n236_));
  OR2_X1    g035(.A1(new_n236_), .A2(KEYINPUT21), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(KEYINPUT21), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G211gat), .B(G218gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n238_), .A2(new_n239_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n235_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT94), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(new_n245_), .A3(KEYINPUT20), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT25), .B(G183gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n207_), .A2(new_n247_), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n218_), .A2(new_n220_), .A3(new_n248_), .ZN(new_n249_));
  AOI22_X1  g048(.A1(new_n229_), .A2(new_n228_), .B1(G169gat), .B2(G176gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT95), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n224_), .B1(G183gat), .B2(G190gat), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n249_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n253_), .A2(new_n243_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n246_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G226gat), .A2(G233gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n245_), .B1(new_n244_), .B2(KEYINPUT20), .ZN(new_n259_));
  NOR3_X1   g058(.A1(new_n255_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n258_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n242_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT96), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT20), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n265_), .B1(new_n253_), .B2(new_n243_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n261_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n206_), .B1(new_n260_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT100), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT100), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n270_), .B(new_n206_), .C1(new_n260_), .C2(new_n267_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n258_), .B1(new_n255_), .B2(new_n259_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n264_), .A2(new_n261_), .A3(new_n266_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(new_n205_), .A3(new_n274_), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n275_), .A2(KEYINPUT27), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n273_), .A2(new_n274_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n206_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(new_n275_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT27), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n272_), .A2(new_n276_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(KEYINPUT90), .A2(KEYINPUT3), .ZN(new_n282_));
  INV_X1    g081(.A(G141gat), .ZN(new_n283_));
  INV_X1    g082(.A(G148gat), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT2), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n286_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n287_));
  OAI22_X1  g086(.A1(KEYINPUT90), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n285_), .A2(new_n287_), .A3(new_n288_), .A4(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT88), .ZN(new_n292_));
  XOR2_X1   g091(.A(G141gat), .B(G148gat), .Z(new_n293_));
  AOI22_X1  g092(.A1(new_n290_), .A2(new_n292_), .B1(KEYINPUT1), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G155gat), .A2(G162gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT89), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n298_), .B1(new_n295_), .B2(KEYINPUT1), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n292_), .A2(new_n299_), .ZN(new_n300_));
  NOR3_X1   g099(.A1(new_n295_), .A2(new_n298_), .A3(KEYINPUT1), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n293_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G127gat), .B(G134gat), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  XOR2_X1   g103(.A(G113gat), .B(G120gat), .Z(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n297_), .A2(new_n302_), .A3(new_n306_), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n307_), .A2(KEYINPUT97), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G225gat), .A2(G233gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(KEYINPUT97), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n297_), .A2(new_n302_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT86), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n312_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n313_), .B1(new_n306_), .B2(new_n312_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n308_), .A2(new_n309_), .A3(new_n310_), .A4(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(KEYINPUT4), .B1(new_n311_), .B2(new_n314_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n308_), .A2(new_n310_), .A3(new_n315_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n317_), .B1(new_n318_), .B2(KEYINPUT4), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n309_), .B(KEYINPUT98), .Z(new_n320_));
  OAI21_X1  g119(.A(new_n316_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G1gat), .B(G29gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(G85gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT0), .B(G57gat), .ZN(new_n324_));
  XOR2_X1   g123(.A(new_n323_), .B(new_n324_), .Z(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n321_), .A2(new_n326_), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n316_), .B(new_n325_), .C1(new_n319_), .C2(new_n320_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n311_), .A2(KEYINPUT29), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n242_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(G78gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G228gat), .A2(G233gat), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT91), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n333_), .B1(new_n242_), .B2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(G106gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n332_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(G78gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n331_), .B(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n336_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n337_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT92), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G22gat), .B(G50gat), .ZN(new_n344_));
  OR3_X1    g143(.A1(new_n311_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT28), .B1(new_n311_), .B2(KEYINPUT29), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n344_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n345_), .A2(new_n346_), .A3(new_n344_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n343_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n348_), .A2(new_n343_), .A3(new_n349_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n342_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n350_), .A2(new_n337_), .A3(new_n341_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G71gat), .B(G99gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT85), .B(G43gat), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n356_), .B(new_n357_), .Z(new_n358_));
  NAND2_X1  g157(.A1(G227gat), .A2(G233gat), .ZN(new_n359_));
  INV_X1    g158(.A(G15gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT30), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n235_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n235_), .A2(new_n363_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n358_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n366_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n358_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n369_), .A3(new_n364_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n367_), .A2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n314_), .B(KEYINPUT31), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT87), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT87), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n367_), .A2(new_n370_), .A3(new_n375_), .A4(new_n372_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n355_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n374_), .A2(new_n376_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n329_), .B1(new_n378_), .B2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n326_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n319_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n382_), .B1(new_n383_), .B2(new_n309_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT33), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n328_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  OR2_X1    g185(.A1(new_n328_), .A2(new_n385_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n278_), .A2(new_n386_), .A3(new_n275_), .A4(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n389_));
  NOR3_X1   g188(.A1(new_n260_), .A2(new_n267_), .A3(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n273_), .A2(KEYINPUT99), .A3(new_n274_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT99), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n273_), .A2(new_n392_), .A3(new_n274_), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n390_), .A2(new_n391_), .B1(new_n389_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n329_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n388_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n355_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n397_), .A2(new_n377_), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n281_), .A2(new_n381_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT8), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NOR3_X1   g201(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT6), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT64), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT64), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT6), .ZN(new_n408_));
  AND2_X1   g207(.A1(G99gat), .A2(G106gat), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n406_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n409_), .B1(new_n406_), .B2(new_n408_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n404_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  XOR2_X1   g211(.A(G85gat), .B(G92gat), .Z(new_n413_));
  AOI21_X1  g212(.A(new_n400_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT65), .ZN(new_n415_));
  NOR3_X1   g214(.A1(new_n410_), .A2(new_n411_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G99gat), .A2(G106gat), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n407_), .A2(KEYINPUT6), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n405_), .A2(KEYINPUT64), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n417_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n406_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n421_));
  AOI21_X1  g220(.A(KEYINPUT65), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n404_), .B1(new_n416_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n413_), .A2(new_n400_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n414_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  XOR2_X1   g225(.A(KEYINPUT10), .B(G99gat), .Z(new_n427_));
  INV_X1    g226(.A(G106gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n413_), .A2(KEYINPUT9), .ZN(new_n430_));
  INV_X1    g229(.A(G85gat), .ZN(new_n431_));
  INV_X1    g230(.A(G92gat), .ZN(new_n432_));
  OR3_X1    g231(.A1(new_n431_), .A2(new_n432_), .A3(KEYINPUT9), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n429_), .A2(new_n430_), .A3(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n415_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n420_), .A2(KEYINPUT65), .A3(new_n421_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n434_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT66), .B1(new_n426_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT66), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n424_), .B1(new_n437_), .B2(new_n404_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n441_), .B(new_n438_), .C1(new_n442_), .C2(new_n414_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G57gat), .B(G64gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT11), .ZN(new_n445_));
  XOR2_X1   g244(.A(G71gat), .B(G78gat), .Z(new_n446_));
  OR2_X1    g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n446_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n444_), .A2(KEYINPUT11), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n447_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT12), .ZN(new_n451_));
  OR2_X1    g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n440_), .A2(new_n443_), .A3(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT67), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n426_), .A2(new_n439_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n451_), .B1(new_n457_), .B2(new_n450_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n440_), .A2(KEYINPUT67), .A3(new_n443_), .A4(new_n453_), .ZN(new_n459_));
  AND2_X1   g258(.A1(G230gat), .A2(G233gat), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n460_), .B1(new_n457_), .B2(new_n450_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n456_), .A2(new_n458_), .A3(new_n459_), .A4(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n457_), .A2(new_n450_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n457_), .A2(new_n450_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n460_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G120gat), .B(G148gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT5), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G176gat), .B(G204gat), .ZN(new_n469_));
  XOR2_X1   g268(.A(new_n468_), .B(new_n469_), .Z(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n462_), .A2(new_n466_), .A3(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n471_), .B1(new_n462_), .B2(new_n466_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT68), .ZN(new_n475_));
  OAI22_X1  g274(.A1(new_n473_), .A2(new_n474_), .B1(new_n475_), .B2(KEYINPUT13), .ZN(new_n476_));
  INV_X1    g275(.A(new_n474_), .ZN(new_n477_));
  XOR2_X1   g276(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(new_n472_), .A3(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n476_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G113gat), .B(G141gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G169gat), .B(G197gat), .ZN(new_n483_));
  XOR2_X1   g282(.A(new_n482_), .B(new_n483_), .Z(new_n484_));
  NAND2_X1  g283(.A1(G229gat), .A2(G233gat), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT77), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G29gat), .B(G36gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G43gat), .B(G50gat), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n488_), .A2(new_n489_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(G1gat), .ZN(new_n493_));
  INV_X1    g292(.A(G8gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G1gat), .A2(G8gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  AND2_X1   g296(.A1(G15gat), .A2(G22gat), .ZN(new_n498_));
  NOR2_X1   g297(.A1(G15gat), .A2(G22gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT14), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n501_), .B1(G1gat), .B2(G8gat), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n497_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G15gat), .B(G22gat), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n504_), .A2(new_n501_), .A3(new_n496_), .A4(new_n495_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n487_), .B1(new_n492_), .B2(new_n506_), .ZN(new_n507_));
  XOR2_X1   g306(.A(G29gat), .B(G36gat), .Z(new_n508_));
  XOR2_X1   g307(.A(G43gat), .B(G50gat), .Z(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n488_), .A2(new_n489_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n512_), .A2(KEYINPUT77), .A3(new_n503_), .A4(new_n505_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n507_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n492_), .A2(new_n506_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n514_), .A2(KEYINPUT78), .A3(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT78), .B1(new_n514_), .B2(new_n515_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n486_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT79), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT79), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n520_), .B(new_n486_), .C1(new_n516_), .C2(new_n517_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT15), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n523_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n510_), .A2(KEYINPUT15), .A3(new_n511_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n524_), .A2(new_n506_), .A3(new_n525_), .ZN(new_n526_));
  AND4_X1   g325(.A1(KEYINPUT80), .A2(new_n514_), .A3(new_n485_), .A4(new_n526_), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n526_), .A2(new_n485_), .ZN(new_n528_));
  AOI21_X1  g327(.A(KEYINPUT80), .B1(new_n528_), .B2(new_n514_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n484_), .B1(new_n522_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n484_), .ZN(new_n533_));
  AOI211_X1 g332(.A(new_n530_), .B(new_n533_), .C1(new_n519_), .C2(new_n521_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n532_), .A2(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n481_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n399_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT74), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n524_), .A2(new_n525_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n440_), .A2(new_n540_), .A3(new_n443_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G232gat), .A2(G233gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT70), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(KEYINPUT71), .B(KEYINPUT35), .Z(new_n547_));
  NOR2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n457_), .A2(new_n512_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n541_), .A2(KEYINPUT72), .A3(new_n548_), .A4(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G190gat), .B(G218gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G134gat), .B(G162gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  XOR2_X1   g352(.A(new_n553_), .B(KEYINPUT36), .Z(new_n554_));
  NAND2_X1  g353(.A1(new_n546_), .A2(new_n547_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n541_), .A2(new_n555_), .A3(new_n549_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n548_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT72), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n558_), .B1(new_n541_), .B2(new_n559_), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n550_), .B(new_n554_), .C1(new_n557_), .C2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT73), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n553_), .A2(KEYINPUT36), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n541_), .A2(new_n559_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n556_), .B1(new_n566_), .B2(new_n558_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n565_), .B1(new_n567_), .B2(new_n550_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n563_), .A2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(KEYINPUT37), .B1(new_n561_), .B2(new_n562_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n539_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n567_), .A2(KEYINPUT75), .A3(new_n550_), .A4(new_n554_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT75), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n561_), .A2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n572_), .B1(new_n574_), .B2(new_n568_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT37), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n570_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n550_), .B1(new_n557_), .B2(new_n560_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(new_n564_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n580_), .A2(new_n562_), .A3(new_n561_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n578_), .A2(KEYINPUT74), .A3(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n571_), .A2(new_n577_), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(G127gat), .B(G155gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT16), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G183gat), .B(G211gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n506_), .A2(G231gat), .A3(G233gat), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n503_), .A2(new_n505_), .A3(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n592_), .A2(new_n450_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n450_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n588_), .B1(new_n595_), .B2(KEYINPUT17), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n593_), .A2(KEYINPUT76), .A3(new_n594_), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n588_), .A2(KEYINPUT17), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n596_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n597_), .B1(new_n596_), .B2(new_n598_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n584_), .A2(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n538_), .A2(new_n603_), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n604_), .A2(new_n493_), .A3(new_n329_), .ZN(new_n605_));
  XOR2_X1   g404(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n606_));
  AND2_X1   g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NOR4_X1   g406(.A1(new_n399_), .A2(new_n602_), .A3(new_n575_), .A4(new_n537_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n493_), .B1(new_n608_), .B2(new_n329_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n610_), .B1(new_n605_), .B2(new_n606_), .ZN(G1324gat));
  INV_X1    g410(.A(new_n281_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n604_), .A2(new_n494_), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT39), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n608_), .A2(new_n612_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n614_), .B1(new_n615_), .B2(G8gat), .ZN(new_n616_));
  AOI211_X1 g415(.A(KEYINPUT39), .B(new_n494_), .C1(new_n608_), .C2(new_n612_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n613_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT40), .Z(G1325gat));
  NAND2_X1  g418(.A1(new_n608_), .A2(new_n377_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(G15gat), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n621_), .A2(KEYINPUT102), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(KEYINPUT102), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT41), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n604_), .A2(new_n360_), .A3(new_n377_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n622_), .A2(KEYINPUT41), .A3(new_n623_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n626_), .A2(new_n627_), .A3(new_n628_), .ZN(G1326gat));
  INV_X1    g428(.A(G22gat), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n630_), .B1(new_n608_), .B2(new_n397_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT42), .Z(new_n632_));
  NAND3_X1  g431(.A1(new_n604_), .A2(new_n630_), .A3(new_n397_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(G1327gat));
  OAI21_X1  g433(.A(KEYINPUT43), .B1(new_n399_), .B2(new_n583_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n272_), .A2(new_n276_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n279_), .A2(new_n280_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n381_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n396_), .A2(new_n398_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT43), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(new_n641_), .A3(new_n584_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n635_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n536_), .A2(new_n602_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT44), .B1(new_n643_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT44), .ZN(new_n647_));
  AOI211_X1 g446(.A(new_n647_), .B(new_n644_), .C1(new_n635_), .C2(new_n642_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(G29gat), .B1(new_n650_), .B2(new_n395_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n580_), .A2(new_n573_), .A3(new_n561_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n601_), .B1(new_n652_), .B2(new_n572_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n538_), .A2(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n395_), .A2(G29gat), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT103), .Z(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n651_), .A2(new_n657_), .ZN(G1328gat));
  INV_X1    g457(.A(KEYINPUT46), .ZN(new_n659_));
  INV_X1    g458(.A(G36gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n660_), .B1(new_n649_), .B2(new_n612_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n281_), .A2(G36gat), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n640_), .A2(new_n662_), .A3(new_n536_), .A4(new_n653_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n663_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT45), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n663_), .A2(new_n665_), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n666_), .A2(new_n667_), .A3(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n667_), .B1(new_n666_), .B2(new_n668_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n659_), .B1(new_n661_), .B2(new_n671_), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n646_), .A2(new_n648_), .A3(new_n281_), .ZN(new_n673_));
  OAI221_X1 g472(.A(KEYINPUT46), .B1(new_n669_), .B2(new_n670_), .C1(new_n673_), .C2(new_n660_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(G1329gat));
  AOI21_X1  g474(.A(G43gat), .B1(new_n654_), .B2(new_n377_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n377_), .A2(G43gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n649_), .B2(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n678_), .B(new_n679_), .ZN(G1330gat));
  AOI21_X1  g479(.A(G50gat), .B1(new_n654_), .B2(new_n397_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n397_), .A2(G50gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n649_), .B2(new_n682_), .ZN(G1331gat));
  NOR2_X1   g482(.A1(new_n399_), .A2(new_n575_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n535_), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n480_), .A2(new_n602_), .A3(new_n685_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n684_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(G57gat), .B1(new_n688_), .B2(new_n395_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n480_), .A2(new_n685_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n640_), .A2(new_n690_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n691_), .A2(new_n603_), .ZN(new_n692_));
  INV_X1    g491(.A(G57gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(new_n693_), .A3(new_n329_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n689_), .A2(new_n694_), .ZN(G1332gat));
  OAI21_X1  g494(.A(G64gat), .B1(new_n688_), .B2(new_n281_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(KEYINPUT107), .B(KEYINPUT48), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n696_), .B(new_n697_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n281_), .A2(G64gat), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT108), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n692_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n698_), .A2(new_n701_), .ZN(G1333gat));
  NOR2_X1   g501(.A1(new_n379_), .A2(G71gat), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT109), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n692_), .A2(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(G71gat), .B1(new_n688_), .B2(new_n379_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n706_), .A2(KEYINPUT49), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(KEYINPUT49), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n705_), .B1(new_n707_), .B2(new_n708_), .ZN(G1334gat));
  AOI21_X1  g508(.A(new_n338_), .B1(new_n687_), .B2(new_n397_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT50), .Z(new_n711_));
  NAND3_X1  g510(.A1(new_n692_), .A2(new_n338_), .A3(new_n397_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1335gat));
  NAND2_X1  g512(.A1(new_n691_), .A2(new_n653_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n715_), .A2(new_n431_), .A3(new_n329_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n643_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n690_), .A2(new_n602_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n717_), .A2(new_n395_), .A3(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n716_), .B1(new_n719_), .B2(new_n431_), .ZN(G1336gat));
  NAND3_X1  g519(.A1(new_n715_), .A2(new_n432_), .A3(new_n612_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n717_), .A2(new_n281_), .A3(new_n718_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n722_), .B2(new_n432_), .ZN(G1337gat));
  NAND2_X1  g522(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT111), .Z(new_n725_));
  NAND4_X1  g524(.A1(new_n643_), .A2(new_n602_), .A3(new_n377_), .A4(new_n690_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(G99gat), .ZN(new_n727_));
  INV_X1    g526(.A(new_n427_), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n714_), .A2(new_n728_), .A3(new_n379_), .ZN(new_n729_));
  OAI221_X1 g528(.A(new_n725_), .B1(KEYINPUT110), .B2(KEYINPUT51), .C1(new_n727_), .C2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n725_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n729_), .B1(G99gat), .B2(new_n726_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n731_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n730_), .A2(new_n734_), .ZN(G1338gat));
  NAND4_X1  g534(.A1(new_n643_), .A2(new_n602_), .A3(new_n397_), .A4(new_n690_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(G106gat), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT52), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n736_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n691_), .A2(new_n428_), .A3(new_n397_), .A4(new_n653_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT112), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n741_), .B(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n739_), .A2(new_n740_), .A3(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT53), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT53), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n739_), .A2(new_n743_), .A3(new_n746_), .A4(new_n740_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(G1339gat));
  INV_X1    g547(.A(KEYINPUT119), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n612_), .A2(new_n395_), .A3(new_n378_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n522_), .A2(new_n531_), .A3(new_n484_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n514_), .A2(new_n515_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT78), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n514_), .A2(KEYINPUT78), .A3(new_n515_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n485_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n514_), .A2(new_n486_), .A3(new_n526_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n758_), .A2(new_n533_), .A3(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n752_), .A2(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n761_), .A2(new_n473_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n456_), .A2(new_n463_), .A3(new_n458_), .A4(new_n459_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n460_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n462_), .A2(new_n765_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n459_), .A2(new_n458_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n767_), .A2(KEYINPUT55), .A3(new_n456_), .A4(new_n461_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n764_), .A2(new_n766_), .A3(new_n768_), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n769_), .A2(KEYINPUT56), .A3(new_n470_), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT56), .B1(new_n769_), .B2(new_n470_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n762_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT58), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n769_), .A2(new_n470_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT56), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n769_), .A2(KEYINPUT56), .A3(new_n470_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(KEYINPUT58), .A3(new_n762_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n584_), .A2(new_n774_), .A3(new_n780_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n535_), .A2(new_n473_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n782_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n761_), .B1(new_n477_), .B2(new_n472_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n652_), .A2(KEYINPUT57), .A3(new_n572_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT118), .B1(new_n786_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT118), .ZN(new_n790_));
  AOI211_X1 g589(.A(new_n790_), .B(new_n787_), .C1(new_n783_), .C2(new_n785_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n781_), .B1(new_n789_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT117), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n575_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n794_));
  XOR2_X1   g593(.A(KEYINPUT116), .B(KEYINPUT57), .Z(new_n795_));
  OAI21_X1  g594(.A(new_n793_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n795_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n784_), .B1(new_n779_), .B2(new_n782_), .ZN(new_n798_));
  OAI211_X1 g597(.A(KEYINPUT117), .B(new_n797_), .C1(new_n798_), .C2(new_n575_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n796_), .A2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n602_), .B1(new_n792_), .B2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT113), .B1(new_n535_), .B2(new_n601_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n520_), .B1(new_n757_), .B2(new_n486_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n521_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n531_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n533_), .ZN(new_n806_));
  AND4_X1   g605(.A1(KEYINPUT113), .A2(new_n806_), .A3(new_n601_), .A4(new_n752_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n802_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT114), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n808_), .A2(new_n809_), .A3(new_n480_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(new_n808_), .B2(new_n480_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n583_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n583_), .B(new_n813_), .C1(new_n810_), .C2(new_n811_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  AOI211_X1 g617(.A(new_n535_), .B(new_n751_), .C1(new_n801_), .C2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n749_), .B1(new_n819_), .B2(G113gat), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n751_), .B1(new_n801_), .B2(new_n818_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n685_), .ZN(new_n822_));
  INV_X1    g621(.A(G113gat), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n822_), .A2(KEYINPUT119), .A3(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n820_), .A2(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n751_), .A2(KEYINPUT59), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n790_), .B1(new_n798_), .B2(new_n787_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n786_), .A2(KEYINPUT118), .A3(new_n788_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n583_), .B1(new_n773_), .B2(new_n772_), .ZN(new_n829_));
  AOI22_X1  g628(.A1(new_n827_), .A2(new_n828_), .B1(new_n829_), .B2(new_n780_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n797_), .B1(new_n798_), .B2(new_n575_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n601_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n826_), .B1(new_n832_), .B2(new_n817_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT120), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT59), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n833_), .B(new_n834_), .C1(new_n821_), .C2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n827_), .A2(new_n828_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n838_), .A2(new_n781_), .A3(new_n796_), .A4(new_n799_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n817_), .B1(new_n839_), .B2(new_n602_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT59), .B1(new_n840_), .B2(new_n751_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n834_), .B1(new_n841_), .B2(new_n833_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n837_), .A2(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n535_), .A2(new_n823_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n825_), .B1(new_n843_), .B2(new_n844_), .ZN(G1340gat));
  INV_X1    g644(.A(G120gat), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(new_n480_), .B2(KEYINPUT60), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n821_), .B(new_n847_), .C1(KEYINPUT60), .C2(new_n846_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n841_), .A2(new_n481_), .A3(new_n833_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n848_), .B1(new_n850_), .B2(new_n846_), .ZN(G1341gat));
  AOI21_X1  g650(.A(G127gat), .B1(new_n821_), .B2(new_n601_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n601_), .A2(G127gat), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n843_), .B2(new_n853_), .ZN(G1342gat));
  AOI21_X1  g653(.A(G134gat), .B1(new_n821_), .B2(new_n575_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n584_), .A2(G134gat), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n855_), .B1(new_n843_), .B2(new_n856_), .ZN(G1343gat));
  NAND2_X1  g656(.A1(new_n801_), .A2(new_n818_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n612_), .A2(new_n395_), .A3(new_n380_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(KEYINPUT121), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(new_n535_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(new_n283_), .ZN(G1344gat));
  NOR2_X1   g662(.A1(new_n861_), .A2(new_n480_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT122), .B(G148gat), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1345gat));
  OAI21_X1  g665(.A(KEYINPUT123), .B1(new_n861_), .B2(new_n602_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT123), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n858_), .A2(new_n868_), .A3(new_n860_), .A4(new_n601_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(KEYINPUT61), .B(G155gat), .ZN(new_n870_));
  AND3_X1   g669(.A1(new_n867_), .A2(new_n869_), .A3(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n867_), .B2(new_n869_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1346gat));
  OAI21_X1  g672(.A(G162gat), .B1(new_n861_), .B2(new_n583_), .ZN(new_n874_));
  INV_X1    g673(.A(G162gat), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n575_), .A2(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n874_), .B1(new_n861_), .B2(new_n876_), .ZN(G1347gat));
  XNOR2_X1  g676(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n830_), .A2(new_n831_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n602_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n818_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n281_), .A2(new_n329_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(new_n378_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n881_), .A2(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n535_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n878_), .B1(new_n886_), .B2(new_n215_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n878_), .ZN(new_n888_));
  OAI211_X1 g687(.A(G169gat), .B(new_n888_), .C1(new_n885_), .C2(new_n535_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n886_), .A2(new_n229_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n887_), .A2(new_n889_), .A3(new_n890_), .ZN(G1348gat));
  INV_X1    g690(.A(new_n885_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n481_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n840_), .A2(new_n397_), .ZN(new_n894_));
  NOR4_X1   g693(.A1(new_n883_), .A2(new_n216_), .A3(new_n379_), .A4(new_n480_), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n893_), .A2(new_n228_), .B1(new_n894_), .B2(new_n895_), .ZN(G1349gat));
  NOR3_X1   g695(.A1(new_n885_), .A2(new_n602_), .A3(new_n247_), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n894_), .A2(new_n601_), .A3(new_n377_), .A4(new_n882_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n897_), .B1(new_n208_), .B2(new_n898_), .ZN(G1350gat));
  OAI21_X1  g698(.A(G190gat), .B1(new_n885_), .B2(new_n583_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n575_), .A2(new_n207_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n885_), .B2(new_n901_), .ZN(G1351gat));
  NOR3_X1   g701(.A1(new_n840_), .A2(new_n380_), .A3(new_n883_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n685_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(KEYINPUT125), .A2(G197gat), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT125), .B(G197gat), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n904_), .B2(new_n907_), .ZN(G1352gat));
  NAND2_X1  g707(.A1(new_n903_), .A2(new_n481_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g709(.A(new_n602_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n903_), .A2(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(KEYINPUT126), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n912_), .B(new_n914_), .ZN(G1354gat));
  NAND2_X1  g714(.A1(new_n903_), .A2(new_n575_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(KEYINPUT127), .B(G218gat), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n583_), .A2(new_n917_), .ZN(new_n918_));
  AOI22_X1  g717(.A1(new_n916_), .A2(new_n917_), .B1(new_n903_), .B2(new_n918_), .ZN(G1355gat));
endmodule


