//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 0 0 1 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n788_, new_n789_, new_n790_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n921_, new_n922_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(G169gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT84), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n208_), .B1(new_n209_), .B2(KEYINPUT23), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(KEYINPUT23), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G183gat), .A3(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n210_), .B1(new_n214_), .B2(new_n208_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n207_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT25), .B(G183gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT26), .B(G190gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  OR2_X1    g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n221_), .A2(KEYINPUT24), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n221_), .A2(KEYINPUT24), .A3(new_n224_), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n220_), .A2(new_n223_), .A3(new_n214_), .A4(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n217_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT85), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n217_), .A2(KEYINPUT85), .A3(new_n226_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(G71gat), .B(G99gat), .Z(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(G43gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT30), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n231_), .B(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G227gat), .A2(G233gat), .ZN(new_n237_));
  INV_X1    g036(.A(G15gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(KEYINPUT86), .B1(new_n236_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT31), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n235_), .A2(new_n239_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n242_), .B1(new_n241_), .B2(new_n243_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n205_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n241_), .A2(new_n243_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT31), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(new_n204_), .A3(new_n244_), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n247_), .A2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G211gat), .B(G218gat), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT89), .ZN(new_n254_));
  INV_X1    g053(.A(G197gat), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n254_), .B1(new_n255_), .B2(G204gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(G204gat), .ZN(new_n257_));
  INV_X1    g056(.A(G204gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(KEYINPUT89), .A3(G197gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n256_), .A2(new_n257_), .A3(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n253_), .A2(new_n260_), .A3(KEYINPUT21), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT90), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT21), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n256_), .A2(new_n259_), .A3(new_n264_), .A4(new_n257_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G197gat), .B(G204gat), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n252_), .B1(new_n267_), .B2(new_n264_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n263_), .B1(new_n266_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n257_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n255_), .A2(G204gat), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT21), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n272_), .A2(new_n265_), .A3(KEYINPUT90), .A4(new_n252_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n262_), .B1(new_n269_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G141gat), .A2(G148gat), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT87), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT2), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT2), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n275_), .A2(new_n276_), .A3(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(G141gat), .A2(G148gat), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT3), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n278_), .A2(new_n280_), .A3(new_n283_), .A4(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(G155gat), .B(G162gat), .Z(new_n286_));
  INV_X1    g085(.A(KEYINPUT1), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n281_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n290_));
  AND3_X1   g089(.A1(new_n289_), .A2(new_n275_), .A3(new_n290_), .ZN(new_n291_));
  AOI22_X1  g090(.A1(new_n285_), .A2(new_n286_), .B1(new_n288_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT29), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G228gat), .A2(G233gat), .ZN(new_n295_));
  AOI211_X1 g094(.A(new_n274_), .B(new_n294_), .C1(KEYINPUT88), .C2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n295_), .B1(new_n274_), .B2(KEYINPUT88), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n294_), .A2(new_n274_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G78gat), .B(G106gat), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NOR3_X1   g100(.A1(new_n296_), .A2(new_n299_), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n301_), .B1(new_n296_), .B2(new_n299_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n292_), .A2(new_n293_), .ZN(new_n306_));
  XOR2_X1   g105(.A(G22gat), .B(G50gat), .Z(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT28), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n306_), .B(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT91), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n309_), .B1(new_n302_), .B2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n305_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G1gat), .B(G29gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT97), .B(G85gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT0), .B(G57gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G225gat), .A2(G233gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT96), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n292_), .A2(new_n320_), .A3(new_n204_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n204_), .B1(new_n292_), .B2(new_n320_), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT4), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NOR3_X1   g122(.A1(new_n205_), .A2(new_n292_), .A3(KEYINPUT4), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n319_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n285_), .A2(new_n286_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n288_), .A2(new_n291_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n205_), .B1(new_n329_), .B2(KEYINPUT96), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n292_), .A2(new_n320_), .A3(new_n204_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n319_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n318_), .B1(new_n326_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT4), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n336_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n333_), .B1(new_n337_), .B2(new_n324_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n334_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n338_), .A2(new_n339_), .A3(new_n317_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n335_), .A2(new_n340_), .A3(KEYINPUT98), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT98), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n338_), .A2(new_n339_), .A3(new_n342_), .A4(new_n317_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n303_), .A2(new_n310_), .A3(new_n304_), .A4(new_n309_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n312_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT93), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n347_), .B1(new_n215_), .B2(new_n222_), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT84), .B1(new_n211_), .B2(new_n213_), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n223_), .B(KEYINPUT93), .C1(new_n349_), .C2(new_n210_), .ZN(new_n350_));
  XOR2_X1   g149(.A(KEYINPUT26), .B(G190gat), .Z(new_n351_));
  INV_X1    g150(.A(KEYINPUT92), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n219_), .A2(KEYINPUT92), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(new_n218_), .A3(new_n354_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n348_), .A2(new_n225_), .A3(new_n350_), .A4(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n214_), .B1(G183gat), .B2(G190gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(new_n207_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n356_), .A2(new_n274_), .A3(new_n358_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n359_), .A2(KEYINPUT20), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT19), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n269_), .A2(new_n273_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(new_n261_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n217_), .A2(KEYINPUT85), .A3(new_n226_), .ZN(new_n366_));
  AOI21_X1  g165(.A(KEYINPUT85), .B1(new_n217_), .B2(new_n226_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n365_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n360_), .A2(KEYINPUT95), .A3(new_n363_), .A4(new_n368_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n368_), .A2(KEYINPUT20), .A3(new_n363_), .A4(new_n359_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT95), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n369_), .A2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G8gat), .B(G36gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT18), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G64gat), .B(G92gat), .ZN(new_n376_));
  XOR2_X1   g175(.A(new_n375_), .B(new_n376_), .Z(new_n377_));
  NAND2_X1  g176(.A1(new_n356_), .A2(new_n358_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(new_n365_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n229_), .A2(new_n274_), .A3(new_n230_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(KEYINPUT20), .A3(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(KEYINPUT94), .B1(new_n381_), .B2(new_n362_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT94), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT20), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n384_), .B1(new_n378_), .B2(new_n365_), .ZN(new_n385_));
  AOI211_X1 g184(.A(new_n383_), .B(new_n363_), .C1(new_n385_), .C2(new_n380_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n373_), .B(new_n377_), .C1(new_n382_), .C2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT27), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n359_), .A2(KEYINPUT20), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n274_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n362_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n391_), .B1(new_n362_), .B2(new_n381_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n377_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n388_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n387_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT99), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n387_), .A2(KEYINPUT99), .A3(new_n394_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n346_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n386_), .A2(new_n382_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n370_), .B(KEYINPUT95), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n393_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n387_), .ZN(new_n403_));
  AOI21_X1  g202(.A(KEYINPUT100), .B1(new_n403_), .B2(new_n388_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT100), .ZN(new_n405_));
  AOI211_X1 g204(.A(new_n405_), .B(KEYINPUT27), .C1(new_n402_), .C2(new_n387_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n399_), .B1(new_n404_), .B2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n323_), .A2(new_n319_), .A3(new_n325_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n318_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n317_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n410_), .B1(new_n411_), .B2(KEYINPUT33), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n412_), .B1(KEYINPUT33), .B2(new_n411_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n413_), .A2(new_n387_), .A3(new_n402_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n344_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n377_), .A2(KEYINPUT32), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n373_), .B(new_n416_), .C1(new_n382_), .C2(new_n386_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n392_), .A2(KEYINPUT32), .A3(new_n377_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n415_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n414_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n312_), .A2(new_n345_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n251_), .B1(new_n407_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n397_), .A2(new_n398_), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n421_), .B(new_n424_), .C1(new_n404_), .C2(new_n406_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n247_), .A2(new_n250_), .A3(new_n344_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n423_), .A2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G29gat), .B(G36gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT73), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G43gat), .B(G50gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT73), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n429_), .B(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n431_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n432_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G15gat), .B(G22gat), .ZN(new_n438_));
  INV_X1    g237(.A(G1gat), .ZN(new_n439_));
  INV_X1    g238(.A(G8gat), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT14), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n438_), .A2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G1gat), .B(G8gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  XOR2_X1   g243(.A(new_n437_), .B(new_n444_), .Z(new_n445_));
  NAND2_X1  g244(.A1(G229gat), .A2(G233gat), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n432_), .A2(new_n436_), .A3(KEYINPUT15), .ZN(new_n449_));
  AOI21_X1  g248(.A(KEYINPUT15), .B1(new_n432_), .B2(new_n436_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n444_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT82), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n437_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n456_), .A2(new_n444_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n446_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n448_), .B1(new_n455_), .B2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G113gat), .B(G141gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G169gat), .B(G197gat), .ZN(new_n462_));
  XOR2_X1   g261(.A(new_n461_), .B(new_n462_), .Z(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n460_), .A2(new_n464_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n448_), .B(new_n463_), .C1(new_n455_), .C2(new_n459_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT83), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n465_), .A2(KEYINPUT83), .A3(new_n466_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n428_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT79), .ZN(new_n473_));
  XOR2_X1   g272(.A(G190gat), .B(G218gat), .Z(new_n474_));
  XNOR2_X1  g273(.A(G134gat), .B(G162gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT36), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G232gat), .A2(G233gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT34), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT35), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT8), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G99gat), .A2(G106gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT6), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n489_), .A2(G99gat), .A3(G106gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT70), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT70), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n488_), .A2(new_n490_), .A3(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(G99gat), .A2(G106gat), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT68), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n496_), .A2(KEYINPUT7), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(KEYINPUT7), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n495_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n498_), .A2(new_n495_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n492_), .A2(new_n494_), .A3(new_n499_), .A4(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G85gat), .B(G92gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT69), .ZN(new_n503_));
  INV_X1    g302(.A(G85gat), .ZN(new_n504_));
  INV_X1    g303(.A(G92gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT69), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G85gat), .A2(G92gat), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n506_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n503_), .A2(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n486_), .B1(new_n501_), .B2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(KEYINPUT8), .B1(new_n503_), .B2(new_n509_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n499_), .A2(new_n500_), .A3(new_n491_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n515_), .A2(KEYINPUT67), .ZN(new_n516_));
  INV_X1    g315(.A(new_n515_), .ZN(new_n517_));
  AOI21_X1  g316(.A(KEYINPUT67), .B1(new_n504_), .B2(new_n505_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n516_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT66), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n505_), .A2(KEYINPUT65), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT65), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(G92gat), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n504_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n520_), .B1(new_n524_), .B2(KEYINPUT9), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT9), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT65), .B(G92gat), .ZN(new_n527_));
  OAI211_X1 g326(.A(KEYINPUT66), .B(new_n526_), .C1(new_n527_), .C2(new_n504_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n519_), .B1(new_n525_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT64), .ZN(new_n530_));
  XOR2_X1   g329(.A(KEYINPUT10), .B(G99gat), .Z(new_n531_));
  INV_X1    g330(.A(G106gat), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n530_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT10), .B(G99gat), .ZN(new_n534_));
  NOR3_X1   g333(.A1(new_n534_), .A2(KEYINPUT64), .A3(G106gat), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n491_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n536_));
  OAI22_X1  g335(.A1(new_n511_), .A2(new_n514_), .B1(new_n529_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT71), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  OAI221_X1 g338(.A(KEYINPUT71), .B1(new_n529_), .B2(new_n536_), .C1(new_n511_), .C2(new_n514_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n539_), .A2(new_n437_), .A3(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT74), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT74), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n539_), .A2(new_n540_), .A3(new_n543_), .A4(new_n437_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n537_), .ZN(new_n546_));
  OAI22_X1  g345(.A1(new_n451_), .A2(new_n546_), .B1(KEYINPUT35), .B2(new_n481_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n485_), .B1(new_n545_), .B2(new_n548_), .ZN(new_n549_));
  AOI211_X1 g348(.A(new_n484_), .B(new_n547_), .C1(new_n542_), .C2(new_n544_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n479_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n545_), .A2(new_n548_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(new_n484_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n545_), .A2(new_n485_), .A3(new_n548_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n478_), .ZN(new_n556_));
  XOR2_X1   g355(.A(KEYINPUT77), .B(KEYINPUT36), .Z(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n554_), .A2(new_n555_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT78), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n549_), .A2(new_n550_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n562_), .A2(KEYINPUT78), .A3(new_n558_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n552_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT37), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n473_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT78), .B1(new_n562_), .B2(new_n558_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n558_), .ZN(new_n568_));
  NOR4_X1   g367(.A1(new_n549_), .A2(new_n550_), .A3(new_n560_), .A4(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n551_), .B1(new_n567_), .B2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(KEYINPUT79), .A3(KEYINPUT37), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n561_), .A2(new_n563_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n551_), .A2(KEYINPUT80), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n551_), .A2(KEYINPUT80), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(KEYINPUT81), .B(KEYINPUT37), .Z(new_n576_));
  AOI22_X1  g375(.A1(new_n566_), .A2(new_n571_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n539_), .A2(new_n540_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G57gat), .B(G64gat), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n579_), .A2(KEYINPUT11), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(KEYINPUT11), .ZN(new_n581_));
  XOR2_X1   g380(.A(G71gat), .B(G78gat), .Z(new_n582_));
  NAND3_X1  g381(.A1(new_n580_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n581_), .A2(new_n582_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n578_), .A2(new_n585_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n537_), .A2(KEYINPUT12), .A3(new_n584_), .A4(new_n583_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G230gat), .A2(G233gat), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n578_), .A2(new_n585_), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n588_), .B(new_n589_), .C1(KEYINPUT12), .C2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n589_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n586_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n592_), .B1(new_n593_), .B2(new_n590_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n591_), .A2(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(G120gat), .B(G148gat), .Z(new_n596_));
  XNOR2_X1  g395(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G176gat), .B(G204gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n595_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n600_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n591_), .A2(new_n594_), .A3(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT13), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(KEYINPUT13), .B1(new_n601_), .B2(new_n603_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n585_), .B(new_n444_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n609_), .B(new_n610_), .Z(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT17), .ZN(new_n613_));
  XOR2_X1   g412(.A(G127gat), .B(G155gat), .Z(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT16), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G183gat), .B(G211gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  OR3_X1    g416(.A1(new_n612_), .A2(new_n613_), .A3(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(KEYINPUT17), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n612_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n608_), .A2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n577_), .A2(new_n623_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n472_), .A2(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n625_), .A2(new_n439_), .A3(new_n415_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT38), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT101), .Z(new_n629_));
  NOR4_X1   g428(.A1(new_n428_), .A2(new_n623_), .A3(new_n471_), .A4(new_n575_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G1gat), .B1(new_n631_), .B2(new_n344_), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n629_), .B(new_n632_), .C1(new_n627_), .C2(new_n626_), .ZN(G1324gat));
  NAND2_X1  g432(.A1(new_n403_), .A2(new_n388_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(new_n405_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n403_), .A2(KEYINPUT100), .A3(new_n388_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(new_n424_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n440_), .B1(new_n630_), .B2(new_n638_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT39), .Z(new_n640_));
  NAND3_X1  g439(.A1(new_n625_), .A2(new_n440_), .A3(new_n638_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT40), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(G1325gat));
  NAND2_X1  g443(.A1(new_n630_), .A2(new_n251_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(G15gat), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT102), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n645_), .A2(new_n648_), .A3(G15gat), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT41), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n625_), .A2(new_n238_), .A3(new_n251_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n647_), .A2(KEYINPUT41), .A3(new_n649_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n652_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT103), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT103), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n652_), .A2(new_n657_), .A3(new_n653_), .A4(new_n654_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(G1326gat));
  INV_X1    g458(.A(G22gat), .ZN(new_n660_));
  INV_X1    g459(.A(new_n421_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n630_), .B2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n625_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1327gat));
  INV_X1    g465(.A(new_n608_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n575_), .A2(new_n621_), .ZN(new_n668_));
  NOR4_X1   g467(.A1(new_n428_), .A2(new_n667_), .A3(new_n471_), .A4(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(G29gat), .B1(new_n669_), .B2(new_n415_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n471_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n608_), .A2(new_n671_), .A3(new_n621_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .A4(new_n576_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n564_), .A2(new_n473_), .A3(new_n565_), .ZN(new_n675_));
  AOI21_X1  g474(.A(KEYINPUT79), .B1(new_n570_), .B2(KEYINPUT37), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n674_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n428_), .A2(new_n677_), .A3(KEYINPUT43), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n247_), .A2(new_n250_), .A3(new_n344_), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n637_), .A2(new_n680_), .A3(new_n421_), .A4(new_n424_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n661_), .B1(new_n414_), .B2(new_n419_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n637_), .B2(new_n399_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n681_), .B1(new_n683_), .B2(new_n251_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n679_), .B1(new_n684_), .B2(new_n577_), .ZN(new_n685_));
  OAI211_X1 g484(.A(KEYINPUT44), .B(new_n673_), .C1(new_n678_), .C2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(KEYINPUT43), .B1(new_n428_), .B2(new_n677_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n684_), .A2(new_n577_), .A3(new_n679_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n672_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n691_), .A2(KEYINPUT105), .A3(KEYINPUT44), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n688_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n415_), .A2(G29gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n673_), .B1(new_n678_), .B2(new_n685_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n694_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n670_), .B1(new_n693_), .B2(new_n697_), .ZN(G1328gat));
  INV_X1    g497(.A(G36gat), .ZN(new_n699_));
  AOI22_X1  g498(.A1(new_n688_), .A2(new_n692_), .B1(new_n696_), .B2(new_n695_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n700_), .B2(new_n638_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n669_), .A2(new_n699_), .A3(new_n638_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT45), .Z(new_n703_));
  NOR2_X1   g502(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n704_));
  OR3_X1    g503(.A1(new_n701_), .A2(new_n703_), .A3(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n704_), .B1(new_n701_), .B2(new_n703_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1329gat));
  XNOR2_X1  g506(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n251_), .A2(G43gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n686_), .A2(new_n687_), .ZN(new_n711_));
  AOI21_X1  g510(.A(KEYINPUT105), .B1(new_n691_), .B2(KEYINPUT44), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n710_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT107), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n693_), .A2(new_n715_), .A3(new_n710_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(G43gat), .B1(new_n669_), .B2(new_n251_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n708_), .B1(new_n717_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n708_), .ZN(new_n721_));
  AOI211_X1 g520(.A(new_n718_), .B(new_n721_), .C1(new_n714_), .C2(new_n716_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1330gat));
  AOI21_X1  g522(.A(G50gat), .B1(new_n669_), .B2(new_n661_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n661_), .A2(G50gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n700_), .B2(new_n725_), .ZN(G1331gat));
  NOR2_X1   g525(.A1(new_n428_), .A2(new_n671_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n608_), .A2(new_n621_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT109), .ZN(new_n730_));
  INV_X1    g529(.A(new_n575_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n729_), .A2(new_n730_), .A3(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n727_), .A2(new_n728_), .ZN(new_n733_));
  OAI21_X1  g532(.A(KEYINPUT109), .B1(new_n733_), .B2(new_n575_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(KEYINPUT110), .B(G57gat), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n344_), .A2(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n732_), .A2(new_n734_), .A3(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT111), .ZN(new_n738_));
  INV_X1    g537(.A(G57gat), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n729_), .A2(new_n677_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n740_), .B2(new_n344_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n738_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT112), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n738_), .A2(KEYINPUT112), .A3(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1332gat));
  INV_X1    g545(.A(KEYINPUT48), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n732_), .A2(new_n734_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(new_n638_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n747_), .B1(new_n749_), .B2(G64gat), .ZN(new_n750_));
  INV_X1    g549(.A(G64gat), .ZN(new_n751_));
  AOI211_X1 g550(.A(KEYINPUT48), .B(new_n751_), .C1(new_n748_), .C2(new_n638_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n638_), .A2(new_n751_), .ZN(new_n753_));
  OAI22_X1  g552(.A1(new_n750_), .A2(new_n752_), .B1(new_n740_), .B2(new_n753_), .ZN(G1333gat));
  INV_X1    g553(.A(new_n251_), .ZN(new_n755_));
  OR3_X1    g554(.A1(new_n740_), .A2(G71gat), .A3(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n732_), .A2(new_n251_), .A3(new_n734_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT49), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n757_), .A2(new_n758_), .A3(G71gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n757_), .B2(G71gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n756_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  OAI211_X1 g562(.A(KEYINPUT113), .B(new_n756_), .C1(new_n759_), .C2(new_n760_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(G1334gat));
  OR3_X1    g564(.A1(new_n740_), .A2(G78gat), .A3(new_n421_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n748_), .A2(new_n661_), .ZN(new_n767_));
  XOR2_X1   g566(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n768_));
  AND3_X1   g567(.A1(new_n767_), .A2(G78gat), .A3(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(new_n767_), .B2(G78gat), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n766_), .B1(new_n769_), .B2(new_n770_), .ZN(G1335gat));
  NOR2_X1   g570(.A1(new_n668_), .A2(new_n608_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n727_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(G85gat), .B1(new_n774_), .B2(new_n415_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n608_), .A2(new_n671_), .A3(new_n622_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT115), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n689_), .A2(new_n690_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT116), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT116), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n777_), .A2(new_n781_), .A3(new_n778_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n344_), .A2(new_n504_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT117), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n775_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT118), .ZN(G1336gat));
  AOI21_X1  g586(.A(G92gat), .B1(new_n774_), .B2(new_n638_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n638_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n789_), .A2(new_n527_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n788_), .B1(new_n783_), .B2(new_n790_), .ZN(G1337gat));
  NOR3_X1   g590(.A1(new_n773_), .A2(new_n755_), .A3(new_n534_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(KEYINPUT119), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n755_), .B1(new_n780_), .B2(new_n782_), .ZN(new_n794_));
  INV_X1    g593(.A(G99gat), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n793_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n797_), .A2(KEYINPUT120), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n796_), .B(new_n798_), .ZN(G1338gat));
  NAND3_X1  g598(.A1(new_n774_), .A2(new_n532_), .A3(new_n661_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n777_), .A2(new_n661_), .A3(new_n778_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(G106gat), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n802_), .A2(KEYINPUT52), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n802_), .A2(KEYINPUT52), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n800_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n586_), .B(new_n587_), .C1(new_n590_), .C2(KEYINPUT12), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n807_), .B1(new_n808_), .B2(new_n592_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n808_), .A2(new_n592_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n808_), .A2(new_n807_), .A3(new_n592_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n600_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT56), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT122), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n813_), .A2(KEYINPUT122), .A3(new_n814_), .ZN(new_n818_));
  OAI211_X1 g617(.A(KEYINPUT56), .B(new_n600_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n817_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n603_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n463_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n458_), .A2(new_n447_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n455_), .B2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n466_), .A2(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n821_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n820_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT58), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n820_), .A2(KEYINPUT58), .A3(new_n826_), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n829_), .A2(new_n577_), .A3(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n469_), .A2(new_n470_), .A3(new_n603_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n832_), .B1(new_n819_), .B2(new_n815_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n825_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n602_), .B1(new_n591_), .B2(new_n594_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n821_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT121), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n604_), .A2(KEYINPUT121), .A3(new_n834_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n731_), .B1(new_n833_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  OAI211_X1 g642(.A(KEYINPUT57), .B(new_n731_), .C1(new_n833_), .C2(new_n840_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n621_), .B1(new_n831_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n847_), .B1(new_n624_), .B2(new_n471_), .ZN(new_n848_));
  NOR4_X1   g647(.A1(new_n577_), .A2(new_n623_), .A3(KEYINPUT54), .A4(new_n671_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n846_), .A2(new_n851_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n755_), .A2(new_n425_), .A3(new_n344_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(G113gat), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n854_), .A2(new_n855_), .A3(new_n671_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n852_), .A2(KEYINPUT123), .A3(new_n853_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n852_), .A2(KEYINPUT123), .A3(KEYINPUT59), .A4(new_n853_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n471_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n856_), .B1(new_n861_), .B2(new_n855_), .ZN(G1340gat));
  INV_X1    g661(.A(G120gat), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n608_), .B2(KEYINPUT60), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n854_), .B(new_n864_), .C1(KEYINPUT60), .C2(new_n863_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n608_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(new_n863_), .ZN(G1341gat));
  INV_X1    g666(.A(G127gat), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n854_), .A2(new_n868_), .A3(new_n622_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n621_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n870_), .B2(new_n868_), .ZN(G1342gat));
  INV_X1    g670(.A(G134gat), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n854_), .A2(new_n872_), .A3(new_n575_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n677_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n874_), .B2(new_n872_), .ZN(G1343gat));
  NAND3_X1  g674(.A1(new_n789_), .A2(new_n661_), .A3(new_n415_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n843_), .A2(new_n844_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n829_), .A2(new_n577_), .A3(new_n830_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n622_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n755_), .B(new_n877_), .C1(new_n880_), .C2(new_n850_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n471_), .ZN(new_n882_));
  XOR2_X1   g681(.A(new_n882_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g682(.A1(new_n881_), .A2(new_n608_), .ZN(new_n884_));
  XOR2_X1   g683(.A(new_n884_), .B(G148gat), .Z(G1345gat));
  OAI21_X1  g684(.A(KEYINPUT124), .B1(new_n881_), .B2(new_n621_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n251_), .B1(new_n846_), .B2(new_n851_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT124), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n887_), .A2(new_n888_), .A3(new_n622_), .A4(new_n877_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n886_), .A2(new_n889_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(KEYINPUT61), .B(G155gat), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n892_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n886_), .A2(new_n889_), .A3(new_n891_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1346gat));
  OAI21_X1  g694(.A(G162gat), .B1(new_n881_), .B2(new_n677_), .ZN(new_n896_));
  OR2_X1    g695(.A1(new_n731_), .A2(G162gat), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n881_), .B2(new_n897_), .ZN(G1347gat));
  NOR3_X1   g697(.A1(new_n789_), .A2(new_n661_), .A3(new_n426_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n852_), .A2(new_n671_), .A3(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(KEYINPUT62), .B1(new_n900_), .B2(KEYINPUT22), .ZN(new_n901_));
  OAI21_X1  g700(.A(G169gat), .B1(new_n900_), .B2(KEYINPUT62), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(G169gat), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n904_), .B2(new_n901_), .ZN(G1348gat));
  AND2_X1   g704(.A1(KEYINPUT125), .A2(G176gat), .ZN(new_n906_));
  NOR2_X1   g705(.A1(KEYINPUT125), .A2(G176gat), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n852_), .A2(new_n667_), .A3(new_n899_), .ZN(new_n909_));
  MUX2_X1   g708(.A(new_n908_), .B(new_n906_), .S(new_n909_), .Z(G1349gat));
  NAND2_X1  g709(.A1(new_n852_), .A2(new_n899_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(G183gat), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(KEYINPUT126), .ZN(new_n914_));
  NAND4_X1  g713(.A1(new_n912_), .A2(new_n218_), .A3(new_n622_), .A4(new_n914_), .ZN(new_n915_));
  OAI22_X1  g714(.A1(new_n911_), .A2(new_n621_), .B1(KEYINPUT126), .B2(G183gat), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1350gat));
  OAI21_X1  g716(.A(G190gat), .B1(new_n911_), .B2(new_n677_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n575_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n911_), .B2(new_n919_), .ZN(G1351gat));
  NOR2_X1   g719(.A1(new_n789_), .A2(new_n346_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n887_), .A2(new_n671_), .A3(new_n921_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g722(.A1(new_n887_), .A2(new_n667_), .A3(new_n921_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g724(.A(new_n621_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(KEYINPUT127), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n887_), .A2(new_n921_), .A3(new_n928_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n930_));
  XOR2_X1   g729(.A(new_n929_), .B(new_n930_), .Z(G1354gat));
  NAND2_X1  g730(.A1(new_n887_), .A2(new_n921_), .ZN(new_n932_));
  OAI21_X1  g731(.A(G218gat), .B1(new_n932_), .B2(new_n677_), .ZN(new_n933_));
  OR2_X1    g732(.A1(new_n731_), .A2(G218gat), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n933_), .B1(new_n932_), .B2(new_n934_), .ZN(G1355gat));
endmodule


