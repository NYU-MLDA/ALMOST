//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n903_, new_n904_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n931_, new_n932_, new_n933_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n944_,
    new_n945_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT31), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT23), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT80), .B(G183gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT81), .B(G190gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n205_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G176gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT22), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n209_), .B1(new_n210_), .B2(KEYINPUT84), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G169gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n213_), .B1(KEYINPUT84), .B2(new_n210_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n208_), .A2(new_n212_), .A3(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT82), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT24), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT82), .B1(G169gat), .B2(G176gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n221_), .B1(new_n206_), .B2(KEYINPUT25), .ZN(new_n222_));
  NOR2_X1   g021(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n223_), .B1(new_n207_), .B2(KEYINPUT26), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n205_), .B(new_n220_), .C1(new_n222_), .C2(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n218_), .B1(G169gat), .B2(G176gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n219_), .ZN(new_n227_));
  NOR3_X1   g026(.A1(KEYINPUT82), .A2(G169gat), .A3(G176gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n226_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT83), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n217_), .A2(new_n219_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n232_), .A2(KEYINPUT83), .A3(new_n226_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n215_), .B1(new_n225_), .B2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT30), .ZN(new_n236_));
  INV_X1    g035(.A(G71gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT30), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n238_), .B(new_n215_), .C1(new_n225_), .C2(new_n234_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n236_), .A2(new_n237_), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n237_), .B1(new_n236_), .B2(new_n239_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT85), .B(G99gat), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NOR3_X1   g043(.A1(new_n241_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n236_), .A2(new_n239_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(G71gat), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n243_), .B1(new_n247_), .B2(new_n240_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n203_), .B1(new_n245_), .B2(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(G127gat), .B(G134gat), .Z(new_n250_));
  INV_X1    g049(.A(G113gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G127gat), .B(G134gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(G113gat), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n252_), .A2(G120gat), .A3(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(G120gat), .B1(new_n252_), .B2(new_n254_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G227gat), .A2(G233gat), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n257_), .B(new_n258_), .Z(new_n259_));
  OAI21_X1  g058(.A(new_n244_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n247_), .A2(new_n240_), .A3(new_n243_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n203_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n249_), .A2(new_n259_), .A3(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n259_), .B1(new_n249_), .B2(new_n263_), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G226gat), .A2(G233gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT19), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G211gat), .B(G218gat), .ZN(new_n270_));
  INV_X1    g069(.A(G197gat), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n271_), .A2(G204gat), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n270_), .B(KEYINPUT21), .C1(KEYINPUT91), .C2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G197gat), .B(G204gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  OR2_X1    g074(.A1(new_n270_), .A2(KEYINPUT21), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n272_), .A2(KEYINPUT91), .ZN(new_n277_));
  INV_X1    g076(.A(new_n274_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n277_), .A2(new_n278_), .A3(KEYINPUT21), .A4(new_n270_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n275_), .A2(new_n276_), .A3(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n235_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT99), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(KEYINPUT22), .B(G169gat), .Z(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT97), .B1(new_n285_), .B2(G176gat), .ZN(new_n286_));
  INV_X1    g085(.A(G169gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n286_), .B1(new_n287_), .B2(new_n209_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n205_), .B1(G183gat), .B2(G190gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT98), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n205_), .B(KEYINPUT98), .C1(G183gat), .C2(G190gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(KEYINPUT97), .A2(G169gat), .A3(G176gat), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n288_), .A2(new_n291_), .A3(new_n292_), .A4(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT100), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT96), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n226_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n226_), .A2(new_n296_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(new_n232_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n213_), .A2(new_n218_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT25), .B(G183gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT26), .B(G190gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n299_), .A2(new_n205_), .A3(new_n300_), .A4(new_n303_), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n294_), .A2(new_n295_), .A3(new_n280_), .A4(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n235_), .A2(KEYINPUT99), .A3(new_n281_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n284_), .A2(KEYINPUT20), .A3(new_n305_), .A4(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n294_), .A2(new_n304_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n295_), .B1(new_n309_), .B2(new_n280_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n269_), .B1(new_n307_), .B2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n281_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n235_), .A2(new_n281_), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n312_), .A2(new_n313_), .A3(KEYINPUT20), .A4(new_n268_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT18), .B(G64gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(G92gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G8gat), .B(G36gat), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n317_), .B(new_n318_), .Z(new_n319_));
  NAND2_X1  g118(.A1(new_n315_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n319_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n311_), .A2(new_n314_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT0), .B(G57gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(G85gat), .ZN(new_n325_));
  XOR2_X1   g124(.A(G1gat), .B(G29gat), .Z(new_n326_));
  XOR2_X1   g125(.A(new_n325_), .B(new_n326_), .Z(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G225gat), .A2(G233gat), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT101), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G155gat), .A2(G162gat), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333_));
  OR3_X1    g132(.A1(new_n332_), .A2(new_n333_), .A3(KEYINPUT1), .ZN(new_n334_));
  NOR2_X1   g133(.A1(G141gat), .A2(G148gat), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  AOI22_X1  g135(.A1(new_n332_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n334_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT87), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT86), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n339_), .B1(new_n340_), .B2(KEYINPUT3), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(new_n335_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G141gat), .A2(G148gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT2), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT2), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n345_), .A2(G141gat), .A3(G148gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  OAI221_X1 g146(.A(new_n339_), .B1(G141gat), .B2(G148gat), .C1(new_n340_), .C2(KEYINPUT3), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n339_), .A2(KEYINPUT3), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n342_), .A2(new_n347_), .A3(new_n348_), .A4(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT89), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT88), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n352_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n353_));
  OR2_X1    g152(.A1(G155gat), .A2(G162gat), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n354_), .A2(KEYINPUT88), .A3(new_n331_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n350_), .A2(new_n351_), .A3(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n351_), .B1(new_n350_), .B2(new_n356_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n330_), .B(new_n338_), .C1(new_n357_), .C2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n257_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n350_), .A2(new_n356_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT89), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n350_), .A2(new_n351_), .A3(new_n356_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n365_), .A2(new_n330_), .A3(new_n338_), .A4(new_n257_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n361_), .A2(new_n366_), .A3(KEYINPUT4), .ZN(new_n367_));
  INV_X1    g166(.A(new_n338_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n368_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n369_));
  OR3_X1    g168(.A1(new_n369_), .A2(KEYINPUT4), .A3(new_n257_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n329_), .B1(new_n367_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n329_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n372_), .B1(new_n361_), .B2(new_n366_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n328_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT33), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n367_), .A2(new_n329_), .A3(new_n370_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n361_), .A2(new_n366_), .A3(new_n372_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(new_n327_), .A3(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n375_), .B1(new_n374_), .B2(new_n379_), .ZN(new_n380_));
  NOR3_X1   g179(.A1(new_n323_), .A2(new_n376_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n371_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n373_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(new_n327_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n374_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT32), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n315_), .B1(new_n386_), .B2(new_n321_), .ZN(new_n387_));
  OR2_X1    g186(.A1(new_n308_), .A2(KEYINPUT102), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n308_), .A2(KEYINPUT102), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(new_n280_), .A3(new_n389_), .ZN(new_n390_));
  AND3_X1   g189(.A1(new_n284_), .A2(KEYINPUT20), .A3(new_n306_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n269_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  AND4_X1   g191(.A1(KEYINPUT20), .A2(new_n312_), .A3(new_n269_), .A4(new_n313_), .ZN(new_n393_));
  OAI211_X1 g192(.A(KEYINPUT32), .B(new_n319_), .C1(new_n392_), .C2(new_n393_), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n385_), .A2(new_n387_), .A3(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n266_), .B1(new_n381_), .B2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G22gat), .B(G50gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  XOR2_X1   g197(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT29), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n400_), .B1(new_n369_), .B2(new_n401_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n401_), .B(new_n338_), .C1(new_n357_), .C2(new_n358_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n403_), .A2(new_n399_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n398_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n369_), .A2(new_n401_), .A3(new_n400_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n403_), .A2(new_n399_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(new_n407_), .A3(new_n397_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n405_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT94), .ZN(new_n411_));
  XOR2_X1   g210(.A(G78gat), .B(G106gat), .Z(new_n412_));
  OAI21_X1  g211(.A(new_n281_), .B1(new_n369_), .B2(new_n401_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G228gat), .A2(G233gat), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT92), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n413_), .A2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n414_), .B(KEYINPUT92), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n281_), .B(new_n419_), .C1(new_n369_), .C2(new_n401_), .ZN(new_n420_));
  AOI211_X1 g219(.A(new_n411_), .B(new_n412_), .C1(new_n417_), .C2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n338_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n280_), .B1(new_n422_), .B2(KEYINPUT29), .ZN(new_n423_));
  INV_X1    g222(.A(new_n416_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n420_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n412_), .ZN(new_n426_));
  AOI21_X1  g225(.A(KEYINPUT94), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n421_), .A2(new_n427_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n420_), .B(new_n412_), .C1(new_n423_), .C2(new_n424_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT93), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n417_), .A2(KEYINPUT93), .A3(new_n412_), .A4(new_n420_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n410_), .B1(new_n428_), .B2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n429_), .A2(new_n408_), .A3(new_n405_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n412_), .B1(new_n417_), .B2(new_n420_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT95), .B1(new_n434_), .B2(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n423_), .A2(new_n424_), .ZN(new_n439_));
  AOI211_X1 g238(.A(new_n280_), .B(new_n418_), .C1(new_n422_), .C2(KEYINPUT29), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n426_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n411_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n425_), .A2(KEYINPUT94), .A3(new_n426_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n442_), .A2(new_n431_), .A3(new_n432_), .A4(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n409_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT95), .ZN(new_n446_));
  INV_X1    g245(.A(new_n437_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n438_), .A2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n396_), .A2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT104), .B(KEYINPUT27), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n323_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n321_), .A2(KEYINPUT103), .ZN(new_n453_));
  OR2_X1    g252(.A1(new_n321_), .A2(KEYINPUT103), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n453_), .B(new_n454_), .C1(new_n392_), .C2(new_n393_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n455_), .A2(KEYINPUT27), .A3(new_n320_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n452_), .A2(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n446_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n458_));
  AOI211_X1 g257(.A(KEYINPUT95), .B(new_n437_), .C1(new_n444_), .C2(new_n409_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n266_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n264_), .A2(new_n265_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n438_), .A2(new_n448_), .A3(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n457_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n385_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n450_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G57gat), .B(G64gat), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n466_), .A2(KEYINPUT11), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(KEYINPUT11), .ZN(new_n468_));
  XOR2_X1   g267(.A(G71gat), .B(G78gat), .Z(new_n469_));
  NAND3_X1  g268(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  OR2_X1    g269(.A1(new_n468_), .A2(new_n469_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G231gat), .A2(G233gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(G15gat), .ZN(new_n475_));
  INV_X1    g274(.A(G22gat), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n476_), .A2(KEYINPUT75), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(KEYINPUT75), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n475_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT75), .B(G22gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(G15gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G1gat), .A2(G8gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT14), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n479_), .A2(new_n481_), .A3(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(G1gat), .A2(G8gat), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT76), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n486_), .A2(new_n487_), .A3(new_n482_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n482_), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT76), .B1(new_n489_), .B2(new_n485_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n484_), .B(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n474_), .B(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT17), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT16), .B(G183gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(G211gat), .ZN(new_n497_));
  XOR2_X1   g296(.A(G127gat), .B(G155gat), .Z(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  OR3_X1    g298(.A1(new_n494_), .A2(new_n495_), .A3(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(KEYINPUT17), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n494_), .A2(new_n501_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G190gat), .B(G218gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(G134gat), .ZN(new_n506_));
  INV_X1    g305(.A(G162gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n508_), .A2(KEYINPUT36), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G232gat), .A2(G233gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT34), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G29gat), .A2(G36gat), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(G29gat), .A2(G36gat), .ZN(new_n515_));
  OAI21_X1  g314(.A(G43gat), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(G29gat), .ZN(new_n517_));
  INV_X1    g316(.A(G36gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(G43gat), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n519_), .A2(new_n520_), .A3(new_n513_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n516_), .A2(G50gat), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(G50gat), .B1(new_n516_), .B2(new_n521_), .ZN(new_n524_));
  OAI21_X1  g323(.A(KEYINPUT73), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n524_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT73), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n526_), .A2(new_n527_), .A3(new_n522_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n525_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT15), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n525_), .A2(new_n528_), .A3(KEYINPUT15), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT7), .ZN(new_n533_));
  INV_X1    g332(.A(G99gat), .ZN(new_n534_));
  INV_X1    g333(.A(G106gat), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n533_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G99gat), .A2(G106gat), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT6), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n540_));
  NAND3_X1  g339(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n536_), .A2(new_n539_), .A3(new_n540_), .A4(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(G85gat), .ZN(new_n543_));
  INV_X1    g342(.A(G92gat), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G85gat), .A2(G92gat), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n542_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT8), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT69), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT67), .ZN(new_n551_));
  AND3_X1   g350(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n552_));
  AOI21_X1  g351(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n551_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n539_), .A2(KEYINPUT67), .A3(new_n541_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n536_), .A2(new_n540_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(KEYINPUT68), .B(KEYINPUT8), .Z(new_n559_));
  NAND3_X1  g358(.A1(new_n558_), .A2(new_n547_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT69), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n548_), .A2(new_n561_), .A3(KEYINPUT8), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n550_), .A2(new_n560_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT9), .ZN(new_n564_));
  AND3_X1   g363(.A1(new_n546_), .A2(KEYINPUT65), .A3(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n564_), .B1(new_n546_), .B2(KEYINPUT65), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(new_n545_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT66), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT10), .B(G99gat), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n570_), .A2(KEYINPUT64), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(KEYINPUT64), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n535_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT66), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n567_), .A2(new_n574_), .A3(new_n545_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n569_), .A2(new_n573_), .A3(new_n556_), .A4(new_n575_), .ZN(new_n576_));
  AOI22_X1  g375(.A1(new_n531_), .A2(new_n532_), .B1(new_n563_), .B2(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n523_), .A2(new_n524_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n563_), .A2(new_n578_), .A3(new_n576_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  OAI211_X1 g379(.A(KEYINPUT35), .B(new_n512_), .C1(new_n577_), .C2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n563_), .A2(new_n576_), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n525_), .A2(new_n528_), .A3(KEYINPUT15), .ZN(new_n583_));
  AOI21_X1  g382(.A(KEYINPUT15), .B1(new_n525_), .B2(new_n528_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n582_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n512_), .A2(KEYINPUT35), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n512_), .A2(KEYINPUT35), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n585_), .A2(new_n579_), .A3(new_n586_), .A4(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n508_), .B1(new_n581_), .B2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT36), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n510_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n581_), .A2(new_n588_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT74), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n591_), .A2(new_n594_), .ZN(new_n595_));
  OAI211_X1 g394(.A(new_n593_), .B(new_n510_), .C1(new_n590_), .C2(new_n589_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT37), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n465_), .A2(new_n504_), .A3(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n563_), .A2(new_n472_), .A3(new_n576_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G230gat), .A2(G233gat), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT70), .ZN(new_n603_));
  INV_X1    g402(.A(new_n472_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n582_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT12), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n582_), .A2(KEYINPUT12), .A3(new_n604_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT70), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n600_), .A2(new_n609_), .A3(new_n601_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n603_), .A2(new_n607_), .A3(new_n608_), .A4(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n601_), .B1(new_n605_), .B2(new_n600_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(G120gat), .B(G148gat), .Z(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(G204gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT5), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(new_n209_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n611_), .A2(new_n613_), .A3(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT71), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT71), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n611_), .A2(new_n620_), .A3(new_n613_), .A4(new_n617_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n611_), .A2(new_n613_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n617_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n622_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n600_), .A2(new_n609_), .A3(new_n601_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n609_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(KEYINPUT12), .B1(new_n582_), .B2(new_n604_), .ZN(new_n631_));
  AOI211_X1 g430(.A(new_n606_), .B(new_n472_), .C1(new_n563_), .C2(new_n576_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n612_), .B1(new_n630_), .B2(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n620_), .B1(new_n634_), .B2(new_n617_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n621_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n625_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  XOR2_X1   g437(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n639_));
  OAI21_X1  g438(.A(new_n627_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n578_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n493_), .A2(new_n641_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n484_), .A2(new_n491_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n484_), .A2(new_n491_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n578_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT77), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT77), .B1(new_n492_), .B2(new_n578_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n642_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(G229gat), .A2(G233gat), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n493_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n645_), .A2(new_n646_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n492_), .A2(KEYINPUT77), .A3(new_n578_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n653_), .A2(new_n656_), .A3(new_n650_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n652_), .A2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(G113gat), .B(G141gat), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(new_n287_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(new_n271_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n662_), .A2(KEYINPUT78), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n658_), .B(new_n663_), .Z(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT79), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT79), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n664_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n640_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n599_), .A2(new_n671_), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n672_), .A2(G1gat), .A3(new_n464_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n465_), .A2(new_n597_), .A3(new_n504_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n640_), .A2(new_n664_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n676_), .A2(new_n385_), .A3(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(G1gat), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n675_), .A2(new_n680_), .ZN(G1324gat));
  INV_X1    g480(.A(new_n457_), .ZN(new_n682_));
  OR3_X1    g481(.A1(new_n672_), .A2(G8gat), .A3(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n676_), .A2(new_n678_), .A3(new_n457_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT39), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n684_), .A2(new_n685_), .A3(G8gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n684_), .B2(G8gat), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n683_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g488(.A1(new_n676_), .A2(new_n678_), .A3(new_n461_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(G15gat), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n691_), .A2(KEYINPUT106), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(KEYINPUT106), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT41), .ZN(new_n694_));
  OR3_X1    g493(.A1(new_n692_), .A2(new_n693_), .A3(new_n694_), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n599_), .A2(new_n475_), .A3(new_n461_), .A4(new_n671_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n694_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n695_), .A2(new_n696_), .A3(new_n697_), .ZN(G1326gat));
  NAND3_X1  g497(.A1(new_n676_), .A2(new_n678_), .A3(new_n449_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n699_), .A2(new_n700_), .A3(G22gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n699_), .B2(G22gat), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n449_), .A2(new_n476_), .ZN(new_n703_));
  OAI22_X1  g502(.A1(new_n701_), .A2(new_n702_), .B1(new_n672_), .B2(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT107), .ZN(G1327gat));
  NAND2_X1  g504(.A1(KEYINPUT108), .A2(KEYINPUT43), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(KEYINPUT108), .A2(KEYINPUT43), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n595_), .A2(new_n596_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT37), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n709_), .B1(new_n465_), .B2(new_n711_), .ZN(new_n712_));
  AOI211_X1 g511(.A(new_n385_), .B(new_n457_), .C1(new_n460_), .C2(new_n462_), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n598_), .B(new_n707_), .C1(new_n713_), .C2(new_n450_), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n712_), .A2(new_n678_), .A3(new_n714_), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n715_), .A2(KEYINPUT109), .A3(KEYINPUT44), .A4(new_n504_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n712_), .A2(new_n678_), .A3(new_n504_), .A4(new_n714_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n717_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n716_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n718_), .A2(new_n719_), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n721_), .A2(G29gat), .A3(new_n385_), .A4(new_n722_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n465_), .A2(new_n710_), .A3(new_n503_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(new_n671_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n517_), .B1(new_n725_), .B2(new_n464_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n723_), .A2(new_n726_), .ZN(G1328gat));
  INV_X1    g526(.A(KEYINPUT46), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n682_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n518_), .B1(new_n721_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n725_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n731_), .A2(KEYINPUT45), .A3(new_n518_), .A4(new_n457_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n724_), .A2(new_n518_), .A3(new_n671_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n734_), .B2(new_n682_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n732_), .A2(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n728_), .B1(new_n730_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n736_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n729_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n720_), .B2(new_n716_), .ZN(new_n740_));
  OAI211_X1 g539(.A(KEYINPUT46), .B(new_n738_), .C1(new_n740_), .C2(new_n518_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n737_), .A2(new_n741_), .ZN(G1329gat));
  NOR2_X1   g541(.A1(new_n266_), .A2(new_n520_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  AOI221_X4 g543(.A(new_n744_), .B1(new_n719_), .B2(new_n718_), .C1(new_n716_), .C2(new_n720_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n725_), .A2(new_n266_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n746_), .A2(G43gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(KEYINPUT47), .B1(new_n745_), .B2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n721_), .A2(new_n722_), .A3(new_n743_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT47), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n749_), .B(new_n750_), .C1(G43gat), .C2(new_n746_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n748_), .A2(new_n751_), .ZN(G1330gat));
  AND3_X1   g551(.A1(new_n721_), .A2(new_n449_), .A3(new_n722_), .ZN(new_n753_));
  INV_X1    g552(.A(G50gat), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n449_), .A2(new_n754_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT110), .Z(new_n756_));
  OAI22_X1  g555(.A1(new_n753_), .A2(new_n754_), .B1(new_n725_), .B2(new_n756_), .ZN(G1331gat));
  NOR2_X1   g556(.A1(new_n640_), .A2(new_n664_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n599_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(G57gat), .B1(new_n760_), .B2(new_n385_), .ZN(new_n761_));
  OAI21_X1  g560(.A(G57gat), .B1(new_n464_), .B2(KEYINPUT111), .ZN(new_n762_));
  INV_X1    g561(.A(new_n640_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n676_), .A2(new_n763_), .A3(new_n666_), .A4(new_n668_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(KEYINPUT111), .A2(G57gat), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n761_), .B1(new_n762_), .B2(new_n766_), .ZN(G1332gat));
  OAI21_X1  g566(.A(G64gat), .B1(new_n764_), .B2(new_n682_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT48), .ZN(new_n769_));
  OR2_X1    g568(.A1(new_n682_), .A2(G64gat), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(new_n759_), .B2(new_n770_), .ZN(G1333gat));
  NAND3_X1  g570(.A1(new_n760_), .A2(new_n237_), .A3(new_n461_), .ZN(new_n772_));
  OAI21_X1  g571(.A(G71gat), .B1(new_n764_), .B2(new_n266_), .ZN(new_n773_));
  OR2_X1    g572(.A1(new_n773_), .A2(KEYINPUT112), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(KEYINPUT112), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n774_), .A2(KEYINPUT49), .A3(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT49), .B1(new_n774_), .B2(new_n775_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n772_), .B1(new_n776_), .B2(new_n777_), .ZN(G1334gat));
  INV_X1    g577(.A(new_n449_), .ZN(new_n779_));
  OR3_X1    g578(.A1(new_n759_), .A2(G78gat), .A3(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(G78gat), .B1(new_n764_), .B2(new_n779_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n781_), .A2(KEYINPUT50), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n783_), .B(G78gat), .C1(new_n764_), .C2(new_n779_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n780_), .B1(new_n782_), .B2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT113), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n780_), .B(new_n788_), .C1(new_n782_), .C2(new_n785_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(G1335gat));
  AND2_X1   g589(.A1(new_n724_), .A2(new_n758_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n791_), .A2(new_n543_), .A3(new_n385_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n712_), .A2(new_n504_), .A3(new_n714_), .A4(new_n758_), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n793_), .A2(KEYINPUT114), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(KEYINPUT114), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n464_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n792_), .B1(new_n796_), .B2(new_n543_), .ZN(G1336gat));
  NAND3_X1  g596(.A1(new_n791_), .A2(new_n544_), .A3(new_n457_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n682_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(new_n544_), .ZN(G1337gat));
  OAI211_X1 g599(.A(new_n791_), .B(new_n461_), .C1(new_n572_), .C2(new_n571_), .ZN(new_n801_));
  OAI21_X1  g600(.A(G99gat), .B1(new_n793_), .B2(new_n266_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g603(.A(G106gat), .B1(new_n793_), .B2(new_n779_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT52), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n807_), .B(G106gat), .C1(new_n793_), .C2(new_n779_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n791_), .A2(new_n535_), .A3(new_n449_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n809_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n810_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n812_), .A2(new_n813_), .ZN(G1339gat));
  AND3_X1   g613(.A1(new_n666_), .A2(new_n503_), .A3(new_n668_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n711_), .A2(new_n815_), .A3(new_n640_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT54), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT119), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n611_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n607_), .A2(new_n600_), .A3(new_n608_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n821_), .A2(G230gat), .A3(G233gat), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n633_), .A2(KEYINPUT55), .A3(new_n603_), .A4(new_n610_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n820_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n624_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT56), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n824_), .A2(KEYINPUT56), .A3(new_n624_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n827_), .A2(KEYINPUT118), .A3(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n649_), .A2(new_n650_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n653_), .A2(new_n656_), .A3(new_n651_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n662_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n661_), .B1(new_n652_), .B2(new_n657_), .ZN(new_n833_));
  OAI21_X1  g632(.A(KEYINPUT117), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n831_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n651_), .B1(new_n656_), .B2(new_n642_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n661_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n653_), .A2(new_n656_), .A3(new_n650_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n650_), .B1(new_n656_), .B2(new_n642_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n662_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n837_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n622_), .A2(new_n834_), .A3(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT118), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n825_), .A2(new_n844_), .A3(new_n826_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n829_), .A2(new_n843_), .A3(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT58), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n829_), .A2(KEYINPUT58), .A3(new_n843_), .A4(new_n845_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n598_), .A3(new_n849_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n834_), .A2(new_n842_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n637_), .A2(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n824_), .A2(new_n624_), .A3(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n854_), .A2(new_n664_), .A3(new_n622_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n853_), .B1(new_n824_), .B2(new_n624_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n852_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT57), .B1(new_n857_), .B2(new_n710_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n857_), .A2(KEYINPUT57), .A3(new_n710_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n850_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n818_), .B1(new_n861_), .B2(new_n504_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863_));
  INV_X1    g662(.A(new_n853_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n825_), .A2(new_n864_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n865_), .A2(new_n664_), .A3(new_n622_), .A4(new_n854_), .ZN(new_n866_));
  AOI211_X1 g665(.A(new_n863_), .B(new_n597_), .C1(new_n866_), .C2(new_n852_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(new_n858_), .ZN(new_n868_));
  AOI211_X1 g667(.A(KEYINPUT119), .B(new_n503_), .C1(new_n868_), .C2(new_n850_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n817_), .B1(new_n862_), .B2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT59), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n462_), .A2(new_n464_), .A3(new_n457_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n870_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n861_), .A2(new_n504_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n817_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n872_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT59), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n873_), .A2(G113gat), .A3(new_n669_), .A4(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n251_), .B1(new_n876_), .B2(new_n665_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1340gat));
  INV_X1    g679(.A(G120gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n881_), .B1(new_n640_), .B2(KEYINPUT60), .ZN(new_n882_));
  OR2_X1    g681(.A1(new_n881_), .A2(KEYINPUT60), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n875_), .A2(new_n872_), .A3(new_n882_), .A4(new_n883_), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n873_), .A2(new_n763_), .A3(new_n877_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(new_n881_), .ZN(G1341gat));
  NAND4_X1  g685(.A1(new_n873_), .A2(G127gat), .A3(new_n503_), .A4(new_n877_), .ZN(new_n887_));
  INV_X1    g686(.A(G127gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n888_), .B1(new_n876_), .B2(new_n504_), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n887_), .A2(new_n889_), .ZN(G1342gat));
  NAND4_X1  g689(.A1(new_n873_), .A2(G134gat), .A3(new_n598_), .A4(new_n877_), .ZN(new_n891_));
  INV_X1    g690(.A(G134gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n892_), .B1(new_n876_), .B2(new_n710_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n891_), .A2(new_n893_), .ZN(G1343gat));
  AOI21_X1  g693(.A(new_n460_), .B1(new_n874_), .B2(new_n817_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n457_), .A2(new_n464_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n664_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n763_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g701(.A1(new_n897_), .A2(new_n504_), .ZN(new_n903_));
  XOR2_X1   g702(.A(KEYINPUT61), .B(G155gat), .Z(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1346gat));
  NOR3_X1   g704(.A1(new_n897_), .A2(new_n507_), .A3(new_n711_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n898_), .A2(new_n597_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n507_), .B2(new_n907_), .ZN(G1347gat));
  NOR3_X1   g707(.A1(new_n682_), .A2(new_n385_), .A3(new_n266_), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n870_), .A2(new_n664_), .A3(new_n779_), .A4(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(G169gat), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n910_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n914_));
  OAI211_X1 g713(.A(new_n913_), .B(new_n914_), .C1(new_n285_), .C2(new_n910_), .ZN(G1348gat));
  NAND4_X1  g714(.A1(new_n870_), .A2(new_n763_), .A3(new_n779_), .A4(new_n909_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n209_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n449_), .B1(new_n874_), .B2(new_n817_), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n918_), .A2(G176gat), .A3(new_n763_), .A4(new_n909_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(KEYINPUT120), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT120), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n917_), .A2(new_n922_), .A3(new_n919_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n923_), .ZN(G1349gat));
  NAND2_X1  g723(.A1(new_n909_), .A2(new_n503_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n925_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n206_), .B1(new_n918_), .B2(new_n926_), .ZN(new_n927_));
  AND2_X1   g726(.A1(new_n870_), .A2(new_n779_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n925_), .A2(new_n301_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n927_), .B1(new_n928_), .B2(new_n929_), .ZN(G1350gat));
  NAND3_X1  g729(.A1(new_n928_), .A2(new_n598_), .A3(new_n909_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(G190gat), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n928_), .A2(new_n302_), .A3(new_n909_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n710_), .B2(new_n933_), .ZN(G1351gat));
  INV_X1    g733(.A(new_n460_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n682_), .A2(new_n385_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT54), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n816_), .B(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n503_), .B1(new_n868_), .B2(new_n850_), .ZN(new_n939_));
  OAI211_X1 g738(.A(new_n935_), .B(new_n936_), .C1(new_n938_), .C2(new_n939_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n940_), .A2(new_n665_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(KEYINPUT121), .B(G197gat), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n941_), .B(new_n942_), .ZN(G1352gat));
  INV_X1    g742(.A(new_n940_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(new_n763_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g745(.A(new_n504_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n947_));
  OR2_X1    g746(.A1(new_n947_), .A2(KEYINPUT122), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(KEYINPUT122), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n944_), .A2(new_n948_), .A3(new_n949_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n950_), .A2(KEYINPUT123), .ZN(new_n951_));
  NOR2_X1   g750(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n952_));
  INV_X1    g751(.A(KEYINPUT123), .ZN(new_n953_));
  NAND4_X1  g752(.A1(new_n944_), .A2(new_n953_), .A3(new_n948_), .A4(new_n949_), .ZN(new_n954_));
  AND3_X1   g753(.A1(new_n951_), .A2(new_n952_), .A3(new_n954_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n952_), .B1(new_n951_), .B2(new_n954_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n955_), .A2(new_n956_), .ZN(G1354gat));
  XNOR2_X1  g756(.A(KEYINPUT125), .B(G218gat), .ZN(new_n958_));
  INV_X1    g757(.A(new_n958_), .ZN(new_n959_));
  NOR3_X1   g758(.A1(new_n940_), .A2(new_n711_), .A3(new_n959_), .ZN(new_n960_));
  INV_X1    g759(.A(KEYINPUT124), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n961_), .B1(new_n940_), .B2(new_n710_), .ZN(new_n962_));
  NAND4_X1  g761(.A1(new_n895_), .A2(KEYINPUT124), .A3(new_n597_), .A4(new_n936_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n962_), .A2(new_n963_), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n960_), .B1(new_n964_), .B2(new_n959_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n965_), .A2(KEYINPUT126), .ZN(new_n966_));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n958_), .B1(new_n962_), .B2(new_n963_), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n967_), .B1(new_n968_), .B2(new_n960_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n966_), .A2(new_n969_), .ZN(G1355gat));
endmodule


