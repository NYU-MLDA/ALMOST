//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 1 0 1 0 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 1 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n825_, new_n826_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n835_, new_n836_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n869_, new_n870_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_;
  NOR2_X1   g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT7), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n205_));
  AND2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT65), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT6), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n204_), .A2(new_n205_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n207_), .A2(new_n209_), .A3(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(G85gat), .B(G92gat), .Z(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT66), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n213_), .A2(new_n217_), .A3(new_n214_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(KEYINPUT8), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n206_), .A2(new_n209_), .ZN(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT8), .B1(new_n220_), .B2(KEYINPUT64), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n221_), .B(new_n214_), .C1(KEYINPUT64), .C2(new_n220_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n219_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n209_), .ZN(new_n224_));
  INV_X1    g023(.A(G85gat), .ZN(new_n225_));
  INV_X1    g024(.A(G92gat), .ZN(new_n226_));
  NOR3_X1   g025(.A1(new_n225_), .A2(new_n226_), .A3(KEYINPUT9), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n224_), .A2(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(KEYINPUT10), .B(G99gat), .Z(new_n229_));
  INV_X1    g028(.A(G106gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n214_), .A2(KEYINPUT9), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n228_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n223_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT67), .ZN(new_n235_));
  INV_X1    g034(.A(new_n233_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n236_), .B1(new_n219_), .B2(new_n222_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n235_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G29gat), .B(G36gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT69), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(G43gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(G50gat), .ZN(new_n244_));
  INV_X1    g043(.A(G50gat), .ZN(new_n245_));
  INV_X1    g044(.A(G43gat), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n242_), .A2(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n242_), .A2(new_n246_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n245_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n244_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n240_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n244_), .A2(KEYINPUT15), .A3(new_n249_), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT15), .B1(new_n244_), .B2(new_n249_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n253_), .B1(new_n256_), .B2(new_n237_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n256_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(KEYINPUT70), .A3(new_n234_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n252_), .A2(new_n257_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G232gat), .A2(G233gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT34), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT35), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n260_), .A2(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n262_), .A2(KEYINPUT35), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n252_), .B(new_n267_), .C1(new_n256_), .C2(new_n237_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G190gat), .B(G218gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(G134gat), .ZN(new_n271_));
  INV_X1    g070(.A(G162gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT36), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n273_), .A2(new_n274_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n269_), .A2(new_n275_), .A3(new_n277_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n265_), .A2(new_n274_), .A3(new_n273_), .A4(new_n268_), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n278_), .A2(KEYINPUT37), .A3(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(KEYINPUT37), .B1(new_n278_), .B2(new_n279_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT71), .B(G8gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(G1gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT14), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G15gat), .B(G22gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(G1gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(G8gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n286_), .B(G1gat), .ZN(new_n290_));
  INV_X1    g089(.A(G8gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  XOR2_X1   g093(.A(G71gat), .B(G78gat), .Z(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT11), .ZN(new_n297_));
  XOR2_X1   g096(.A(G57gat), .B(G64gat), .Z(new_n298_));
  OR3_X1    g097(.A1(new_n296_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n297_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n296_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n299_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G231gat), .A2(G233gat), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n302_), .B(new_n303_), .Z(new_n304_));
  XNOR2_X1  g103(.A(new_n294_), .B(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G183gat), .B(G211gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(G155gat), .ZN(new_n308_));
  XOR2_X1   g107(.A(KEYINPUT73), .B(KEYINPUT16), .Z(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT74), .B(G127gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n312_), .A2(KEYINPUT72), .A3(KEYINPUT17), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n306_), .A2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n313_), .B1(KEYINPUT17), .B2(new_n312_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n305_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n317_), .B(KEYINPUT75), .Z(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NOR3_X1   g118(.A1(new_n280_), .A2(new_n281_), .A3(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n320_), .B(KEYINPUT76), .Z(new_n321_));
  NOR2_X1   g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT79), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT24), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G169gat), .A2(G176gat), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n327_), .B(KEYINPUT80), .Z(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G183gat), .A2(G190gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT23), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n324_), .A2(new_n325_), .ZN(new_n332_));
  INV_X1    g131(.A(G183gat), .ZN(new_n333_));
  OR3_X1    g132(.A1(new_n333_), .A2(KEYINPUT78), .A3(KEYINPUT25), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT26), .B(G190gat), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT25), .B1(new_n333_), .B2(KEYINPUT78), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n334_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n329_), .A2(new_n331_), .A3(new_n332_), .A4(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n331_), .B1(G183gat), .B2(G190gat), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n339_), .A2(new_n328_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT22), .B(G169gat), .ZN(new_n341_));
  INV_X1    g140(.A(G176gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n338_), .A2(new_n344_), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n345_), .B(KEYINPUT81), .Z(new_n346_));
  XOR2_X1   g145(.A(new_n346_), .B(KEYINPUT30), .Z(new_n347_));
  NOR2_X1   g146(.A1(new_n347_), .A2(KEYINPUT82), .ZN(new_n348_));
  XOR2_X1   g147(.A(G15gat), .B(G43gat), .Z(new_n349_));
  XNOR2_X1  g148(.A(G71gat), .B(G99gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G227gat), .A2(G233gat), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n351_), .B(new_n352_), .Z(new_n353_));
  XNOR2_X1  g152(.A(new_n346_), .B(KEYINPUT30), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT82), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n353_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  OR2_X1    g155(.A1(new_n348_), .A2(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(G127gat), .A2(G134gat), .ZN(new_n358_));
  AND2_X1   g157(.A1(G127gat), .A2(G134gat), .ZN(new_n359_));
  AND2_X1   g158(.A1(G113gat), .A2(G120gat), .ZN(new_n360_));
  NOR2_X1   g159(.A1(G113gat), .A2(G120gat), .ZN(new_n361_));
  OAI22_X1  g160(.A1(new_n358_), .A2(new_n359_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT84), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G127gat), .B(G134gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G113gat), .B(G120gat), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(new_n366_), .A3(KEYINPUT84), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n364_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT85), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n369_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n359_), .A2(new_n358_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n360_), .A2(new_n361_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(new_n372_), .A3(KEYINPUT85), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n370_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT86), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n368_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n375_), .B1(new_n368_), .B2(new_n374_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n378_), .B(KEYINPUT31), .Z(new_n379_));
  NOR2_X1   g178(.A1(new_n379_), .A2(KEYINPUT83), .ZN(new_n380_));
  NOR3_X1   g179(.A1(new_n347_), .A2(KEYINPUT82), .A3(new_n353_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n357_), .A2(new_n380_), .A3(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n348_), .A2(new_n356_), .ZN(new_n384_));
  OAI22_X1  g183(.A1(new_n384_), .A2(new_n381_), .B1(KEYINPUT83), .B2(new_n379_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G8gat), .B(G36gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT18), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(G64gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(new_n226_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G211gat), .B(G218gat), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT91), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT90), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  XOR2_X1   g195(.A(G197gat), .B(G204gat), .Z(new_n397_));
  NAND3_X1  g196(.A1(new_n396_), .A2(KEYINPUT21), .A3(new_n397_), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n397_), .A2(KEYINPUT21), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(KEYINPUT21), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n394_), .A2(new_n395_), .A3(new_n399_), .A4(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n398_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n345_), .A2(new_n402_), .ZN(new_n403_));
  XOR2_X1   g202(.A(new_n341_), .B(KEYINPUT95), .Z(new_n404_));
  OAI21_X1  g203(.A(new_n340_), .B1(G176gat), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n326_), .A2(new_n327_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT25), .B(G183gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n335_), .A2(new_n407_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n406_), .A2(new_n331_), .A3(new_n408_), .A4(new_n332_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n405_), .A2(new_n409_), .A3(new_n398_), .A4(new_n401_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G226gat), .A2(G233gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(KEYINPUT19), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n403_), .A2(KEYINPUT20), .A3(new_n410_), .A4(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT20), .B1(new_n345_), .B2(new_n402_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT94), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n405_), .A2(new_n409_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n402_), .ZN(new_n420_));
  OAI211_X1 g219(.A(KEYINPUT94), .B(KEYINPUT20), .C1(new_n345_), .C2(new_n402_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n418_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  AOI211_X1 g221(.A(new_n391_), .B(new_n415_), .C1(new_n422_), .C2(new_n412_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(KEYINPUT98), .A2(KEYINPUT20), .ZN(new_n425_));
  OR2_X1    g224(.A1(KEYINPUT98), .A2(KEYINPUT20), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n403_), .A2(new_n410_), .A3(new_n425_), .A4(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(KEYINPUT99), .A3(new_n412_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n428_), .B1(new_n422_), .B2(new_n412_), .ZN(new_n429_));
  AOI21_X1  g228(.A(KEYINPUT99), .B1(new_n427_), .B2(new_n412_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n391_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n424_), .A2(new_n431_), .A3(KEYINPUT27), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT27), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n422_), .A2(new_n412_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n390_), .B1(new_n434_), .B2(new_n414_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n433_), .B1(new_n435_), .B2(new_n423_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n432_), .A2(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(KEYINPUT87), .B1(G155gat), .B2(G162gat), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT1), .ZN(new_n440_));
  NAND3_X1  g239(.A1(KEYINPUT87), .A2(G155gat), .A3(G162gat), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n439_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n441_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT1), .B1(new_n443_), .B2(new_n438_), .ZN(new_n444_));
  OR2_X1    g243(.A1(G155gat), .A2(G162gat), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n442_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  XOR2_X1   g245(.A(G141gat), .B(G148gat), .Z(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(G141gat), .ZN(new_n449_));
  INV_X1    g248(.A(G148gat), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT88), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n449_), .B(new_n450_), .C1(new_n451_), .C2(KEYINPUT3), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT3), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n453_), .B(KEYINPUT88), .C1(G141gat), .C2(G148gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G141gat), .A2(G148gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT2), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT2), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(G141gat), .A3(G148gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n455_), .A2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n445_), .B1(new_n461_), .B2(KEYINPUT89), .ZN(new_n462_));
  AOI22_X1  g261(.A1(new_n452_), .A2(new_n454_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT89), .ZN(new_n464_));
  OAI22_X1  g263(.A1(new_n463_), .A2(new_n464_), .B1(new_n438_), .B2(new_n443_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n448_), .B1(new_n462_), .B2(new_n465_), .ZN(new_n466_));
  AOI22_X1  g265(.A1(new_n398_), .A2(new_n401_), .B1(new_n466_), .B2(KEYINPUT29), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G228gat), .A2(G233gat), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT92), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n468_), .A2(new_n469_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n467_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G78gat), .B(G106gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(new_n245_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n472_), .A2(new_n474_), .A3(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n477_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n466_), .A2(KEYINPUT29), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT28), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT93), .B(G22gat), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(new_n483_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n480_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n482_), .B(new_n483_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n487_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n437_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G1gat), .B(G29gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(G85gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT0), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(G57gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n371_), .A2(new_n372_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n362_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n448_), .B(new_n496_), .C1(new_n462_), .C2(new_n465_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT96), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n466_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n497_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n499_), .B1(new_n501_), .B2(KEYINPUT96), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G225gat), .A2(G233gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n501_), .A2(KEYINPUT96), .ZN(new_n506_));
  INV_X1    g305(.A(new_n499_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n506_), .A2(KEYINPUT97), .A3(KEYINPUT4), .A4(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n498_), .B1(new_n500_), .B2(new_n497_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT4), .ZN(new_n510_));
  NOR3_X1   g309(.A1(new_n509_), .A2(new_n510_), .A3(new_n499_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT97), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n512_), .B1(new_n500_), .B2(KEYINPUT4), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n508_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n503_), .ZN(new_n515_));
  AOI211_X1 g314(.A(new_n494_), .B(new_n505_), .C1(new_n514_), .C2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n494_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n513_), .B1(new_n502_), .B2(KEYINPUT4), .ZN(new_n518_));
  NOR4_X1   g317(.A1(new_n509_), .A2(new_n512_), .A3(new_n510_), .A4(new_n499_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n515_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n517_), .B1(new_n520_), .B2(new_n504_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n516_), .A2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n386_), .A2(new_n490_), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n520_), .A2(new_n517_), .A3(new_n504_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT33), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n435_), .A2(new_n423_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n514_), .A2(new_n503_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n502_), .A2(new_n515_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(new_n494_), .A3(new_n530_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n520_), .A2(KEYINPUT33), .A3(new_n517_), .A4(new_n504_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n527_), .A2(new_n528_), .A3(new_n531_), .A4(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n390_), .A2(KEYINPUT32), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n434_), .A2(new_n414_), .A3(new_n534_), .ZN(new_n535_));
  OAI211_X1 g334(.A(KEYINPUT32), .B(new_n390_), .C1(new_n429_), .C2(new_n430_), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n535_), .B(new_n536_), .C1(new_n516_), .C2(new_n521_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n533_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n486_), .A2(new_n488_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT100), .ZN(new_n541_));
  INV_X1    g340(.A(new_n522_), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n542_), .A2(new_n437_), .A3(new_n539_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT100), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n538_), .A2(new_n545_), .A3(new_n539_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n541_), .A2(new_n544_), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n386_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n524_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n235_), .A2(new_n239_), .A3(new_n302_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT12), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n302_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n240_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G230gat), .A2(G233gat), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n234_), .A2(KEYINPUT12), .A3(new_n302_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n552_), .A2(new_n554_), .A3(new_n555_), .A4(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n554_), .A2(new_n550_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n557_), .B1(new_n558_), .B2(new_n555_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G120gat), .B(G148gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT5), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(G176gat), .ZN(new_n562_));
  INV_X1    g361(.A(G204gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n559_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n559_), .A2(new_n564_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  XOR2_X1   g366(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT13), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n565_), .B(new_n566_), .C1(KEYINPUT68), .C2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n251_), .A2(new_n293_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT77), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n575_), .B1(new_n258_), .B2(new_n294_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G229gat), .A2(G233gat), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n251_), .A2(new_n293_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n575_), .A2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n578_), .B1(new_n577_), .B2(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(G113gat), .B(G141gat), .Z(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(G169gat), .ZN(new_n583_));
  INV_X1    g382(.A(G197gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n581_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n585_), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n578_), .B(new_n587_), .C1(new_n577_), .C2(new_n580_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n572_), .A2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n549_), .A2(new_n590_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n321_), .A2(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n592_), .A2(new_n287_), .A3(new_n542_), .ZN(new_n593_));
  XOR2_X1   g392(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n275_), .ZN(new_n596_));
  AOI211_X1 g395(.A(new_n596_), .B(new_n276_), .C1(new_n265_), .C2(new_n268_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n279_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n591_), .A2(new_n600_), .A3(new_n317_), .ZN(new_n601_));
  OAI21_X1  g400(.A(G1gat), .B1(new_n601_), .B2(new_n522_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n595_), .A2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT102), .ZN(G1324gat));
  INV_X1    g403(.A(new_n437_), .ZN(new_n605_));
  OAI21_X1  g404(.A(G8gat), .B1(new_n601_), .B2(new_n605_), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n606_), .B(KEYINPUT39), .Z(new_n607_));
  INV_X1    g406(.A(new_n592_), .ZN(new_n608_));
  NOR3_X1   g407(.A1(new_n608_), .A2(new_n282_), .A3(new_n605_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT40), .ZN(G1325gat));
  OAI21_X1  g410(.A(G15gat), .B1(new_n601_), .B2(new_n548_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT103), .Z(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT41), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n548_), .A2(G15gat), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n614_), .B1(new_n608_), .B2(new_n615_), .ZN(G1326gat));
  OAI21_X1  g415(.A(G22gat), .B1(new_n601_), .B2(new_n539_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT42), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n539_), .A2(G22gat), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n619_), .B(KEYINPUT104), .Z(new_n620_));
  OAI21_X1  g419(.A(new_n618_), .B1(new_n608_), .B2(new_n620_), .ZN(G1327gat));
  NOR2_X1   g420(.A1(new_n600_), .A2(new_n318_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n591_), .A2(new_n622_), .ZN(new_n623_));
  OR3_X1    g422(.A1(new_n623_), .A2(G29gat), .A3(new_n522_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT44), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n280_), .A2(new_n281_), .ZN(new_n626_));
  NOR3_X1   g425(.A1(new_n549_), .A2(KEYINPUT43), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT105), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n628_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT37), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n630_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n278_), .A2(KEYINPUT37), .A3(new_n279_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n631_), .A2(KEYINPUT105), .A3(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n629_), .A2(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(KEYINPUT43), .B1(new_n549_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT106), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n545_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n638_));
  AOI211_X1 g437(.A(KEYINPUT100), .B(new_n489_), .C1(new_n533_), .C2(new_n537_), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n638_), .A2(new_n639_), .A3(new_n543_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n523_), .B1(new_n640_), .B2(new_n386_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n280_), .A2(new_n281_), .A3(new_n628_), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT105), .B1(new_n631_), .B2(new_n632_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n641_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n645_), .A2(KEYINPUT106), .A3(KEYINPUT43), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n627_), .B1(new_n637_), .B2(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n590_), .A2(new_n318_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n625_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n627_), .ZN(new_n651_));
  AOI21_X1  g450(.A(KEYINPUT106), .B1(new_n645_), .B2(KEYINPUT43), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT43), .ZN(new_n653_));
  AOI211_X1 g452(.A(new_n636_), .B(new_n653_), .C1(new_n641_), .C2(new_n644_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n651_), .B1(new_n652_), .B2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(KEYINPUT44), .A3(new_n648_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n650_), .A2(new_n656_), .A3(new_n542_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT107), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n657_), .A2(new_n658_), .A3(G29gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n657_), .B2(G29gat), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n624_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT108), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT108), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n663_), .B(new_n624_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(G1328gat));
  NOR3_X1   g464(.A1(new_n623_), .A2(G36gat), .A3(new_n605_), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n666_), .B(KEYINPUT45), .Z(new_n667_));
  AND3_X1   g466(.A1(new_n650_), .A2(new_n656_), .A3(new_n437_), .ZN(new_n668_));
  INV_X1    g467(.A(G36gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n667_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT46), .Z(G1329gat));
  NAND4_X1  g470(.A1(new_n650_), .A2(new_n656_), .A3(G43gat), .A4(new_n386_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n246_), .B1(new_n623_), .B2(new_n548_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g474(.A1(new_n650_), .A2(new_n656_), .A3(G50gat), .A4(new_n489_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n245_), .B1(new_n623_), .B2(new_n539_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1331gat));
  INV_X1    g477(.A(new_n572_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n321_), .A2(new_n679_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT109), .Z(new_n681_));
  INV_X1    g480(.A(new_n589_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n681_), .A2(new_n682_), .A3(new_n641_), .ZN(new_n683_));
  AOI21_X1  g482(.A(G57gat), .B1(new_n683_), .B2(new_n542_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n549_), .A2(new_n589_), .A3(new_n572_), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n685_), .A2(new_n600_), .A3(new_n318_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n542_), .A2(G57gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n684_), .B1(new_n686_), .B2(new_n687_), .ZN(G1332gat));
  INV_X1    g487(.A(G64gat), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n683_), .A2(new_n689_), .A3(new_n437_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n686_), .B2(new_n437_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT48), .Z(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(G1333gat));
  INV_X1    g492(.A(G71gat), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n386_), .A2(new_n694_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT110), .Z(new_n696_));
  NAND2_X1  g495(.A1(new_n683_), .A2(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n694_), .B1(new_n686_), .B2(new_n386_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT49), .Z(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(G1334gat));
  INV_X1    g499(.A(G78gat), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n683_), .A2(new_n701_), .A3(new_n489_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n686_), .B2(new_n489_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT50), .Z(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT111), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n702_), .A2(KEYINPUT111), .A3(new_n704_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1335gat));
  AND2_X1   g508(.A1(new_n685_), .A2(new_n622_), .ZN(new_n710_));
  AOI21_X1  g509(.A(G85gat), .B1(new_n710_), .B2(new_n542_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n572_), .A2(new_n318_), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n655_), .A2(new_n682_), .A3(new_n712_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n522_), .A2(new_n225_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n711_), .B1(new_n713_), .B2(new_n714_), .ZN(G1336gat));
  AOI21_X1  g514(.A(G92gat), .B1(new_n710_), .B2(new_n437_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n605_), .A2(new_n226_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n713_), .B2(new_n717_), .ZN(G1337gat));
  NAND2_X1  g517(.A1(new_n713_), .A2(new_n386_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(G99gat), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT113), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT51), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n710_), .A2(new_n229_), .A3(new_n386_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT112), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n720_), .A2(new_n722_), .A3(new_n724_), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n721_), .A2(KEYINPUT51), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n725_), .B(new_n726_), .ZN(G1338gat));
  NAND3_X1  g526(.A1(new_n710_), .A2(new_n230_), .A3(new_n489_), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n655_), .A2(new_n682_), .A3(new_n489_), .A4(new_n712_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT52), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n729_), .A2(new_n730_), .A3(G106gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n729_), .B2(G106gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n733_), .B(new_n734_), .Z(G1339gat));
  INV_X1    g534(.A(G113gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n386_), .A2(new_n490_), .A3(new_n542_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT57), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT119), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT115), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n557_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT55), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n552_), .A2(new_n554_), .A3(new_n556_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n744_), .A2(G230gat), .A3(G233gat), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT55), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n557_), .A2(new_n741_), .A3(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n743_), .A2(new_n745_), .A3(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT116), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT116), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n743_), .A2(new_n745_), .A3(new_n750_), .A4(new_n747_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n749_), .A2(new_n564_), .A3(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT56), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n753_), .A2(KEYINPUT117), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n565_), .A2(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n682_), .B1(new_n752_), .B2(new_n755_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n749_), .A2(new_n564_), .A3(new_n751_), .A4(new_n754_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n577_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n585_), .B1(new_n580_), .B2(new_n758_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT118), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n576_), .A2(new_n758_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n588_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  AOI22_X1  g563(.A1(new_n756_), .A2(new_n757_), .B1(new_n567_), .B2(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n740_), .B1(new_n765_), .B2(new_n599_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n752_), .A2(new_n755_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n767_), .A2(new_n589_), .A3(new_n757_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n764_), .A2(new_n567_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n740_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n770_), .A2(new_n600_), .A3(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n766_), .A2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n763_), .B1(new_n752_), .B2(KEYINPUT56), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n749_), .A2(new_n753_), .A3(new_n564_), .A4(new_n751_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(new_n565_), .A3(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT58), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n626_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n774_), .A2(KEYINPUT58), .A3(new_n565_), .A4(new_n775_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n778_), .A2(new_n779_), .A3(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n317_), .B1(new_n773_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n320_), .A2(new_n682_), .ZN(new_n783_));
  OR3_X1    g582(.A1(new_n783_), .A2(KEYINPUT54), .A3(new_n679_), .ZN(new_n784_));
  OAI21_X1  g583(.A(KEYINPUT54), .B1(new_n783_), .B2(new_n679_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n738_), .B1(new_n782_), .B2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n736_), .B1(new_n788_), .B2(new_n682_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT120), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  OAI211_X1 g590(.A(KEYINPUT120), .B(new_n736_), .C1(new_n788_), .C2(new_n682_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n318_), .B1(new_n773_), .B2(new_n781_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n794_), .A2(new_n787_), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n795_), .A2(KEYINPUT59), .A3(new_n737_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT121), .B1(new_n788_), .B2(KEYINPUT59), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n765_), .A2(new_n599_), .A3(new_n740_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n771_), .B1(new_n770_), .B2(new_n600_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n781_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n317_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n787_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(KEYINPUT121), .B(KEYINPUT59), .C1(new_n803_), .C2(new_n737_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n796_), .B1(new_n798_), .B2(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n682_), .A2(new_n736_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n793_), .B1(new_n805_), .B2(new_n806_), .ZN(G1340gat));
  OR3_X1    g606(.A1(new_n795_), .A2(KEYINPUT59), .A3(new_n737_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n804_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n808_), .B(new_n679_), .C1(new_n809_), .C2(new_n797_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(G120gat), .ZN(new_n811_));
  INV_X1    g610(.A(new_n788_), .ZN(new_n812_));
  INV_X1    g611(.A(G120gat), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n572_), .B2(KEYINPUT60), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n812_), .B(new_n814_), .C1(KEYINPUT60), .C2(new_n813_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n811_), .A2(new_n815_), .ZN(G1341gat));
  INV_X1    g615(.A(G127gat), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n788_), .B2(new_n319_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT122), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  OAI211_X1 g619(.A(KEYINPUT122), .B(new_n817_), .C1(new_n788_), .C2(new_n319_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n802_), .A2(new_n817_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n805_), .B2(new_n823_), .ZN(G1342gat));
  AOI21_X1  g623(.A(G134gat), .B1(new_n812_), .B2(new_n599_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n779_), .A2(G134gat), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n825_), .B1(new_n805_), .B2(new_n826_), .ZN(G1343gat));
  NOR3_X1   g626(.A1(new_n803_), .A2(new_n539_), .A3(new_n386_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n437_), .A2(new_n522_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(new_n449_), .A3(new_n589_), .ZN(new_n832_));
  OAI21_X1  g631(.A(G141gat), .B1(new_n830_), .B2(new_n682_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(G1344gat));
  NAND3_X1  g633(.A1(new_n831_), .A2(new_n450_), .A3(new_n679_), .ZN(new_n835_));
  OAI21_X1  g634(.A(G148gat), .B1(new_n830_), .B2(new_n572_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(G1345gat));
  XNOR2_X1  g636(.A(KEYINPUT61), .B(G155gat), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(KEYINPUT123), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n839_), .B1(new_n831_), .B2(new_n318_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n839_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n830_), .A2(new_n319_), .A3(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n840_), .A2(new_n842_), .ZN(G1346gat));
  NAND2_X1  g642(.A1(new_n831_), .A2(new_n599_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n634_), .A2(new_n272_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(KEYINPUT124), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n844_), .A2(new_n272_), .B1(new_n831_), .B2(new_n846_), .ZN(G1347gat));
  NOR4_X1   g646(.A1(new_n548_), .A2(new_n542_), .A3(new_n489_), .A4(new_n605_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n801_), .A2(new_n319_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(new_n786_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n589_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(G169gat), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(new_n404_), .B2(new_n852_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(KEYINPUT62), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT62), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n853_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(G1348gat));
  NOR2_X1   g657(.A1(new_n803_), .A2(new_n849_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n342_), .B1(new_n859_), .B2(new_n679_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n848_), .B1(new_n794_), .B2(new_n787_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n861_), .A2(G176gat), .A3(new_n572_), .ZN(new_n862_));
  OR3_X1    g661(.A1(new_n860_), .A2(new_n862_), .A3(KEYINPUT125), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT125), .B1(new_n860_), .B2(new_n862_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(G1349gat));
  AOI21_X1  g664(.A(G183gat), .B1(new_n859_), .B2(new_n318_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n861_), .A2(new_n407_), .A3(new_n802_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1350gat));
  NAND3_X1  g667(.A1(new_n851_), .A2(new_n599_), .A3(new_n335_), .ZN(new_n869_));
  OAI21_X1  g668(.A(G190gat), .B1(new_n861_), .B2(new_n626_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1351gat));
  INV_X1    g670(.A(new_n803_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n548_), .A2(new_n522_), .A3(new_n489_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT126), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n605_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n872_), .A2(new_n875_), .A3(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n584_), .B1(new_n877_), .B2(new_n682_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT127), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n877_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n881_), .A2(G197gat), .A3(new_n589_), .ZN(new_n882_));
  OAI211_X1 g681(.A(KEYINPUT127), .B(new_n584_), .C1(new_n877_), .C2(new_n682_), .ZN(new_n883_));
  AND3_X1   g682(.A1(new_n880_), .A2(new_n882_), .A3(new_n883_), .ZN(G1352gat));
  NOR2_X1   g683(.A1(new_n877_), .A2(new_n572_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(new_n563_), .ZN(G1353gat));
  AOI211_X1 g685(.A(KEYINPUT63), .B(G211gat), .C1(new_n881_), .C2(new_n317_), .ZN(new_n887_));
  XOR2_X1   g686(.A(KEYINPUT63), .B(G211gat), .Z(new_n888_));
  AND3_X1   g687(.A1(new_n881_), .A2(new_n317_), .A3(new_n888_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n887_), .A2(new_n889_), .ZN(G1354gat));
  AND3_X1   g689(.A1(new_n881_), .A2(G218gat), .A3(new_n779_), .ZN(new_n891_));
  AOI21_X1  g690(.A(G218gat), .B1(new_n881_), .B2(new_n599_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1355gat));
endmodule


