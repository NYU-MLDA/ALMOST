//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 1 0 0 1 1 1 0 0 0 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n774_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT23), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G183gat), .A3(G190gat), .ZN(new_n205_));
  AND2_X1   g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT82), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT82), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G190gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(new_n210_), .A3(KEYINPUT26), .ZN(new_n211_));
  OR2_X1    g010(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT25), .B(G183gat), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n206_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT24), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n216_), .B1(G169gat), .B2(G176gat), .ZN(new_n217_));
  INV_X1    g016(.A(G169gat), .ZN(new_n218_));
  INV_X1    g017(.A(G176gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n218_), .A2(new_n219_), .A3(KEYINPUT83), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT83), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n221_), .B1(G169gat), .B2(G176gat), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n220_), .A2(new_n222_), .A3(KEYINPUT84), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT84), .B1(new_n220_), .B2(new_n222_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n217_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT84), .ZN(new_n226_));
  NOR3_X1   g025(.A1(new_n221_), .A2(G169gat), .A3(G176gat), .ZN(new_n227_));
  AOI21_X1  g026(.A(KEYINPUT83), .B1(new_n218_), .B2(new_n219_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n226_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n220_), .A2(new_n222_), .A3(KEYINPUT84), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(new_n216_), .A3(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n215_), .A2(new_n225_), .A3(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(KEYINPUT85), .A2(G169gat), .ZN(new_n234_));
  AOI21_X1  g033(.A(G176gat), .B1(new_n234_), .B2(KEYINPUT22), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n235_), .B1(KEYINPUT22), .B2(new_n234_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n205_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT86), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n203_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n202_), .A2(KEYINPUT86), .A3(KEYINPUT23), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n237_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(G183gat), .B1(new_n208_), .B2(new_n210_), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n233_), .B(new_n236_), .C1(new_n241_), .C2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n232_), .A2(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n244_), .A2(KEYINPUT30), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT30), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n246_), .B1(new_n232_), .B2(new_n243_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT90), .B1(new_n248_), .B2(KEYINPUT87), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT87), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT90), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n250_), .B(new_n251_), .C1(new_n245_), .C2(new_n247_), .ZN(new_n252_));
  INV_X1    g051(.A(G127gat), .ZN(new_n253_));
  INV_X1    g052(.A(G134gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(G113gat), .ZN(new_n256_));
  INV_X1    g055(.A(G120gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G127gat), .A2(G134gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G113gat), .A2(G120gat), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n255_), .A2(new_n258_), .A3(new_n259_), .A4(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT89), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n255_), .A2(new_n259_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n258_), .A2(new_n260_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(new_n261_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n263_), .B1(KEYINPUT89), .B2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT31), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT88), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n249_), .A2(new_n252_), .A3(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n272_), .B1(new_n249_), .B2(new_n252_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G71gat), .B(G99gat), .ZN(new_n276_));
  INV_X1    g075(.A(G43gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G227gat), .A2(G233gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(G15gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n278_), .B(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n282_), .B1(new_n248_), .B2(KEYINPUT87), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NOR3_X1   g083(.A1(new_n274_), .A2(new_n275_), .A3(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n249_), .A2(new_n252_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(new_n271_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n283_), .B1(new_n287_), .B2(new_n273_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n285_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G226gat), .A2(G233gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT19), .ZN(new_n291_));
  INV_X1    g090(.A(G204gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(G197gat), .ZN(new_n293_));
  INV_X1    g092(.A(G197gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(G204gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(G211gat), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n297_), .A2(G218gat), .ZN(new_n298_));
  INV_X1    g097(.A(G218gat), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n299_), .A2(G211gat), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n296_), .B(KEYINPUT21), .C1(new_n298_), .C2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G211gat), .B(G218gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G197gat), .B(G204gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT21), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n302_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n296_), .A2(KEYINPUT21), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n301_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n232_), .A2(new_n308_), .A3(new_n243_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT20), .ZN(new_n310_));
  AOI21_X1  g109(.A(KEYINPUT24), .B1(new_n220_), .B2(new_n222_), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT97), .B1(new_n241_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n240_), .ZN(new_n313_));
  AOI21_X1  g112(.A(KEYINPUT86), .B1(new_n202_), .B2(KEYINPUT23), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n205_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT97), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n216_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT26), .B(G190gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n214_), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n312_), .A2(new_n318_), .A3(new_n320_), .A4(new_n225_), .ZN(new_n321_));
  XOR2_X1   g120(.A(KEYINPUT22), .B(G169gat), .Z(new_n322_));
  NOR2_X1   g121(.A1(G183gat), .A2(G190gat), .ZN(new_n323_));
  OAI221_X1 g122(.A(new_n233_), .B1(new_n322_), .B2(G176gat), .C1(new_n206_), .C2(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n308_), .B1(new_n321_), .B2(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n291_), .B1(new_n310_), .B2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G8gat), .B(G36gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G64gat), .B(G92gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n244_), .A2(new_n307_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n321_), .A2(new_n308_), .A3(new_n324_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n291_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n332_), .A2(new_n333_), .A3(KEYINPUT20), .A4(new_n334_), .ZN(new_n335_));
  AND3_X1   g134(.A1(new_n326_), .A2(new_n331_), .A3(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n331_), .B1(new_n326_), .B2(new_n335_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT27), .ZN(new_n340_));
  INV_X1    g139(.A(new_n331_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n332_), .A2(new_n333_), .A3(KEYINPUT20), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n291_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n309_), .A2(KEYINPUT20), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n321_), .A2(new_n324_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(new_n307_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT102), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n344_), .A2(new_n346_), .A3(new_n347_), .A4(new_n334_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n343_), .A2(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n310_), .A2(new_n325_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n347_), .B1(new_n350_), .B2(new_n334_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n341_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n336_), .A2(new_n340_), .ZN(new_n353_));
  AOI22_X1  g152(.A1(new_n339_), .A2(new_n340_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n289_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT96), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G78gat), .B(G106gat), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n357_), .B(KEYINPUT95), .Z(new_n358_));
  XOR2_X1   g157(.A(G155gat), .B(G162gat), .Z(new_n359_));
  INV_X1    g158(.A(KEYINPUT93), .ZN(new_n360_));
  INV_X1    g159(.A(G141gat), .ZN(new_n361_));
  INV_X1    g160(.A(G148gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT3), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT3), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n360_), .A2(new_n365_), .A3(new_n361_), .A4(new_n362_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n364_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G141gat), .A2(G148gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT92), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT92), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n371_), .A2(G141gat), .A3(G148gat), .ZN(new_n372_));
  AOI21_X1  g171(.A(KEYINPUT2), .B1(new_n370_), .B2(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n359_), .B1(new_n368_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(G155gat), .ZN(new_n375_));
  INV_X1    g174(.A(G162gat), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT1), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT1), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n378_), .A2(G155gat), .A3(G162gat), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n377_), .B(new_n379_), .C1(G155gat), .C2(G162gat), .ZN(new_n380_));
  AOI22_X1  g179(.A1(new_n370_), .A2(new_n372_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n374_), .A2(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n308_), .B1(new_n383_), .B2(KEYINPUT29), .ZN(new_n384_));
  INV_X1    g183(.A(G228gat), .ZN(new_n385_));
  INV_X1    g184(.A(G233gat), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n384_), .A2(new_n388_), .ZN(new_n389_));
  AOI211_X1 g188(.A(new_n387_), .B(new_n308_), .C1(KEYINPUT29), .C2(new_n383_), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n356_), .B(new_n358_), .C1(new_n389_), .C2(new_n390_), .ZN(new_n391_));
  OR2_X1    g190(.A1(new_n384_), .A2(new_n388_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n384_), .A2(new_n388_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n358_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n392_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n391_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n384_), .B(new_n388_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n356_), .B1(new_n397_), .B2(new_n358_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n370_), .A2(new_n372_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT2), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n401_), .A2(new_n366_), .A3(new_n364_), .A4(new_n367_), .ZN(new_n402_));
  AOI22_X1  g201(.A1(new_n402_), .A2(new_n359_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT28), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT29), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n403_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT28), .B1(new_n383_), .B2(KEYINPUT29), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G22gat), .B(G50gat), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n406_), .A2(new_n407_), .A3(new_n409_), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n411_), .A2(KEYINPUT94), .A3(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(KEYINPUT94), .B1(new_n411_), .B2(new_n412_), .ZN(new_n414_));
  OAI22_X1  g213(.A1(new_n396_), .A2(new_n398_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n397_), .A2(new_n357_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n416_), .A2(new_n412_), .A3(new_n411_), .A4(new_n395_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G1gat), .B(G29gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G57gat), .B(G85gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G225gat), .A2(G233gat), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n374_), .A2(new_n382_), .A3(new_n267_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n267_), .A2(KEYINPUT89), .ZN(new_n426_));
  INV_X1    g225(.A(new_n263_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n425_), .B1(new_n403_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT4), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT4), .B1(new_n383_), .B2(new_n268_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n424_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n425_), .B(new_n424_), .C1(new_n403_), .C2(new_n428_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT100), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n383_), .A2(new_n268_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n437_), .A2(KEYINPUT100), .A3(new_n424_), .A4(new_n425_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n423_), .B1(new_n433_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n424_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT4), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n442_), .B1(new_n437_), .B2(new_n425_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n441_), .B1(new_n443_), .B2(new_n431_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n423_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n444_), .A2(new_n445_), .A3(new_n438_), .A4(new_n436_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n440_), .A2(new_n446_), .A3(KEYINPUT103), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT103), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n448_), .B(new_n423_), .C1(new_n433_), .C2(new_n439_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NOR3_X1   g250(.A1(new_n355_), .A2(new_n418_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT105), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n331_), .A2(KEYINPUT32), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n455_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n331_), .A2(KEYINPUT32), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n326_), .A2(new_n457_), .A3(new_n335_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n447_), .A2(new_n456_), .A3(new_n449_), .A4(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n441_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n437_), .A2(new_n441_), .A3(new_n425_), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n461_), .A2(KEYINPUT101), .A3(new_n423_), .ZN(new_n462_));
  AOI21_X1  g261(.A(KEYINPUT101), .B1(new_n461_), .B2(new_n423_), .ZN(new_n463_));
  OR3_X1    g262(.A1(new_n460_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT33), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n446_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n439_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n467_), .A2(KEYINPUT33), .A3(new_n445_), .A4(new_n444_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n338_), .A2(new_n464_), .A3(new_n466_), .A4(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n418_), .B1(new_n459_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT104), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n415_), .A2(new_n417_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n470_), .A2(new_n471_), .B1(new_n472_), .B2(new_n354_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n459_), .A2(new_n469_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n418_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT104), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n473_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT91), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n479_), .B1(new_n285_), .B2(new_n288_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n284_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n287_), .A2(new_n283_), .A3(new_n273_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n481_), .A2(new_n482_), .A3(KEYINPUT91), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n480_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n454_), .B1(new_n478_), .B2(new_n485_), .ZN(new_n486_));
  AOI211_X1 g285(.A(KEYINPUT105), .B(new_n484_), .C1(new_n473_), .C2(new_n477_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n453_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G71gat), .B(G78gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G57gat), .B(G64gat), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n489_), .B1(KEYINPUT11), .B2(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n491_), .B1(KEYINPUT11), .B2(new_n490_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n489_), .A3(KEYINPUT11), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT78), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G231gat), .A2(G233gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT76), .B(G1gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(G8gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT14), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT77), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G15gat), .B(G22gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G1gat), .B(G8gat), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n504_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n497_), .B(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G127gat), .B(G155gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(new_n297_), .ZN(new_n512_));
  XOR2_X1   g311(.A(KEYINPUT16), .B(G183gat), .Z(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n514_), .A2(KEYINPUT17), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n514_), .A2(KEYINPUT17), .ZN(new_n516_));
  OR3_X1    g315(.A1(new_n510_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  OR2_X1    g316(.A1(new_n517_), .A2(KEYINPUT79), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n510_), .A2(new_n515_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n517_), .A2(KEYINPUT79), .A3(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT66), .B(KEYINPUT6), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G99gat), .A2(G106gat), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n523_), .B(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(G106gat), .ZN(new_n527_));
  XOR2_X1   g326(.A(KEYINPUT10), .B(G99gat), .Z(new_n528_));
  AOI21_X1  g327(.A(new_n526_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT64), .B(G92gat), .ZN(new_n530_));
  AOI21_X1  g329(.A(KEYINPUT9), .B1(new_n530_), .B2(G85gat), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n531_), .A2(KEYINPUT65), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(KEYINPUT65), .ZN(new_n533_));
  NOR2_X1   g332(.A1(G85gat), .A2(G92gat), .ZN(new_n534_));
  AND2_X1   g333(.A1(G85gat), .A2(G92gat), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n534_), .B1(new_n535_), .B2(KEYINPUT9), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n533_), .A2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n529_), .B1(new_n532_), .B2(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(G99gat), .A2(G106gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT7), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n526_), .A2(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n535_), .A2(new_n534_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n542_), .A2(KEYINPUT8), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT8), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n523_), .B(new_n524_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n540_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n546_), .B1(new_n548_), .B2(new_n543_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n538_), .B1(new_n545_), .B2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G29gat), .B(G36gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G43gat), .B(G50gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT15), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT35), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G232gat), .A2(G233gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT34), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  AOI22_X1  g357(.A1(new_n550_), .A2(new_n554_), .B1(new_n555_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n553_), .ZN(new_n560_));
  OAI21_X1  g359(.A(KEYINPUT71), .B1(new_n550_), .B2(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT8), .B1(new_n542_), .B2(new_n544_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n548_), .A2(new_n546_), .A3(new_n543_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT71), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n564_), .A2(new_n565_), .A3(new_n538_), .A4(new_n553_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n559_), .A2(new_n561_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT70), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n558_), .A2(new_n555_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT70), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n559_), .A2(new_n561_), .A3(new_n566_), .A4(new_n570_), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n568_), .A2(new_n569_), .A3(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n569_), .B1(new_n568_), .B2(new_n571_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  XOR2_X1   g373(.A(G190gat), .B(G218gat), .Z(new_n575_));
  XNOR2_X1  g374(.A(G134gat), .B(G162gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT36), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n578_), .B(KEYINPUT73), .Z(new_n579_));
  NAND2_X1  g378(.A1(new_n574_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT74), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n574_), .A2(KEYINPUT74), .A3(new_n579_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT36), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n577_), .A2(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n585_), .B(KEYINPUT72), .Z(new_n586_));
  OAI21_X1  g385(.A(new_n586_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n582_), .A2(new_n583_), .A3(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(KEYINPUT37), .ZN(new_n589_));
  INV_X1    g388(.A(new_n573_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n568_), .A2(new_n569_), .A3(new_n571_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n590_), .A2(new_n591_), .A3(new_n578_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(new_n587_), .ZN(new_n593_));
  OAI21_X1  g392(.A(KEYINPUT75), .B1(new_n593_), .B2(KEYINPUT37), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT75), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT37), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n592_), .A2(new_n587_), .A3(new_n595_), .A4(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n594_), .A2(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n522_), .B1(new_n589_), .B2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G230gat), .A2(G233gat), .ZN(new_n600_));
  INV_X1    g399(.A(new_n494_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n550_), .A2(new_n601_), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n538_), .B(new_n494_), .C1(new_n545_), .C2(new_n549_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n600_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n600_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT67), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n603_), .A2(KEYINPUT67), .A3(new_n600_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n550_), .A2(KEYINPUT12), .A3(new_n601_), .ZN(new_n610_));
  AOI21_X1  g409(.A(KEYINPUT12), .B1(new_n550_), .B2(new_n601_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n604_), .B1(new_n609_), .B2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT69), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(G176gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G120gat), .B(G148gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(new_n292_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n616_), .B(new_n618_), .Z(new_n619_));
  XNOR2_X1  g418(.A(new_n613_), .B(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT13), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n621_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT81), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n553_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n502_), .A2(new_n503_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n504_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n629_), .A2(new_n560_), .A3(new_n505_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n626_), .A2(KEYINPUT80), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(G229gat), .A2(G233gat), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT80), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n508_), .A2(new_n634_), .A3(new_n560_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n631_), .A2(new_n633_), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n508_), .A2(new_n554_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n637_), .A2(new_n632_), .A3(new_n626_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(G113gat), .B(G141gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(G169gat), .B(G197gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n625_), .B1(new_n639_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n642_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n636_), .A2(KEYINPUT81), .A3(new_n638_), .A4(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n639_), .A2(new_n642_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n624_), .A2(new_n649_), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n488_), .A2(new_n599_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n498_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n651_), .A2(new_n652_), .A3(new_n451_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT106), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n488_), .A2(new_n650_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT107), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n593_), .B(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n657_), .A2(new_n522_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n655_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(new_n451_), .ZN(new_n660_));
  AOI22_X1  g459(.A1(new_n654_), .A2(KEYINPUT38), .B1(G1gat), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT106), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n653_), .B(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT38), .ZN(new_n664_));
  AND3_X1   g463(.A1(new_n663_), .A2(KEYINPUT108), .A3(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT108), .B1(new_n663_), .B2(new_n664_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n661_), .B1(new_n665_), .B2(new_n666_), .ZN(G1324gat));
  INV_X1    g466(.A(G8gat), .ZN(new_n668_));
  INV_X1    g467(.A(new_n354_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n651_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n488_), .A2(new_n650_), .A3(new_n669_), .A4(new_n658_), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n671_), .A2(KEYINPUT109), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n668_), .B1(new_n671_), .B2(KEYINPUT109), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT39), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n672_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n670_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT40), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n677_), .B(new_n678_), .ZN(G1325gat));
  NAND2_X1  g478(.A1(new_n659_), .A2(new_n484_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(G15gat), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n681_), .A2(KEYINPUT41), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(KEYINPUT41), .ZN(new_n683_));
  INV_X1    g482(.A(G15gat), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n651_), .A2(new_n684_), .A3(new_n484_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n682_), .A2(new_n683_), .A3(new_n685_), .ZN(G1326gat));
  XNOR2_X1  g485(.A(new_n418_), .B(KEYINPUT110), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n659_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(G22gat), .ZN(new_n689_));
  XOR2_X1   g488(.A(KEYINPUT111), .B(KEYINPUT42), .Z(new_n690_));
  OR2_X1    g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n690_), .ZN(new_n692_));
  INV_X1    g491(.A(G22gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n651_), .A2(new_n693_), .A3(new_n687_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n691_), .A2(new_n692_), .A3(new_n694_), .ZN(G1327gat));
  INV_X1    g494(.A(KEYINPUT112), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n696_), .A2(KEYINPUT43), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(KEYINPUT43), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n474_), .A2(new_n471_), .A3(new_n475_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n354_), .A2(new_n472_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n470_), .A2(new_n471_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n485_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT105), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n478_), .A2(new_n454_), .A3(new_n485_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n452_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n589_), .A2(new_n598_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n697_), .B(new_n698_), .C1(new_n706_), .C2(new_n707_), .ZN(new_n708_));
  AOI22_X1  g507(.A1(new_n588_), .A2(KEYINPUT37), .B1(new_n594_), .B2(new_n597_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n488_), .A2(new_n696_), .A3(KEYINPUT43), .A4(new_n709_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n624_), .A2(new_n521_), .A3(new_n649_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n708_), .A2(new_n710_), .A3(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n708_), .A2(new_n710_), .A3(KEYINPUT44), .A4(new_n711_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n714_), .A2(new_n451_), .A3(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(G29gat), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n593_), .B(KEYINPUT107), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n718_), .A2(new_n521_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n655_), .A2(new_n719_), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n450_), .A2(G29gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(G1328gat));
  NAND3_X1  g521(.A1(new_n714_), .A2(new_n669_), .A3(new_n715_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G36gat), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n354_), .A2(G36gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n655_), .A2(new_n719_), .A3(new_n725_), .ZN(new_n726_));
  XOR2_X1   g525(.A(KEYINPUT113), .B(KEYINPUT45), .Z(new_n727_));
  XNOR2_X1  g526(.A(new_n726_), .B(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n724_), .A2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(KEYINPUT114), .B(KEYINPUT46), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n724_), .A2(new_n728_), .A3(new_n730_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1329gat));
  NAND4_X1  g533(.A1(new_n714_), .A2(G43gat), .A3(new_n289_), .A4(new_n715_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n277_), .B1(new_n720_), .B2(new_n485_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g537(.A(G50gat), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n714_), .A2(new_n418_), .A3(new_n715_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT115), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n739_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n742_), .B1(new_n741_), .B2(new_n740_), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n655_), .A2(new_n739_), .A3(new_n687_), .A4(new_n719_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1331gat));
  INV_X1    g544(.A(new_n624_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n706_), .A2(new_n648_), .A3(new_n746_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n747_), .A2(new_n599_), .ZN(new_n748_));
  AOI21_X1  g547(.A(G57gat), .B1(new_n748_), .B2(new_n451_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n747_), .A2(new_n658_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n451_), .A2(G57gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n749_), .B1(new_n750_), .B2(new_n751_), .ZN(G1332gat));
  INV_X1    g551(.A(G64gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n750_), .B2(new_n669_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT48), .Z(new_n755_));
  NAND3_X1  g554(.A1(new_n748_), .A2(new_n753_), .A3(new_n669_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1333gat));
  INV_X1    g556(.A(G71gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n750_), .B2(new_n484_), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT49), .Z(new_n760_));
  NAND3_X1  g559(.A1(new_n748_), .A2(new_n758_), .A3(new_n484_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(G1334gat));
  INV_X1    g561(.A(G78gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n763_), .B1(new_n750_), .B2(new_n687_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT50), .Z(new_n765_));
  NAND3_X1  g564(.A1(new_n748_), .A2(new_n763_), .A3(new_n687_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(G1335gat));
  AND2_X1   g566(.A1(new_n747_), .A2(new_n719_), .ZN(new_n768_));
  AOI21_X1  g567(.A(G85gat), .B1(new_n768_), .B2(new_n451_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n746_), .A2(new_n521_), .A3(new_n648_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n708_), .A2(new_n710_), .A3(new_n770_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n451_), .A2(G85gat), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n769_), .B1(new_n771_), .B2(new_n772_), .ZN(G1336gat));
  AOI21_X1  g572(.A(G92gat), .B1(new_n768_), .B2(new_n669_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n669_), .A2(new_n530_), .ZN(new_n775_));
  XOR2_X1   g574(.A(new_n775_), .B(KEYINPUT116), .Z(new_n776_));
  AOI21_X1  g575(.A(new_n774_), .B1(new_n771_), .B2(new_n776_), .ZN(G1337gat));
  NAND3_X1  g576(.A1(new_n768_), .A2(new_n528_), .A3(new_n289_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n771_), .A2(new_n484_), .ZN(new_n779_));
  INV_X1    g578(.A(G99gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n778_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g581(.A1(new_n768_), .A2(new_n527_), .A3(new_n418_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n708_), .A2(new_n710_), .A3(new_n418_), .A4(new_n770_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n784_), .A2(new_n785_), .A3(G106gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n784_), .B2(G106gat), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n783_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  XOR2_X1   g587(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n789_));
  XNOR2_X1  g588(.A(new_n788_), .B(new_n789_), .ZN(G1339gat));
  INV_X1    g589(.A(KEYINPUT58), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT56), .ZN(new_n792_));
  INV_X1    g591(.A(new_n611_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n550_), .A2(KEYINPUT12), .A3(new_n601_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n603_), .A2(KEYINPUT67), .A3(new_n600_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT67), .B1(new_n603_), .B2(new_n600_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n793_), .B(new_n794_), .C1(new_n795_), .C2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT118), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n609_), .A2(KEYINPUT55), .A3(new_n612_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n793_), .A2(new_n603_), .A3(new_n794_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n600_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n799_), .A2(new_n800_), .A3(new_n801_), .A4(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n619_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  AOI22_X1  g606(.A1(new_n797_), .A2(new_n798_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n800_), .B1(new_n808_), .B2(new_n801_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n792_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT119), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n799_), .A2(new_n801_), .A3(new_n804_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT118), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n813_), .A2(KEYINPUT56), .A3(new_n806_), .A4(new_n805_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n810_), .A2(new_n811_), .A3(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n631_), .A2(new_n632_), .A3(new_n635_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n637_), .A2(new_n633_), .A3(new_n626_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(new_n642_), .A3(new_n817_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n646_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n613_), .A2(new_n619_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n819_), .B(new_n820_), .C1(new_n814_), .C2(new_n811_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n791_), .B1(new_n815_), .B2(new_n821_), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n814_), .A2(new_n811_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n819_), .A2(new_n820_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n810_), .A2(new_n811_), .A3(new_n814_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n823_), .A2(new_n824_), .A3(new_n825_), .A4(KEYINPUT58), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n822_), .A2(new_n709_), .A3(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT57), .ZN(new_n828_));
  AND3_X1   g627(.A1(new_n620_), .A2(new_n646_), .A3(new_n818_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n810_), .A2(new_n814_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n648_), .A2(new_n820_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n829_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n828_), .B1(new_n832_), .B2(new_n657_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n648_), .A2(new_n820_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n834_), .B1(new_n810_), .B2(new_n814_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n718_), .B(KEYINPUT57), .C1(new_n835_), .C2(new_n829_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n833_), .A2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n522_), .B1(new_n827_), .B2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n624_), .A2(new_n648_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n707_), .A2(new_n521_), .A3(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT54), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n599_), .A2(new_n842_), .A3(new_n839_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n838_), .A2(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n355_), .A2(new_n450_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n845_), .A2(new_n475_), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n648_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n256_), .ZN(new_n849_));
  XOR2_X1   g648(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n850_));
  NAND4_X1  g649(.A1(new_n845_), .A2(new_n475_), .A3(new_n846_), .A4(new_n850_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n649_), .A2(new_n256_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(KEYINPUT59), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n851_), .B(new_n852_), .C1(new_n847_), .C2(new_n854_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n849_), .A2(new_n855_), .ZN(G1340gat));
  OAI211_X1 g655(.A(new_n624_), .B(new_n851_), .C1(new_n847_), .C2(new_n854_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(G120gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n257_), .B1(new_n746_), .B2(KEYINPUT60), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n847_), .B(new_n859_), .C1(KEYINPUT60), .C2(new_n257_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(G1341gat));
  NAND2_X1  g660(.A1(new_n847_), .A2(new_n521_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n253_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n522_), .A2(new_n253_), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n851_), .B(new_n864_), .C1(new_n847_), .C2(new_n854_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n863_), .A2(new_n865_), .ZN(G1342gat));
  NAND2_X1  g665(.A1(new_n847_), .A2(new_n657_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n254_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n707_), .A2(new_n254_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n851_), .B(new_n869_), .C1(new_n847_), .C2(new_n854_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n868_), .A2(new_n870_), .ZN(G1343gat));
  NOR4_X1   g670(.A1(new_n484_), .A2(new_n475_), .A3(new_n450_), .A4(new_n669_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n845_), .A2(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n649_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(new_n361_), .ZN(G1344gat));
  NOR2_X1   g674(.A1(new_n873_), .A2(new_n746_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(new_n362_), .ZN(G1345gat));
  OAI21_X1  g676(.A(KEYINPUT121), .B1(new_n873_), .B2(new_n522_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT121), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n845_), .A2(new_n879_), .A3(new_n521_), .A4(new_n872_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(KEYINPUT61), .B(G155gat), .ZN(new_n881_));
  AND3_X1   g680(.A1(new_n878_), .A2(new_n880_), .A3(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n881_), .B1(new_n878_), .B2(new_n880_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1346gat));
  NOR3_X1   g683(.A1(new_n873_), .A2(new_n376_), .A3(new_n707_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n873_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n657_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n885_), .B1(new_n376_), .B2(new_n887_), .ZN(G1347gat));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n484_), .A2(new_n450_), .A3(new_n669_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n687_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n892_), .B1(new_n838_), .B2(new_n844_), .ZN(new_n893_));
  AOI211_X1 g692(.A(KEYINPUT122), .B(new_n218_), .C1(new_n893_), .C2(new_n648_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n895_));
  AND2_X1   g694(.A1(new_n833_), .A2(new_n836_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n822_), .A2(new_n826_), .A3(new_n709_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n521_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n599_), .A2(new_n842_), .A3(new_n839_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n842_), .B1(new_n599_), .B2(new_n839_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n648_), .B(new_n891_), .C1(new_n898_), .C2(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n895_), .B1(new_n902_), .B2(G169gat), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n889_), .B1(new_n894_), .B2(new_n903_), .ZN(new_n904_));
  AOI211_X1 g703(.A(new_n649_), .B(new_n892_), .C1(new_n838_), .C2(new_n844_), .ZN(new_n905_));
  OAI21_X1  g704(.A(KEYINPUT122), .B1(new_n905_), .B2(new_n218_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n902_), .A2(new_n895_), .A3(G169gat), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n906_), .A2(KEYINPUT62), .A3(new_n907_), .ZN(new_n908_));
  OR2_X1    g707(.A1(new_n902_), .A2(new_n322_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n904_), .A2(new_n908_), .A3(new_n909_), .ZN(G1348gat));
  AOI21_X1  g709(.A(G176gat), .B1(new_n893_), .B2(new_n624_), .ZN(new_n911_));
  AOI211_X1 g710(.A(new_n418_), .B(new_n890_), .C1(new_n838_), .C2(new_n844_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n746_), .A2(new_n219_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n911_), .B1(new_n912_), .B2(new_n913_), .ZN(G1349gat));
  AOI21_X1  g713(.A(G183gat), .B1(new_n912_), .B2(new_n521_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n522_), .A2(new_n214_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n915_), .B1(new_n893_), .B2(new_n916_), .ZN(G1350gat));
  NAND3_X1  g716(.A1(new_n893_), .A2(new_n319_), .A3(new_n657_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n893_), .A2(new_n709_), .ZN(new_n919_));
  AND3_X1   g718(.A1(new_n919_), .A2(KEYINPUT123), .A3(G190gat), .ZN(new_n920_));
  AOI21_X1  g719(.A(KEYINPUT123), .B1(new_n919_), .B2(G190gat), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n918_), .B1(new_n920_), .B2(new_n921_), .ZN(G1351gat));
  NOR4_X1   g721(.A1(new_n484_), .A2(new_n475_), .A3(new_n451_), .A4(new_n354_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n845_), .A2(new_n923_), .ZN(new_n924_));
  OAI22_X1  g723(.A1(new_n924_), .A2(new_n649_), .B1(KEYINPUT124), .B2(new_n294_), .ZN(new_n925_));
  AND2_X1   g724(.A1(new_n294_), .A2(KEYINPUT124), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n925_), .B(new_n926_), .ZN(G1352gat));
  NAND3_X1  g726(.A1(new_n845_), .A2(new_n624_), .A3(new_n923_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(KEYINPUT125), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT125), .ZN(new_n930_));
  NAND4_X1  g729(.A1(new_n845_), .A2(new_n930_), .A3(new_n624_), .A4(new_n923_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n929_), .A2(G204gat), .A3(new_n931_), .ZN(new_n932_));
  OAI21_X1  g731(.A(KEYINPUT126), .B1(new_n928_), .B2(G204gat), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  NAND4_X1  g733(.A1(new_n929_), .A2(KEYINPUT126), .A3(G204gat), .A4(new_n931_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(G1353gat));
  NOR2_X1   g735(.A1(new_n924_), .A2(new_n522_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n938_));
  INV_X1    g737(.A(new_n938_), .ZN(new_n939_));
  OAI21_X1  g738(.A(KEYINPUT127), .B1(new_n937_), .B2(new_n939_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT127), .ZN(new_n941_));
  OAI211_X1 g740(.A(new_n941_), .B(new_n938_), .C1(new_n924_), .C2(new_n522_), .ZN(new_n942_));
  XOR2_X1   g741(.A(KEYINPUT63), .B(G211gat), .Z(new_n943_));
  AOI22_X1  g742(.A1(new_n940_), .A2(new_n942_), .B1(new_n937_), .B2(new_n943_), .ZN(G1354gat));
  AND2_X1   g743(.A1(new_n845_), .A2(new_n923_), .ZN(new_n945_));
  AOI21_X1  g744(.A(G218gat), .B1(new_n945_), .B2(new_n657_), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n924_), .A2(new_n299_), .A3(new_n707_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n946_), .A2(new_n947_), .ZN(G1355gat));
endmodule


