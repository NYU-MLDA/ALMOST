//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 1 1 0 1 1 0 0 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n869_, new_n870_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n916_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_, new_n934_;
  INV_X1    g000(.A(KEYINPUT65), .ZN(new_n202_));
  INV_X1    g001(.A(G85gat), .ZN(new_n203_));
  INV_X1    g002(.A(G92gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT64), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G92gat), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n203_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n202_), .B1(new_n208_), .B2(KEYINPUT9), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT9), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G92gat), .ZN(new_n211_));
  OAI211_X1 g010(.A(KEYINPUT65), .B(new_n210_), .C1(new_n211_), .C2(new_n203_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G85gat), .A2(G92gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n203_), .A2(new_n204_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n213_), .B1(new_n214_), .B2(KEYINPUT9), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n209_), .A2(KEYINPUT66), .A3(new_n212_), .A4(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(KEYINPUT10), .B(G99gat), .Z(new_n217_));
  INV_X1    g016(.A(G106gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT6), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT6), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G99gat), .A3(G106gat), .ZN(new_n222_));
  AOI22_X1  g021(.A1(new_n217_), .A2(new_n218_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n216_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT66), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n212_), .A2(new_n215_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n206_), .A2(G92gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n204_), .A2(KEYINPUT64), .ZN(new_n228_));
  OAI21_X1  g027(.A(G85gat), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(KEYINPUT65), .B1(new_n229_), .B2(new_n210_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n225_), .B1(new_n226_), .B2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n220_), .A2(new_n222_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT68), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n235_));
  INV_X1    g034(.A(G99gat), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n235_), .A2(new_n236_), .A3(new_n218_), .A4(KEYINPUT7), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT7), .ZN(new_n238_));
  OAI22_X1  g037(.A1(new_n238_), .A2(KEYINPUT67), .B1(G99gat), .B2(G106gat), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n235_), .A2(KEYINPUT7), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n237_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n220_), .A2(new_n222_), .A3(KEYINPUT68), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n234_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n214_), .A2(new_n213_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT8), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n241_), .A2(new_n232_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT8), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n247_), .A2(new_n248_), .A3(new_n244_), .ZN(new_n249_));
  AOI22_X1  g048(.A1(new_n224_), .A2(new_n231_), .B1(new_n246_), .B2(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(G43gat), .B(G50gat), .Z(new_n251_));
  XNOR2_X1  g050(.A(G29gat), .B(G36gat), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n252_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n250_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n231_), .A2(new_n216_), .A3(new_n223_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n244_), .ZN(new_n257_));
  AND3_X1   g056(.A1(new_n220_), .A2(new_n222_), .A3(KEYINPUT68), .ZN(new_n258_));
  AOI21_X1  g057(.A(KEYINPUT68), .B1(new_n220_), .B2(new_n222_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n257_), .B1(new_n260_), .B2(new_n241_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n249_), .B1(new_n261_), .B2(new_n248_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n256_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n253_), .A2(new_n254_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT15), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n263_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G232gat), .A2(G233gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT34), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT35), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT75), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n255_), .A2(new_n267_), .A3(new_n272_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n270_), .A2(new_n271_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n274_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n255_), .A2(new_n276_), .A3(new_n267_), .A4(new_n272_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(KEYINPUT74), .A3(new_n277_), .ZN(new_n278_));
  XOR2_X1   g077(.A(G190gat), .B(G218gat), .Z(new_n279_));
  XNOR2_X1  g078(.A(G134gat), .B(G162gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT36), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n275_), .A2(new_n277_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n281_), .A2(new_n282_), .ZN(new_n286_));
  AOI22_X1  g085(.A1(new_n278_), .A2(new_n284_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n278_), .A2(new_n284_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT101), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G78gat), .B(G106gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(G197gat), .B(G204gat), .Z(new_n293_));
  XNOR2_X1  g092(.A(G211gat), .B(G218gat), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n293_), .B1(KEYINPUT21), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(KEYINPUT21), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT85), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n299_), .A2(KEYINPUT2), .ZN(new_n300_));
  NOR2_X1   g099(.A1(G141gat), .A2(G148gat), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT3), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT2), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n303_), .B(new_n304_), .C1(new_n305_), .C2(new_n298_), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT86), .B1(new_n300_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT85), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n298_), .B(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(new_n305_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT86), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n298_), .A2(new_n305_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n312_), .B1(new_n302_), .B2(new_n301_), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n310_), .A2(new_n311_), .A3(new_n304_), .A4(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n307_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n315_), .A2(new_n319_), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n316_), .A2(KEYINPUT1), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n316_), .B1(new_n318_), .B2(KEYINPUT1), .ZN(new_n322_));
  AOI211_X1 g121(.A(new_n301_), .B(new_n299_), .C1(new_n321_), .C2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n320_), .A2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n297_), .B1(new_n325_), .B2(KEYINPUT29), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G228gat), .A2(G233gat), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n327_), .B(KEYINPUT88), .Z(new_n328_));
  AND2_X1   g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(KEYINPUT88), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n326_), .A2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n292_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n326_), .A2(new_n328_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n333_), .B(new_n291_), .C1(new_n326_), .C2(new_n330_), .ZN(new_n334_));
  AOI21_X1  g133(.A(KEYINPUT87), .B1(new_n332_), .B2(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(G22gat), .B(G50gat), .Z(new_n336_));
  INV_X1    g135(.A(new_n319_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n337_), .B1(new_n307_), .B2(new_n314_), .ZN(new_n338_));
  OR3_X1    g137(.A1(new_n338_), .A2(KEYINPUT29), .A3(new_n323_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT28), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n339_), .A2(KEYINPUT28), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n336_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n342_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n336_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n344_), .A2(new_n340_), .A3(new_n345_), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n343_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n335_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G1gat), .B(G29gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT0), .ZN(new_n350_));
  INV_X1    g149(.A(G57gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(new_n203_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G127gat), .B(G134gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G113gat), .B(G120gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n320_), .A2(new_n356_), .A3(new_n324_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G225gat), .A2(G233gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n356_), .B(KEYINPUT84), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n359_), .B1(new_n338_), .B2(new_n323_), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n357_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT94), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n338_), .A2(new_n323_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G127gat), .B(G134gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(new_n355_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT84), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT4), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT84), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n356_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n366_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n362_), .B1(new_n363_), .B2(new_n370_), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n366_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n372_), .B(KEYINPUT94), .C1(new_n323_), .C2(new_n338_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n358_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n357_), .A2(new_n360_), .A3(KEYINPUT4), .ZN(new_n375_));
  AOI211_X1 g174(.A(new_n353_), .B(new_n361_), .C1(new_n374_), .C2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT95), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT33), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(KEYINPUT94), .B1(new_n325_), .B2(new_n372_), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n363_), .A2(new_n362_), .A3(new_n370_), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n375_), .B(new_n358_), .C1(new_n379_), .C2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n358_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n357_), .A2(new_n360_), .A3(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n381_), .A2(new_n353_), .A3(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(G64gat), .B(G92gat), .Z(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT93), .ZN(new_n386_));
  XOR2_X1   g185(.A(G8gat), .B(G36gat), .Z(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G183gat), .A2(G190gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT23), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT23), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n393_), .A2(G183gat), .A3(G190gat), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT24), .ZN(new_n395_));
  NOR2_X1   g194(.A1(G169gat), .A2(G176gat), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n392_), .A2(new_n394_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT80), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n398_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n396_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G169gat), .A2(G176gat), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(KEYINPUT24), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT79), .ZN(new_n404_));
  INV_X1    g203(.A(G183gat), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n404_), .B1(new_n405_), .B2(KEYINPUT25), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT26), .B(G190gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT25), .B(G183gat), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n406_), .B(new_n407_), .C1(new_n408_), .C2(new_n404_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n399_), .A2(new_n400_), .A3(new_n403_), .A4(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n392_), .A2(new_n394_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n411_), .B1(G183gat), .B2(G190gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT22), .B(G169gat), .ZN(new_n413_));
  INV_X1    g212(.A(G176gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n412_), .A2(new_n415_), .A3(new_n402_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n410_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT81), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n410_), .A2(KEYINPUT81), .A3(new_n416_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n297_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n408_), .A2(new_n407_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n422_), .A2(new_n397_), .A3(new_n403_), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n423_), .A2(KEYINPUT89), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(KEYINPUT89), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT91), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT90), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n413_), .B(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n414_), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n412_), .A2(new_n402_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n426_), .A2(new_n427_), .A3(new_n432_), .A4(new_n297_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G226gat), .A2(G233gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT19), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT20), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n433_), .A2(new_n437_), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n424_), .A2(new_n425_), .B1(new_n431_), .B2(new_n430_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n427_), .B1(new_n439_), .B2(new_n297_), .ZN(new_n440_));
  NOR3_X1   g239(.A1(new_n421_), .A2(new_n438_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n435_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n426_), .A2(new_n432_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n297_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n436_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n419_), .A2(new_n420_), .A3(new_n297_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n442_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n390_), .B1(new_n441_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n447_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n419_), .A2(new_n420_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n444_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n440_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n451_), .A2(new_n452_), .A3(new_n433_), .A4(new_n437_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n390_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n449_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n384_), .A2(new_n448_), .A3(new_n455_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n375_), .B(new_n382_), .C1(new_n379_), .C2(new_n380_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n353_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n361_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n457_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT33), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n460_), .A2(KEYINPUT95), .A3(new_n461_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n378_), .A2(new_n456_), .A3(KEYINPUT96), .A4(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT32), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n390_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT97), .B(KEYINPUT20), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n297_), .A2(new_n423_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n466_), .B1(new_n467_), .B2(new_n432_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n442_), .B1(new_n451_), .B2(new_n468_), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n445_), .A2(new_n442_), .A3(new_n446_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n465_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n449_), .A2(new_n453_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n458_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n473_));
  OAI221_X1 g272(.A(new_n471_), .B1(new_n472_), .B2(new_n465_), .C1(new_n376_), .C2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n463_), .A2(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n461_), .B1(new_n460_), .B2(KEYINPUT95), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n384_), .A2(new_n448_), .A3(new_n455_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT96), .B1(new_n478_), .B2(new_n462_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n348_), .B1(new_n475_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n343_), .A2(new_n346_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n335_), .B(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n376_), .A2(new_n473_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT27), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n469_), .A2(new_n470_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT98), .ZN(new_n486_));
  AOI22_X1  g285(.A1(new_n485_), .A2(new_n390_), .B1(new_n455_), .B2(new_n486_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n455_), .A2(new_n486_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n484_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n448_), .A2(new_n455_), .A3(new_n484_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n482_), .B(new_n483_), .C1(new_n489_), .C2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n480_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT30), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n450_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n419_), .A2(KEYINPUT30), .A3(new_n420_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G227gat), .A2(G233gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(G15gat), .ZN(new_n498_));
  XOR2_X1   g297(.A(G71gat), .B(G99gat), .Z(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT82), .B(G43gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n496_), .A2(new_n502_), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n496_), .A2(KEYINPUT83), .A3(new_n502_), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT83), .B1(new_n496_), .B2(new_n502_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n503_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT31), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT31), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n508_), .B(new_n503_), .C1(new_n504_), .C2(new_n505_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(new_n359_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n359_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n507_), .A2(new_n509_), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n492_), .A2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n511_), .A2(new_n513_), .A3(new_n483_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n348_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n290_), .B1(new_n515_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n264_), .B(KEYINPUT78), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G15gat), .B(G22gat), .ZN(new_n523_));
  INV_X1    g322(.A(G1gat), .ZN(new_n524_));
  INV_X1    g323(.A(G8gat), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT14), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G1gat), .B(G8gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n527_), .B(new_n528_), .Z(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n522_), .B(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G229gat), .A2(G233gat), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n522_), .A2(new_n529_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n266_), .A2(new_n530_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(new_n532_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n534_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G113gat), .B(G141gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G169gat), .B(G197gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n539_), .A2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n534_), .A2(new_n538_), .A3(new_n542_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G57gat), .B(G64gat), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n548_), .A2(KEYINPUT11), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(KEYINPUT11), .ZN(new_n550_));
  XOR2_X1   g349(.A(G71gat), .B(G78gat), .Z(new_n551_));
  NAND3_X1  g350(.A1(new_n549_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n550_), .A2(new_n551_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n263_), .A2(KEYINPUT12), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT71), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n554_), .B1(new_n256_), .B2(new_n262_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n559_), .A2(KEYINPUT71), .A3(KEYINPUT12), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT12), .ZN(new_n562_));
  OAI211_X1 g361(.A(KEYINPUT72), .B(new_n562_), .C1(new_n250_), .C2(new_n554_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT72), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n564_), .B1(new_n559_), .B2(KEYINPUT12), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G230gat), .A2(G233gat), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n250_), .A2(new_n554_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n561_), .A2(new_n566_), .A3(new_n567_), .A4(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n263_), .A2(new_n555_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT70), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n559_), .A2(KEYINPUT70), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT69), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n574_), .B1(new_n263_), .B2(new_n555_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n250_), .A2(KEYINPUT69), .A3(new_n554_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n572_), .A2(new_n573_), .A3(new_n575_), .A4(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n567_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G120gat), .B(G148gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT5), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G176gat), .B(G204gat), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n581_), .B(new_n582_), .Z(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n569_), .A2(new_n579_), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n584_), .B1(new_n569_), .B2(new_n579_), .ZN(new_n587_));
  OAI21_X1  g386(.A(KEYINPUT13), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n587_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT13), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n589_), .A2(new_n590_), .A3(new_n585_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n588_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT73), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n588_), .A2(new_n591_), .A3(KEYINPUT73), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n547_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G127gat), .B(G155gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT16), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G183gat), .B(G211gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n600_), .A2(KEYINPUT17), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n529_), .B(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(new_n555_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n600_), .A2(KEYINPUT17), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n601_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(KEYINPUT77), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n607_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n596_), .A2(KEYINPUT100), .A3(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(KEYINPUT100), .B1(new_n596_), .B2(new_n610_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n521_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n483_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(G1gat), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT38), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n594_), .A2(new_n595_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n546_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n620_), .B1(new_n515_), .B2(new_n519_), .ZN(new_n621_));
  OR2_X1    g420(.A1(KEYINPUT76), .A2(KEYINPUT37), .ZN(new_n622_));
  NAND2_X1  g421(.A1(KEYINPUT76), .A2(KEYINPUT37), .ZN(new_n623_));
  AND4_X1   g422(.A1(new_n288_), .A2(new_n287_), .A3(new_n622_), .A4(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n623_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n610_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n621_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n629_), .A2(new_n524_), .A3(new_n615_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT99), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n632_), .A2(KEYINPUT102), .A3(new_n618_), .ZN(new_n633_));
  AOI21_X1  g432(.A(KEYINPUT102), .B1(new_n632_), .B2(new_n618_), .ZN(new_n634_));
  OAI221_X1 g433(.A(new_n617_), .B1(new_n618_), .B2(new_n632_), .C1(new_n633_), .C2(new_n634_), .ZN(G1324gat));
  INV_X1    g434(.A(KEYINPUT40), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n489_), .A2(new_n490_), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n520_), .B(new_n637_), .C1(new_n611_), .C2(new_n612_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT39), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(new_n639_), .A3(G8gat), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(KEYINPUT103), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT103), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n638_), .A2(new_n642_), .A3(new_n639_), .A4(G8gat), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n638_), .A2(G8gat), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT39), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n641_), .A2(new_n643_), .A3(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT104), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n629_), .A2(new_n525_), .A3(new_n637_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n646_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n647_), .B1(new_n646_), .B2(new_n648_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n636_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n646_), .A2(new_n648_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT104), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n646_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n653_), .A2(KEYINPUT40), .A3(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n651_), .A2(new_n655_), .ZN(G1325gat));
  AND2_X1   g455(.A1(new_n511_), .A2(new_n513_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n614_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(G15gat), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n659_), .A2(KEYINPUT41), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(KEYINPUT41), .ZN(new_n661_));
  INV_X1    g460(.A(G15gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n629_), .A2(new_n662_), .A3(new_n657_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n660_), .A2(new_n661_), .A3(new_n663_), .ZN(G1326gat));
  INV_X1    g463(.A(G22gat), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n665_), .B1(new_n614_), .B2(new_n482_), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n666_), .B(KEYINPUT42), .Z(new_n667_));
  NAND3_X1  g466(.A1(new_n629_), .A2(new_n665_), .A3(new_n482_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1327gat));
  NAND2_X1  g468(.A1(new_n596_), .A2(new_n627_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT105), .Z(new_n671_));
  AOI21_X1  g470(.A(new_n657_), .B1(new_n480_), .B2(new_n491_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n626_), .B1(new_n672_), .B2(new_n518_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT106), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(new_n674_), .A3(KEYINPUT43), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n676_), .B(new_n626_), .C1(new_n672_), .C2(new_n518_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n674_), .B1(new_n673_), .B2(KEYINPUT43), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n671_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n671_), .B(KEYINPUT44), .C1(new_n678_), .C2(new_n679_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(new_n615_), .A3(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(G29gat), .ZN(new_n685_));
  INV_X1    g484(.A(new_n289_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n686_), .A2(new_n610_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n621_), .A2(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n483_), .A2(G29gat), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT107), .Z(new_n690_));
  OAI21_X1  g489(.A(new_n685_), .B1(new_n688_), .B2(new_n690_), .ZN(G1328gat));
  NAND3_X1  g490(.A1(new_n682_), .A2(new_n637_), .A3(new_n683_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(G36gat), .ZN(new_n693_));
  INV_X1    g492(.A(new_n637_), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n688_), .A2(G36gat), .A3(new_n694_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT45), .Z(new_n696_));
  NAND2_X1  g495(.A1(new_n693_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT46), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n693_), .A2(KEYINPUT46), .A3(new_n696_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1329gat));
  NAND4_X1  g500(.A1(new_n682_), .A2(G43gat), .A3(new_n657_), .A4(new_n683_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(KEYINPUT108), .B(G43gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n703_), .B1(new_n688_), .B2(new_n514_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g505(.A1(new_n688_), .A2(new_n348_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n707_), .A2(G50gat), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n682_), .A2(G50gat), .A3(new_n482_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n709_), .B2(new_n683_), .ZN(G1331gat));
  NAND2_X1  g509(.A1(new_n515_), .A2(new_n519_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n711_), .A2(KEYINPUT109), .A3(new_n547_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n619_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(KEYINPUT109), .B1(new_n711_), .B2(new_n547_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(new_n628_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n351_), .B1(new_n717_), .B2(new_n483_), .ZN(new_n718_));
  NOR4_X1   g517(.A1(new_n521_), .A2(new_n627_), .A3(new_n546_), .A4(new_n619_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n719_), .A2(G57gat), .A3(new_n615_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT110), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n721_), .B(new_n722_), .ZN(G1332gat));
  INV_X1    g522(.A(G64gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n724_), .B1(new_n719_), .B2(new_n637_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT48), .Z(new_n726_));
  NAND2_X1  g525(.A1(new_n637_), .A2(new_n724_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n717_), .B2(new_n727_), .ZN(G1333gat));
  INV_X1    g527(.A(G71gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n729_), .B1(new_n719_), .B2(new_n657_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(KEYINPUT111), .B(KEYINPUT49), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n730_), .B(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n657_), .A2(new_n729_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n717_), .B2(new_n733_), .ZN(G1334gat));
  INV_X1    g533(.A(G78gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n735_), .B1(new_n719_), .B2(new_n482_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT50), .Z(new_n737_));
  NAND2_X1  g536(.A1(new_n482_), .A2(new_n735_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n737_), .B1(new_n717_), .B2(new_n738_), .ZN(G1335gat));
  NOR3_X1   g538(.A1(new_n619_), .A2(new_n610_), .A3(new_n546_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n740_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G85gat), .B1(new_n741_), .B2(new_n483_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n716_), .A2(new_n687_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n615_), .A2(new_n203_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n742_), .B1(new_n743_), .B2(new_n744_), .ZN(G1336gat));
  OAI21_X1  g544(.A(new_n204_), .B1(new_n743_), .B2(new_n694_), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n746_), .A2(KEYINPUT112), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(KEYINPUT112), .ZN(new_n748_));
  OR3_X1    g547(.A1(new_n741_), .A2(new_n211_), .A3(new_n694_), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n747_), .A2(new_n748_), .A3(new_n749_), .ZN(G1337gat));
  INV_X1    g549(.A(new_n743_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n657_), .A2(new_n217_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n657_), .B(new_n740_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n754_));
  AOI22_X1  g553(.A1(new_n751_), .A2(new_n753_), .B1(G99gat), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT113), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n755_), .A2(new_n756_), .A3(KEYINPUT51), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n756_), .A2(KEYINPUT51), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n756_), .A2(KEYINPUT51), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n755_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n757_), .A2(new_n760_), .ZN(G1338gat));
  NAND3_X1  g560(.A1(new_n751_), .A2(new_n218_), .A3(new_n482_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n482_), .B(new_n740_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n763_), .A2(new_n764_), .A3(G106gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n763_), .B2(G106gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n762_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT53), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n762_), .B(new_n769_), .C1(new_n765_), .C2(new_n766_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(G1339gat));
  NOR2_X1   g570(.A1(new_n624_), .A2(new_n625_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n772_), .A2(new_n610_), .A3(new_n592_), .A4(new_n547_), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT54), .Z(new_n774_));
  NAND2_X1  g573(.A1(new_n585_), .A2(new_n546_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT114), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n585_), .A2(new_n546_), .A3(KEYINPUT114), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n569_), .A2(new_n780_), .ZN(new_n781_));
  AOI22_X1  g580(.A1(new_n563_), .A2(new_n565_), .B1(new_n250_), .B2(new_n554_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n782_), .A2(KEYINPUT55), .A3(new_n567_), .A4(new_n561_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT72), .B1(new_n570_), .B2(new_n562_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n559_), .A2(new_n564_), .A3(KEYINPUT12), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n568_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n558_), .A2(new_n560_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n578_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n781_), .A2(new_n783_), .A3(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n583_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT56), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n789_), .A2(KEYINPUT56), .A3(new_n583_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n779_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n535_), .A2(new_n536_), .A3(new_n533_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n542_), .B(new_n795_), .C1(new_n531_), .C2(new_n533_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n544_), .A2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n797_), .B1(new_n589_), .B2(new_n585_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n686_), .B1(new_n794_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n585_), .A2(new_n544_), .A3(new_n796_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n803_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n772_), .B1(new_n804_), .B2(KEYINPUT58), .ZN(new_n805_));
  INV_X1    g604(.A(new_n803_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n789_), .A2(KEYINPUT56), .A3(new_n583_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT56), .B1(new_n789_), .B2(new_n583_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n806_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT58), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  AOI22_X1  g610(.A1(new_n799_), .A2(new_n800_), .B1(new_n805_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n802_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n774_), .B1(new_n813_), .B2(new_n627_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n517_), .A2(new_n514_), .A3(new_n483_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n814_), .A2(new_n547_), .A3(new_n816_), .ZN(new_n817_));
  OR2_X1    g616(.A1(new_n817_), .A2(G113gat), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n818_), .A2(KEYINPUT115), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(KEYINPUT115), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n821_));
  OAI211_X1 g620(.A(KEYINPUT58), .B(new_n806_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n626_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n792_), .A2(new_n793_), .ZN(new_n824_));
  AOI21_X1  g623(.A(KEYINPUT58), .B1(new_n824_), .B2(new_n806_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n585_), .A2(KEYINPUT114), .A3(new_n546_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT114), .B1(new_n585_), .B2(new_n546_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n798_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT57), .B1(new_n832_), .B2(new_n686_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n821_), .B1(new_n826_), .B2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n811_), .A2(new_n626_), .A3(new_n822_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n289_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n835_), .B(KEYINPUT116), .C1(KEYINPUT57), .C2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n834_), .A2(new_n802_), .A3(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n774_), .B1(new_n838_), .B2(new_n627_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n816_), .A2(KEYINPUT59), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n814_), .A2(new_n816_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n842_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n546_), .A2(G113gat), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(KEYINPUT117), .ZN(new_n848_));
  AOI22_X1  g647(.A1(new_n819_), .A2(new_n820_), .B1(new_n846_), .B2(new_n848_), .ZN(G1340gat));
  XOR2_X1   g648(.A(KEYINPUT118), .B(G120gat), .Z(new_n850_));
  OAI21_X1  g649(.A(new_n850_), .B1(new_n619_), .B2(KEYINPUT60), .ZN(new_n851_));
  OAI22_X1  g650(.A1(new_n851_), .A2(KEYINPUT119), .B1(KEYINPUT60), .B2(new_n850_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(KEYINPUT119), .B2(new_n851_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n843_), .A2(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n845_), .A2(new_n619_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n850_), .ZN(G1341gat));
  OAI21_X1  g655(.A(G127gat), .B1(new_n845_), .B2(new_n627_), .ZN(new_n857_));
  INV_X1    g656(.A(G127gat), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n843_), .A2(new_n858_), .A3(new_n610_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(G1342gat));
  OAI21_X1  g659(.A(G134gat), .B1(new_n845_), .B2(new_n772_), .ZN(new_n861_));
  INV_X1    g660(.A(G134gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n843_), .A2(new_n862_), .A3(new_n290_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n863_), .ZN(G1343gat));
  NAND2_X1  g663(.A1(new_n514_), .A2(new_n482_), .ZN(new_n865_));
  NOR4_X1   g664(.A1(new_n814_), .A2(new_n483_), .A3(new_n637_), .A4(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n546_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n713_), .ZN(new_n869_));
  XOR2_X1   g668(.A(KEYINPUT120), .B(G148gat), .Z(new_n870_));
  XNOR2_X1  g669(.A(new_n869_), .B(new_n870_), .ZN(G1345gat));
  NAND2_X1  g670(.A1(new_n866_), .A2(new_n610_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT61), .B(G155gat), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1346gat));
  INV_X1    g673(.A(G162gat), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n866_), .A2(new_n875_), .A3(new_n290_), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n866_), .A2(new_n626_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n877_), .B2(new_n875_), .ZN(G1347gat));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n657_), .A2(new_n483_), .A3(new_n637_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n880_), .A2(new_n482_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n879_), .B1(new_n839_), .B2(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n801_), .B1(new_n812_), .B2(KEYINPUT116), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n610_), .B1(new_n884_), .B2(new_n834_), .ZN(new_n885_));
  OAI211_X1 g684(.A(KEYINPUT122), .B(new_n881_), .C1(new_n885_), .C2(new_n774_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n883_), .A2(new_n886_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n887_), .A2(new_n546_), .A3(new_n429_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n839_), .A2(new_n547_), .A3(new_n882_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT62), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n890_), .A2(KEYINPUT121), .A3(new_n891_), .A4(G169gat), .ZN(new_n892_));
  INV_X1    g691(.A(G169gat), .ZN(new_n893_));
  OAI21_X1  g692(.A(KEYINPUT62), .B1(new_n889_), .B2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n889_), .A2(new_n893_), .ZN(new_n896_));
  AOI21_X1  g695(.A(KEYINPUT121), .B1(new_n896_), .B2(new_n891_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n888_), .B1(new_n895_), .B2(new_n897_), .ZN(G1348gat));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n899_));
  AOI21_X1  g698(.A(G176gat), .B1(new_n887_), .B2(new_n713_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n814_), .A2(new_n482_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n880_), .A2(new_n414_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n901_), .A2(new_n713_), .A3(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n899_), .B1(new_n900_), .B2(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n619_), .B1(new_n883_), .B2(new_n886_), .ZN(new_n906_));
  OAI211_X1 g705(.A(KEYINPUT123), .B(new_n903_), .C1(new_n906_), .C2(G176gat), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n905_), .A2(new_n907_), .ZN(G1349gat));
  NOR4_X1   g707(.A1(new_n814_), .A2(new_n627_), .A3(new_n482_), .A4(new_n880_), .ZN(new_n909_));
  OR2_X1    g708(.A1(new_n909_), .A2(KEYINPUT124), .ZN(new_n910_));
  AOI21_X1  g709(.A(G183gat), .B1(new_n909_), .B2(KEYINPUT124), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n627_), .A2(new_n408_), .ZN(new_n912_));
  AOI22_X1  g711(.A1(new_n910_), .A2(new_n911_), .B1(new_n887_), .B2(new_n912_), .ZN(G1350gat));
  INV_X1    g712(.A(new_n887_), .ZN(new_n914_));
  OAI21_X1  g713(.A(G190gat), .B1(new_n914_), .B2(new_n772_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n887_), .A2(new_n407_), .A3(new_n290_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1351gat));
  NOR3_X1   g716(.A1(new_n865_), .A2(new_n615_), .A3(new_n694_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n814_), .A2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n546_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g721(.A1(new_n920_), .A2(new_n713_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g723(.A(new_n627_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n920_), .A2(new_n925_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(KEYINPUT125), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(KEYINPUT126), .ZN(new_n929_));
  XOR2_X1   g728(.A(new_n926_), .B(new_n929_), .Z(G1354gat));
  INV_X1    g729(.A(G218gat), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n920_), .A2(new_n931_), .A3(new_n290_), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n814_), .A2(new_n772_), .A3(new_n919_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n931_), .B2(new_n933_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


