//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 1 0 0 1 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 1 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n913_, new_n915_, new_n917_, new_n918_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n946_, new_n947_, new_n948_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n955_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n965_, new_n966_;
  INV_X1    g000(.A(G169gat), .ZN(new_n202_));
  INV_X1    g001(.A(G176gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205_));
  AND3_X1   g004(.A1(new_n204_), .A2(KEYINPUT24), .A3(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n204_), .A2(KEYINPUT24), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G183gat), .ZN(new_n209_));
  INV_X1    g008(.A(G190gat), .ZN(new_n210_));
  NOR3_X1   g009(.A1(new_n209_), .A2(new_n210_), .A3(KEYINPUT23), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT23), .B1(new_n209_), .B2(new_n210_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT25), .B(G183gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT26), .B(G190gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n208_), .A2(new_n214_), .A3(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT22), .B(G169gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT95), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n219_), .B(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n205_), .B1(new_n221_), .B2(G176gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n213_), .A2(KEYINPUT83), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT83), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n224_), .B(KEYINPUT23), .C1(new_n209_), .C2(new_n210_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n211_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n218_), .B1(new_n222_), .B2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G197gat), .B(G204gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT21), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n231_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G211gat), .B(G218gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT92), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n234_), .A2(new_n235_), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n232_), .B(new_n233_), .C1(new_n237_), .C2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n238_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n230_), .A2(new_n231_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(new_n241_), .A3(new_n236_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n239_), .A2(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT20), .B1(new_n229_), .B2(new_n243_), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n239_), .A2(new_n242_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(KEYINPUT81), .B(G190gat), .Z(new_n248_));
  INV_X1    g047(.A(KEYINPUT26), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n250_), .A2(KEYINPUT82), .A3(new_n215_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT82), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT81), .B(G190gat), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n246_), .B1(new_n253_), .B2(KEYINPUT26), .ZN(new_n254_));
  INV_X1    g053(.A(new_n215_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n252_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n226_), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n251_), .A2(new_n256_), .A3(new_n257_), .A4(new_n208_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n214_), .B1(G183gat), .B2(new_n253_), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT84), .B1(new_n202_), .B2(KEYINPUT22), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n203_), .B(new_n260_), .C1(new_n219_), .C2(KEYINPUT84), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n259_), .A2(new_n205_), .A3(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n245_), .B1(new_n258_), .B2(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n244_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT96), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G226gat), .A2(G233gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT19), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n264_), .A2(new_n265_), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n258_), .A2(new_n262_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(new_n243_), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n245_), .B(new_n218_), .C1(new_n228_), .C2(new_n222_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n271_), .A2(new_n272_), .A3(KEYINPUT20), .A4(new_n268_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT96), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT20), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n275_), .B1(new_n229_), .B2(new_n243_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n245_), .A2(new_n258_), .A3(new_n262_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n268_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n269_), .B1(new_n274_), .B2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G8gat), .B(G36gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT18), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G64gat), .B(G92gat), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n281_), .B(new_n282_), .Z(new_n283_));
  NAND2_X1  g082(.A1(new_n279_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n276_), .A2(new_n277_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n267_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n286_), .A2(KEYINPUT96), .A3(new_n273_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n283_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n287_), .A2(new_n288_), .A3(new_n269_), .ZN(new_n289_));
  AOI21_X1  g088(.A(KEYINPUT27), .B1(new_n284_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT99), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n291_), .B1(new_n279_), .B2(new_n283_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n229_), .A2(new_n243_), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n293_), .A2(new_n277_), .A3(KEYINPUT20), .A4(new_n268_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT98), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT98), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n276_), .A2(new_n296_), .A3(new_n268_), .A4(new_n277_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n267_), .B1(new_n244_), .B2(new_n263_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n295_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n288_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT27), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n292_), .A2(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n288_), .B1(new_n287_), .B2(new_n269_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n291_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n290_), .B1(new_n302_), .B2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT28), .B(G22gat), .ZN(new_n306_));
  INV_X1    g105(.A(G50gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT90), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311_));
  OR2_X1    g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312_));
  AOI21_X1  g111(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT89), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT3), .ZN(new_n315_));
  INV_X1    g114(.A(G141gat), .ZN(new_n316_));
  INV_X1    g115(.A(G148gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT2), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G141gat), .A2(G148gat), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n318_), .B(new_n319_), .C1(new_n320_), .C2(new_n321_), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n311_), .B(new_n312_), .C1(new_n314_), .C2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n316_), .A2(new_n317_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n311_), .A2(KEYINPUT1), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(new_n312_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n311_), .A2(KEYINPUT1), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n321_), .B(new_n324_), .C1(new_n326_), .C2(new_n327_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n323_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT29), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n310_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n323_), .A2(new_n328_), .ZN(new_n332_));
  NOR3_X1   g131(.A1(new_n332_), .A2(KEYINPUT90), .A3(KEYINPUT29), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n309_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n329_), .A2(new_n310_), .A3(new_n330_), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT90), .B1(new_n332_), .B2(KEYINPUT29), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(new_n308_), .A3(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n334_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G78gat), .B(G106gat), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n332_), .A2(KEYINPUT29), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(new_n243_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(KEYINPUT91), .A2(G233gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(KEYINPUT91), .A2(G233gat), .ZN(new_n345_));
  OAI21_X1  g144(.A(G228gat), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n342_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n341_), .A2(new_n243_), .A3(new_n346_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n340_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n338_), .B1(KEYINPUT93), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n349_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n346_), .B1(new_n341_), .B2(new_n243_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n339_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n348_), .A2(new_n349_), .A3(new_n340_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT93), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n338_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT94), .ZN(new_n359_));
  AOI22_X1  g158(.A1(new_n351_), .A2(new_n357_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n358_), .A2(new_n359_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G1gat), .B(G29gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT97), .B(G85gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT0), .B(G57gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT4), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G127gat), .B(G134gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G113gat), .B(G120gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT85), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n371_), .A2(new_n372_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT86), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(new_n332_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n373_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n323_), .B(new_n328_), .C1(new_n379_), .C2(new_n376_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n370_), .B1(new_n378_), .B2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT86), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n376_), .B(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n383_), .A2(new_n374_), .ZN(new_n384_));
  AOI21_X1  g183(.A(KEYINPUT4), .B1(new_n384_), .B2(new_n332_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G225gat), .A2(G233gat), .ZN(new_n386_));
  NOR3_X1   g185(.A1(new_n381_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n378_), .A2(new_n380_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n386_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n369_), .B1(new_n387_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n388_), .A2(KEYINPUT4), .ZN(new_n392_));
  INV_X1    g191(.A(new_n386_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n385_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n392_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n395_), .A2(new_n368_), .A3(new_n389_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n391_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT31), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n384_), .B(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT87), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT88), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G71gat), .B(G99gat), .ZN(new_n403_));
  INV_X1    g202(.A(G43gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n270_), .B(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G227gat), .A2(G233gat), .ZN(new_n407_));
  INV_X1    g206(.A(G15gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT30), .ZN(new_n410_));
  OR2_X1    g209(.A1(new_n406_), .A2(new_n410_), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n399_), .A2(KEYINPUT87), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n406_), .A2(new_n410_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n402_), .A2(new_n411_), .A3(new_n412_), .A4(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n400_), .B(KEYINPUT88), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n411_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n397_), .B1(new_n414_), .B2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n305_), .A2(new_n363_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n393_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n368_), .B1(new_n388_), .B2(new_n386_), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT33), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n391_), .ZN(new_n423_));
  OAI211_X1 g222(.A(KEYINPUT33), .B(new_n369_), .C1(new_n387_), .C2(new_n390_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n284_), .A2(new_n423_), .A3(new_n289_), .A4(new_n424_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n283_), .A2(KEYINPUT32), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n299_), .A2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n273_), .A2(KEYINPUT96), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n265_), .B1(new_n264_), .B2(new_n268_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n428_), .B1(new_n429_), .B2(new_n286_), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n397_), .B(new_n427_), .C1(new_n430_), .C2(new_n426_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n362_), .B1(new_n425_), .B2(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n397_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n432_), .B1(new_n305_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n414_), .A2(new_n417_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n419_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G232gat), .A2(G233gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT34), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT35), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G99gat), .A2(G106gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT6), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT6), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n444_), .A2(G99gat), .A3(G106gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT10), .B(G99gat), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n446_), .B1(new_n447_), .B2(G106gat), .ZN(new_n448_));
  OAI211_X1 g247(.A(KEYINPUT64), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G85gat), .A2(G92gat), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n449_), .B(new_n451_), .C1(KEYINPUT64), .C2(KEYINPUT9), .ZN(new_n452_));
  INV_X1    g251(.A(G85gat), .ZN(new_n453_));
  INV_X1    g252(.A(G92gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n455_), .A2(KEYINPUT64), .A3(KEYINPUT9), .A4(new_n450_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n452_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT65), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n448_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n452_), .A2(KEYINPUT65), .A3(new_n456_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(G85gat), .A2(G92gat), .ZN(new_n462_));
  NOR3_X1   g261(.A1(new_n451_), .A2(new_n462_), .A3(KEYINPUT8), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n443_), .A2(new_n445_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT7), .ZN(new_n465_));
  INV_X1    g264(.A(G99gat), .ZN(new_n466_));
  INV_X1    g265(.A(G106gat), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n463_), .B1(new_n464_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT66), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n446_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT66), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(new_n474_), .A3(new_n463_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n472_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT8), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n446_), .A2(KEYINPUT67), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT67), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n443_), .A2(new_n445_), .A3(new_n479_), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n468_), .A2(new_n469_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n478_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n451_), .A2(new_n462_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n477_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n461_), .B1(new_n476_), .B2(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(G29gat), .B(G36gat), .Z(new_n486_));
  XOR2_X1   g285(.A(G43gat), .B(G50gat), .Z(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G29gat), .B(G36gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G43gat), .B(G50gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  OAI22_X1  g292(.A1(new_n485_), .A2(new_n493_), .B1(KEYINPUT35), .B2(new_n438_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n492_), .B(KEYINPUT15), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n485_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT71), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n485_), .A2(KEYINPUT71), .A3(new_n495_), .ZN(new_n499_));
  AOI211_X1 g298(.A(new_n441_), .B(new_n494_), .C1(new_n498_), .C2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n441_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n498_), .A2(new_n499_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n494_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n501_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT73), .B1(new_n500_), .B2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G190gat), .B(G218gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G134gat), .B(G162gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n508_), .B(KEYINPUT36), .Z(new_n509_));
  INV_X1    g308(.A(new_n499_), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT71), .B1(new_n485_), .B2(new_n495_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n503_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n441_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT73), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n502_), .A2(new_n501_), .A3(new_n503_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n505_), .A2(new_n509_), .A3(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n508_), .A2(KEYINPUT36), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n513_), .A2(new_n515_), .A3(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n436_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT70), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G57gat), .B(G64gat), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n523_), .A2(KEYINPUT11), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(KEYINPUT11), .ZN(new_n525_));
  XOR2_X1   g324(.A(G71gat), .B(G78gat), .Z(new_n526_));
  NAND3_X1  g325(.A1(new_n524_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n525_), .A2(new_n526_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n461_), .B(new_n529_), .C1(new_n476_), .C2(new_n484_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G230gat), .A2(G233gat), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(KEYINPUT69), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n483_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n479_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n534_), .A2(new_n470_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n533_), .B1(new_n535_), .B2(new_n480_), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n472_), .B(new_n475_), .C1(new_n536_), .C2(new_n477_), .ZN(new_n537_));
  AOI211_X1 g336(.A(KEYINPUT12), .B(new_n529_), .C1(new_n537_), .C2(new_n461_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT12), .ZN(new_n539_));
  INV_X1    g338(.A(new_n529_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n539_), .B1(new_n485_), .B2(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n532_), .B1(new_n538_), .B2(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(KEYINPUT69), .B1(new_n530_), .B2(new_n531_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n522_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n473_), .A2(new_n474_), .A3(new_n463_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n474_), .B1(new_n473_), .B2(new_n463_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n443_), .A2(new_n445_), .A3(new_n479_), .ZN(new_n548_));
  NOR3_X1   g347(.A1(new_n548_), .A2(new_n534_), .A3(new_n470_), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT8), .B1(new_n549_), .B2(new_n533_), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n547_), .A2(new_n550_), .B1(new_n460_), .B2(new_n459_), .ZN(new_n551_));
  OAI21_X1  g350(.A(KEYINPUT12), .B1(new_n551_), .B2(new_n529_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n485_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n543_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n554_), .A2(KEYINPUT70), .A3(new_n555_), .A4(new_n532_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n531_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n485_), .A2(KEYINPUT68), .A3(new_n540_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT68), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n559_), .B1(new_n551_), .B2(new_n529_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n530_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n557_), .B(new_n558_), .C1(new_n560_), .C2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n544_), .A2(new_n556_), .A3(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G120gat), .B(G148gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT5), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G176gat), .B(G204gat), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n565_), .B(new_n566_), .Z(new_n567_));
  NAND2_X1  g366(.A1(new_n563_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n567_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n544_), .A2(new_n556_), .A3(new_n562_), .A4(new_n569_), .ZN(new_n570_));
  AND3_X1   g369(.A1(new_n568_), .A2(KEYINPUT13), .A3(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(KEYINPUT13), .B1(new_n568_), .B2(new_n570_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G15gat), .B(G22gat), .ZN(new_n574_));
  INV_X1    g373(.A(G1gat), .ZN(new_n575_));
  INV_X1    g374(.A(G8gat), .ZN(new_n576_));
  OAI21_X1  g375(.A(KEYINPUT14), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n574_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G1gat), .B(G8gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(new_n529_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G127gat), .B(G155gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT16), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G183gat), .B(G211gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n587_), .B(KEYINPUT17), .Z(new_n588_));
  NAND2_X1  g387(.A1(new_n583_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(KEYINPUT17), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n582_), .B(new_n540_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n590_), .B1(new_n591_), .B2(KEYINPUT74), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n592_), .B1(KEYINPUT74), .B2(new_n591_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n593_), .A2(KEYINPUT75), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(KEYINPUT75), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n589_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT76), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n492_), .B(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n580_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n492_), .B(KEYINPUT76), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(new_n580_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G229gat), .A2(G233gat), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n495_), .A2(new_n580_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n605_), .B(KEYINPUT77), .Z(new_n609_));
  NAND3_X1  g408(.A1(new_n601_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(G113gat), .B(G141gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT79), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G169gat), .B(G197gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT80), .ZN(new_n615_));
  AOI22_X1  g414(.A1(new_n607_), .A2(new_n610_), .B1(KEYINPUT78), .B2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n607_), .A2(KEYINPUT78), .A3(new_n610_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(KEYINPUT80), .ZN(new_n618_));
  INV_X1    g417(.A(new_n614_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n616_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n573_), .A2(new_n597_), .A3(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n521_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT101), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n397_), .ZN(new_n625_));
  OAI21_X1  g424(.A(G1gat), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n573_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT72), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n628_), .B(new_n509_), .C1(new_n500_), .C2(new_n504_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(new_n519_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n513_), .A2(new_n515_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n628_), .B1(new_n631_), .B2(new_n509_), .ZN(new_n632_));
  OAI21_X1  g431(.A(KEYINPUT37), .B1(new_n630_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT37), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n517_), .A2(new_n634_), .A3(new_n519_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n596_), .B1(new_n633_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT27), .ZN(new_n638_));
  INV_X1    g437(.A(new_n289_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n638_), .B1(new_n639_), .B2(new_n303_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n304_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n638_), .B1(new_n299_), .B2(new_n288_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n642_), .B1(new_n303_), .B2(new_n291_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n640_), .B(new_n433_), .C1(new_n641_), .C2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n425_), .A2(new_n431_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(new_n363_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n435_), .B1(new_n644_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n292_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n648_), .A2(new_n304_), .A3(new_n642_), .ZN(new_n649_));
  AND4_X1   g448(.A1(new_n363_), .A2(new_n649_), .A3(new_n418_), .A4(new_n640_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n620_), .B1(new_n647_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OAI211_X1 g452(.A(KEYINPUT100), .B(new_n620_), .C1(new_n647_), .C2(new_n650_), .ZN(new_n654_));
  AOI211_X1 g453(.A(new_n627_), .B(new_n637_), .C1(new_n653_), .C2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(new_n575_), .A3(new_n397_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT38), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n657_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n626_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT102), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n626_), .A2(new_n658_), .A3(KEYINPUT102), .A4(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1324gat));
  INV_X1    g463(.A(new_n305_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n576_), .B1(new_n622_), .B2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n666_), .B(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n655_), .A2(new_n576_), .A3(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT40), .Z(G1325gat));
  AOI21_X1  g470(.A(new_n408_), .B1(new_n623_), .B2(new_n435_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n673_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n655_), .A2(new_n408_), .A3(new_n435_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT104), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n674_), .A2(new_n675_), .A3(new_n677_), .ZN(G1326gat));
  INV_X1    g477(.A(G22gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n679_), .B1(new_n623_), .B2(new_n362_), .ZN(new_n680_));
  XOR2_X1   g479(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n655_), .A2(new_n679_), .A3(new_n362_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1327gat));
  INV_X1    g483(.A(new_n520_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(new_n596_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n627_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  OR3_X1    g489(.A1(new_n690_), .A2(G29gat), .A3(new_n625_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n620_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n627_), .A2(new_n692_), .A3(new_n597_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n633_), .A2(new_n635_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n436_), .B2(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n694_), .B(new_n695_), .C1(new_n647_), .C2(new_n650_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n693_), .B1(new_n696_), .B2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n695_), .B1(new_n647_), .B2(new_n650_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT43), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(new_n697_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n704_), .A2(KEYINPUT44), .A3(new_n693_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n701_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(new_n397_), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n707_), .A2(KEYINPUT106), .A3(G29gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT106), .B1(new_n707_), .B2(G29gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n691_), .B1(new_n708_), .B2(new_n709_), .ZN(G1328gat));
  NAND3_X1  g509(.A1(new_n701_), .A2(new_n665_), .A3(new_n705_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(G36gat), .ZN(new_n712_));
  INV_X1    g511(.A(G36gat), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n665_), .A2(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(KEYINPUT107), .B1(new_n690_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT45), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n689_), .A2(new_n717_), .A3(new_n713_), .A4(new_n665_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n715_), .A2(new_n716_), .A3(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n716_), .B1(new_n715_), .B2(new_n718_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n712_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT46), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  OAI211_X1 g522(.A(KEYINPUT46), .B(new_n712_), .C1(new_n719_), .C2(new_n720_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1329gat));
  INV_X1    g524(.A(new_n435_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n726_), .A2(new_n404_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n701_), .A2(new_n705_), .A3(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT100), .B1(new_n436_), .B2(new_n620_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n654_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n435_), .B(new_n687_), .C1(new_n729_), .C2(new_n730_), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n731_), .A2(KEYINPUT108), .A3(new_n404_), .ZN(new_n732_));
  AOI21_X1  g531(.A(KEYINPUT108), .B1(new_n731_), .B2(new_n404_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n728_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT110), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT110), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n728_), .B(new_n736_), .C1(new_n732_), .C2(new_n733_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n735_), .A2(new_n737_), .A3(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n735_), .B2(new_n737_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1330gat));
  AOI21_X1  g540(.A(G50gat), .B1(new_n689_), .B2(new_n362_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n363_), .A2(new_n307_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n706_), .B2(new_n743_), .ZN(G1331gat));
  INV_X1    g543(.A(new_n521_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n745_), .A2(new_n692_), .A3(new_n627_), .A4(new_n597_), .ZN(new_n746_));
  OAI21_X1  g545(.A(G57gat), .B1(new_n746_), .B2(new_n625_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n436_), .A2(new_n692_), .ZN(new_n748_));
  OAI21_X1  g547(.A(KEYINPUT111), .B1(new_n637_), .B2(new_n573_), .ZN(new_n749_));
  OR3_X1    g548(.A1(new_n637_), .A2(KEYINPUT111), .A3(new_n573_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n748_), .A2(new_n749_), .A3(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(G57gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(new_n752_), .A3(new_n397_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n747_), .A2(new_n753_), .ZN(G1332gat));
  OAI21_X1  g553(.A(G64gat), .B1(new_n746_), .B2(new_n305_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT48), .ZN(new_n756_));
  INV_X1    g555(.A(G64gat), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n751_), .A2(new_n757_), .A3(new_n665_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1333gat));
  OAI21_X1  g558(.A(G71gat), .B1(new_n746_), .B2(new_n726_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT49), .ZN(new_n761_));
  INV_X1    g560(.A(G71gat), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n751_), .A2(new_n762_), .A3(new_n435_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1334gat));
  OAI21_X1  g563(.A(G78gat), .B1(new_n746_), .B2(new_n363_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT50), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n363_), .A2(G78gat), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT112), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n751_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n766_), .A2(new_n769_), .ZN(G1335gat));
  NOR3_X1   g569(.A1(new_n573_), .A2(new_n597_), .A3(new_n620_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n772_), .B1(new_n703_), .B2(new_n697_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(G85gat), .B1(new_n774_), .B2(new_n625_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n686_), .A2(new_n573_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n748_), .A2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(new_n453_), .A3(new_n397_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n775_), .A2(new_n779_), .ZN(G1336gat));
  OAI21_X1  g579(.A(G92gat), .B1(new_n774_), .B2(new_n305_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n778_), .A2(new_n454_), .A3(new_n665_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(G1337gat));
  OAI21_X1  g582(.A(G99gat), .B1(new_n774_), .B2(new_n726_), .ZN(new_n784_));
  OR2_X1    g583(.A1(new_n726_), .A2(new_n447_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n784_), .B1(new_n777_), .B2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n787_));
  XOR2_X1   g586(.A(new_n786_), .B(new_n787_), .Z(G1338gat));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n704_), .A2(new_n789_), .A3(new_n362_), .A4(new_n771_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(G106gat), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n789_), .B1(new_n773_), .B2(new_n362_), .ZN(new_n792_));
  OAI21_X1  g591(.A(KEYINPUT115), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n704_), .A2(new_n362_), .A3(new_n771_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT114), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n795_), .A2(new_n796_), .A3(G106gat), .A4(new_n790_), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n793_), .A2(KEYINPUT52), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799_));
  OAI211_X1 g598(.A(KEYINPUT115), .B(new_n799_), .C1(new_n791_), .C2(new_n792_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n778_), .A2(new_n467_), .A3(new_n362_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(KEYINPUT53), .B1(new_n798_), .B2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n793_), .A2(KEYINPUT52), .A3(new_n797_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n804_), .A2(new_n805_), .A3(new_n800_), .A4(new_n801_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n803_), .A2(new_n806_), .ZN(G1339gat));
  NAND2_X1  g606(.A1(new_n568_), .A2(new_n570_), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n607_), .A2(new_n610_), .A3(new_n614_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n601_), .A2(new_n603_), .A3(new_n609_), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n601_), .A2(new_n608_), .A3(KEYINPUT118), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT118), .B1(new_n601_), .B2(new_n608_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n810_), .B1(new_n813_), .B2(new_n609_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n809_), .B1(new_n814_), .B2(new_n619_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n808_), .A2(new_n815_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n570_), .A2(new_n620_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n544_), .A2(new_n818_), .A3(new_n556_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n554_), .A2(KEYINPUT55), .A3(new_n555_), .A4(new_n532_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n530_), .B1(new_n538_), .B2(new_n541_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n557_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n820_), .A2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n569_), .B1(new_n819_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT56), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT117), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n817_), .B1(new_n824_), .B2(new_n827_), .ZN(new_n828_));
  AOI211_X1 g627(.A(new_n569_), .B(new_n826_), .C1(new_n819_), .C2(new_n823_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n816_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n830_), .A2(KEYINPUT57), .A3(new_n520_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n819_), .A2(new_n823_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n833_), .A2(new_n825_), .A3(new_n567_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n815_), .A2(new_n570_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n824_), .A2(new_n825_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n832_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n833_), .A2(new_n567_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT56), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n840_), .A2(KEYINPUT58), .A3(new_n834_), .A4(new_n835_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n838_), .A2(new_n695_), .A3(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT57), .B1(new_n830_), .B2(new_n520_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n831_), .B(new_n842_), .C1(new_n843_), .C2(KEYINPUT119), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT119), .ZN(new_n845_));
  AOI211_X1 g644(.A(new_n845_), .B(KEYINPUT57), .C1(new_n830_), .C2(new_n520_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n596_), .B1(new_n844_), .B2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n636_), .A2(new_n692_), .A3(new_n573_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n850_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n636_), .A2(new_n692_), .A3(new_n573_), .A4(new_n849_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n847_), .A2(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n665_), .A2(new_n362_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n726_), .A2(new_n625_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n854_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(G113gat), .B1(new_n860_), .B2(new_n620_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n851_), .A2(new_n852_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n830_), .A2(new_n520_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n866_), .A2(new_n831_), .A3(new_n842_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n863_), .B1(new_n867_), .B2(new_n596_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n857_), .A2(KEYINPUT59), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n862_), .B1(new_n868_), .B2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n842_), .A2(new_n831_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n596_), .B1(new_n872_), .B2(new_n843_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n853_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(KEYINPUT120), .A3(new_n869_), .ZN(new_n875_));
  AOI22_X1  g674(.A1(new_n859_), .A2(KEYINPUT59), .B1(new_n871_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(G113gat), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n620_), .A2(KEYINPUT121), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n878_), .B1(new_n879_), .B2(G113gat), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n861_), .B1(new_n876_), .B2(new_n880_), .ZN(G1340gat));
  AND2_X1   g680(.A1(new_n876_), .A2(new_n627_), .ZN(new_n882_));
  INV_X1    g681(.A(G120gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n573_), .B2(KEYINPUT60), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(KEYINPUT60), .B2(new_n883_), .ZN(new_n885_));
  OAI22_X1  g684(.A1(new_n882_), .A2(new_n883_), .B1(new_n859_), .B2(new_n885_), .ZN(G1341gat));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n887_));
  INV_X1    g686(.A(G127gat), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n888_), .B1(new_n876_), .B2(new_n597_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n859_), .A2(G127gat), .A3(new_n596_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n887_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n866_), .A2(new_n845_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n843_), .A2(KEYINPUT119), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n892_), .A2(new_n893_), .A3(new_n831_), .A4(new_n842_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n863_), .B1(new_n894_), .B2(new_n596_), .ZN(new_n895_));
  OAI21_X1  g694(.A(KEYINPUT59), .B1(new_n895_), .B2(new_n857_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n871_), .A2(new_n875_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n896_), .A2(new_n897_), .A3(new_n597_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(G127gat), .ZN(new_n899_));
  INV_X1    g698(.A(new_n890_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n899_), .A2(KEYINPUT122), .A3(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n891_), .A2(new_n901_), .ZN(G1342gat));
  INV_X1    g701(.A(G134gat), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n903_), .B1(new_n859_), .B2(new_n520_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n905_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n695_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n908_), .A2(new_n903_), .ZN(new_n909_));
  AOI22_X1  g708(.A1(new_n906_), .A2(new_n907_), .B1(new_n876_), .B2(new_n909_), .ZN(G1343gat));
  NOR3_X1   g709(.A1(new_n363_), .A2(new_n435_), .A3(new_n625_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n854_), .A2(new_n305_), .A3(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(new_n692_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(new_n316_), .ZN(G1344gat));
  NOR2_X1   g713(.A1(new_n912_), .A2(new_n573_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(new_n317_), .ZN(G1345gat));
  NOR2_X1   g715(.A1(new_n912_), .A2(new_n596_), .ZN(new_n917_));
  XOR2_X1   g716(.A(KEYINPUT61), .B(G155gat), .Z(new_n918_));
  XNOR2_X1  g717(.A(new_n917_), .B(new_n918_), .ZN(G1346gat));
  OAI21_X1  g718(.A(G162gat), .B1(new_n912_), .B2(new_n908_), .ZN(new_n920_));
  OR2_X1    g719(.A1(new_n520_), .A2(G162gat), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n912_), .B2(new_n921_), .ZN(G1347gat));
  NAND2_X1  g721(.A1(new_n665_), .A2(new_n418_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n362_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n874_), .A2(new_n924_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n925_), .A2(new_n221_), .A3(new_n692_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n925_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n202_), .B1(new_n927_), .B2(new_n620_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n926_), .B1(new_n928_), .B2(KEYINPUT62), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n929_), .B1(KEYINPUT62), .B2(new_n928_), .ZN(G1348gat));
  AOI21_X1  g729(.A(G176gat), .B1(new_n927_), .B2(new_n627_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT124), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n932_), .B1(new_n895_), .B2(new_n362_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n854_), .A2(KEYINPUT124), .A3(new_n363_), .ZN(new_n934_));
  AND2_X1   g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n935_), .ZN(new_n936_));
  NOR3_X1   g735(.A1(new_n923_), .A2(new_n573_), .A3(new_n203_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n931_), .B1(new_n936_), .B2(new_n937_), .ZN(G1349gat));
  NOR3_X1   g737(.A1(new_n925_), .A2(new_n215_), .A3(new_n596_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n597_), .A2(new_n665_), .A3(new_n418_), .ZN(new_n940_));
  OAI21_X1  g739(.A(KEYINPUT125), .B1(new_n935_), .B2(new_n940_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n940_), .B1(new_n933_), .B2(new_n934_), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n943_));
  AOI21_X1  g742(.A(G183gat), .B1(new_n942_), .B2(new_n943_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n939_), .B1(new_n941_), .B2(new_n944_), .ZN(G1350gat));
  OAI21_X1  g744(.A(G190gat), .B1(new_n925_), .B2(new_n908_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n685_), .A2(new_n216_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(KEYINPUT126), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n946_), .B1(new_n925_), .B2(new_n948_), .ZN(G1351gat));
  NOR4_X1   g748(.A1(new_n305_), .A2(new_n363_), .A3(new_n397_), .A4(new_n435_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n854_), .A2(new_n950_), .ZN(new_n951_));
  INV_X1    g750(.A(new_n951_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n952_), .A2(new_n620_), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n953_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g753(.A1(new_n952_), .A2(new_n627_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n955_), .B(G204gat), .ZN(G1353gat));
  OR2_X1    g755(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n957_));
  NAND2_X1  g756(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n958_));
  NAND4_X1  g757(.A1(new_n952_), .A2(new_n597_), .A3(new_n957_), .A4(new_n958_), .ZN(new_n959_));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n960_));
  AND2_X1   g759(.A1(new_n959_), .A2(new_n960_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n951_), .A2(new_n596_), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n959_), .B1(new_n962_), .B2(new_n957_), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n961_), .B1(new_n963_), .B2(KEYINPUT127), .ZN(G1354gat));
  OR3_X1    g763(.A1(new_n951_), .A2(G218gat), .A3(new_n520_), .ZN(new_n965_));
  OAI21_X1  g764(.A(G218gat), .B1(new_n951_), .B2(new_n908_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n965_), .A2(new_n966_), .ZN(G1355gat));
endmodule


