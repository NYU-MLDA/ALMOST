//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 0 0 1 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n626_, new_n627_, new_n628_, new_n629_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n861_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_;
  INV_X1    g000(.A(KEYINPUT102), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT19), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G197gat), .B(G204gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT21), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n206_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  OR3_X1    g009(.A1(new_n205_), .A2(new_n209_), .A3(new_n206_), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n213_));
  INV_X1    g012(.A(G183gat), .ZN(new_n214_));
  INV_X1    g013(.A(G190gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n213_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n216_), .B(new_n217_), .C1(G183gat), .C2(G190gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(G169gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT25), .B(G183gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT26), .B(G190gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT82), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n227_), .B1(G169gat), .B2(G176gat), .ZN(new_n228_));
  NOR3_X1   g027(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n216_), .A2(new_n217_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT82), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n224_), .A2(new_n233_), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n226_), .A2(new_n230_), .A3(new_n232_), .A4(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n212_), .B1(new_n221_), .B2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n230_), .A2(new_n224_), .A3(new_n232_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(new_n221_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n210_), .A2(new_n211_), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT20), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n204_), .B1(new_n236_), .B2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n218_), .A2(new_n220_), .A3(KEYINPUT96), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(KEYINPUT96), .B1(new_n218_), .B2(new_n220_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n237_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(new_n239_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n212_), .A2(new_n235_), .A3(new_n221_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n204_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n246_), .A2(new_n247_), .A3(KEYINPUT20), .A4(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n241_), .A2(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(G8gat), .B(G36gat), .Z(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G64gat), .B(G92gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT101), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n250_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n248_), .A2(KEYINPUT20), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n235_), .A2(new_n221_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n258_), .B1(new_n259_), .B2(new_n239_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n244_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n225_), .A2(new_n231_), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n261_), .A2(new_n242_), .B1(new_n262_), .B2(new_n230_), .ZN(new_n263_));
  AOI21_X1  g062(.A(KEYINPUT97), .B1(new_n263_), .B2(new_n212_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT97), .ZN(new_n265_));
  NOR3_X1   g064(.A1(new_n245_), .A2(new_n265_), .A3(new_n239_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n260_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n246_), .A2(new_n247_), .A3(KEYINPUT20), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(new_n204_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n255_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n267_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n257_), .A2(new_n271_), .A3(KEYINPUT27), .ZN(new_n272_));
  INV_X1    g071(.A(new_n271_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n270_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n202_), .B(new_n272_), .C1(new_n275_), .C2(KEYINPUT27), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n267_), .A2(new_n269_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n255_), .ZN(new_n278_));
  AOI21_X1  g077(.A(KEYINPUT27), .B1(new_n278_), .B2(new_n271_), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n257_), .A2(KEYINPUT27), .A3(new_n271_), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT102), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n276_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G227gat), .A2(G233gat), .ZN(new_n283_));
  INV_X1    g082(.A(G15gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT30), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n259_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G127gat), .B(G134gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G113gat), .B(G120gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT83), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT83), .B1(new_n288_), .B2(new_n289_), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n287_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G71gat), .B(G99gat), .ZN(new_n297_));
  INV_X1    g096(.A(G43gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT31), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n287_), .A2(new_n295_), .ZN(new_n301_));
  AND3_X1   g100(.A1(new_n296_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n300_), .B1(new_n296_), .B2(new_n301_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n305_));
  XOR2_X1   g104(.A(new_n305_), .B(KEYINPUT88), .Z(new_n306_));
  NOR2_X1   g105(.A1(G141gat), .A2(G148gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT3), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n307_), .A2(KEYINPUT87), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT2), .ZN(new_n310_));
  INV_X1    g109(.A(G141gat), .ZN(new_n311_));
  INV_X1    g110(.A(G148gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n310_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT87), .ZN(new_n314_));
  OAI22_X1  g113(.A1(new_n314_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n315_));
  AND3_X1   g114(.A1(new_n309_), .A2(new_n313_), .A3(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n306_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT85), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT85), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n320_), .A2(G155gat), .A3(G162gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT84), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n317_), .A2(new_n322_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT1), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n319_), .A2(new_n321_), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n324_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n322_), .A2(KEYINPUT1), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT86), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n322_), .A2(KEYINPUT86), .A3(KEYINPUT1), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n328_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n311_), .A2(new_n312_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n334_), .A2(new_n307_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n325_), .B1(new_n333_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n294_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n325_), .B(new_n290_), .C1(new_n333_), .C2(new_n336_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n338_), .A2(KEYINPUT4), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G225gat), .A2(G233gat), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT4), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n337_), .A2(new_n294_), .A3(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n340_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n338_), .A2(new_n341_), .A3(new_n339_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  XOR2_X1   g146(.A(G1gat), .B(G29gat), .Z(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G57gat), .B(G85gat), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n350_), .B(new_n351_), .Z(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n347_), .A2(KEYINPUT100), .A3(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n347_), .A2(new_n353_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT100), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n345_), .A2(new_n352_), .A3(new_n346_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n355_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n304_), .B1(new_n354_), .B2(new_n358_), .ZN(new_n359_));
  XOR2_X1   g158(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n360_));
  AOI21_X1  g159(.A(new_n212_), .B1(new_n337_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(G233gat), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT91), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n364_), .A2(G228gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(G228gat), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n363_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT92), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n337_), .A2(KEYINPUT29), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n212_), .A2(new_n369_), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n362_), .A2(new_n369_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G78gat), .B(G106gat), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT95), .B1(new_n372_), .B2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n372_), .A2(KEYINPUT94), .A3(new_n374_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n370_), .A2(new_n371_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n377_), .B(new_n374_), .C1(new_n361_), .C2(new_n368_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT94), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n377_), .B1(new_n361_), .B2(new_n368_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT95), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n381_), .A2(new_n382_), .A3(new_n373_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n375_), .A2(new_n376_), .A3(new_n380_), .A4(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G22gat), .B(G50gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT90), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n337_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT29), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n387_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  XOR2_X1   g189(.A(KEYINPUT89), .B(KEYINPUT28), .Z(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NOR3_X1   g191(.A1(new_n337_), .A2(KEYINPUT29), .A3(new_n386_), .ZN(new_n393_));
  OR3_X1    g192(.A1(new_n390_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n392_), .B1(new_n390_), .B2(new_n393_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n394_), .A2(new_n395_), .B1(new_n373_), .B2(new_n381_), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n384_), .A2(new_n396_), .B1(new_n397_), .B2(new_n378_), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n282_), .A2(new_n359_), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n384_), .A2(new_n396_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n397_), .A2(new_n378_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n358_), .A2(new_n354_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n279_), .A2(new_n280_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n402_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n250_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n270_), .A2(KEYINPUT32), .ZN(new_n407_));
  MUX2_X1   g206(.A(new_n406_), .B(new_n277_), .S(new_n407_), .Z(new_n408_));
  NAND3_X1  g207(.A1(new_n358_), .A2(new_n354_), .A3(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT33), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n357_), .A2(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n345_), .A2(KEYINPUT33), .A3(new_n352_), .A4(new_n346_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n340_), .A2(new_n341_), .A3(new_n344_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n338_), .A2(new_n342_), .A3(new_n339_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(new_n353_), .A3(new_n414_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n275_), .A2(new_n411_), .A3(new_n412_), .A4(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n409_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n398_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n405_), .A2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n399_), .B1(new_n419_), .B2(new_n304_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G29gat), .B(G36gat), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  XOR2_X1   g221(.A(G43gat), .B(G50gat), .Z(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G43gat), .B(G50gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n421_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT15), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G1gat), .B(G8gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT77), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G15gat), .B(G22gat), .ZN(new_n431_));
  INV_X1    g230(.A(G1gat), .ZN(new_n432_));
  INV_X1    g231(.A(G8gat), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT14), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n431_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n430_), .A2(new_n435_), .ZN(new_n436_));
  OR2_X1    g235(.A1(new_n429_), .A2(KEYINPUT77), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n429_), .A2(KEYINPUT77), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n437_), .A2(new_n434_), .A3(new_n431_), .A4(new_n438_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n436_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n428_), .A2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT80), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G229gat), .A2(G233gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n436_), .A2(new_n439_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n427_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n442_), .A2(new_n443_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(KEYINPUT79), .ZN(new_n447_));
  INV_X1    g246(.A(new_n427_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n440_), .A2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n447_), .B(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n443_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n446_), .A2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G113gat), .B(G141gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G169gat), .B(G197gat), .ZN(new_n455_));
  XOR2_X1   g254(.A(new_n454_), .B(new_n455_), .Z(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n453_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n446_), .A2(new_n452_), .A3(new_n456_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n458_), .A2(KEYINPUT81), .A3(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(KEYINPUT81), .B1(new_n458_), .B2(new_n459_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n420_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT37), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G232gat), .A2(G233gat), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n466_), .B(KEYINPUT34), .Z(new_n467_));
  INV_X1    g266(.A(KEYINPUT35), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n468_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT72), .ZN(new_n471_));
  XOR2_X1   g270(.A(G85gat), .B(G92gat), .Z(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT9), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G85gat), .A2(G92gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT10), .B(G99gat), .ZN(new_n475_));
  OAI221_X1 g274(.A(new_n473_), .B1(KEYINPUT9), .B2(new_n474_), .C1(G106gat), .C2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G99gat), .A2(G106gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT64), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT64), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(G99gat), .A3(G106gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT6), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n478_), .A2(new_n480_), .A3(KEYINPUT6), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n476_), .A2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NOR3_X1   g287(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n483_), .A2(new_n484_), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT8), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(new_n492_), .A3(new_n472_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n481_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT65), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n496_), .A2(KEYINPUT6), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n482_), .A2(KEYINPUT65), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n478_), .B(new_n480_), .C1(new_n497_), .C2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n495_), .A2(new_n499_), .A3(new_n490_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n492_), .B1(new_n500_), .B2(new_n472_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT66), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n493_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  AOI211_X1 g302(.A(KEYINPUT66), .B(new_n492_), .C1(new_n500_), .C2(new_n472_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n486_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n471_), .B1(new_n505_), .B2(new_n448_), .ZN(new_n506_));
  AOI211_X1 g305(.A(new_n469_), .B(new_n506_), .C1(new_n428_), .C2(new_n505_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT73), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT71), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n505_), .A2(new_n509_), .A3(new_n428_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n509_), .B1(new_n505_), .B2(new_n428_), .ZN(new_n512_));
  NOR3_X1   g311(.A1(new_n511_), .A2(new_n506_), .A3(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n469_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n508_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n505_), .A2(new_n428_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT71), .ZN(new_n517_));
  OR2_X1    g316(.A1(new_n505_), .A2(new_n448_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n517_), .A2(new_n518_), .A3(new_n510_), .A4(new_n471_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n519_), .A2(KEYINPUT73), .A3(new_n469_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n507_), .B1(new_n515_), .B2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G190gat), .B(G218gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT74), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G134gat), .B(G162gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT36), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n521_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT36), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n525_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT75), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT76), .ZN(new_n532_));
  AOI211_X1 g331(.A(new_n507_), .B(new_n532_), .C1(new_n515_), .C2(new_n520_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n465_), .B1(new_n528_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n507_), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n531_), .B(KEYINPUT76), .Z(new_n536_));
  NOR3_X1   g335(.A1(new_n513_), .A2(new_n508_), .A3(new_n514_), .ZN(new_n537_));
  AOI21_X1  g336(.A(KEYINPUT73), .B1(new_n519_), .B2(new_n469_), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n535_), .B(new_n536_), .C1(new_n537_), .C2(new_n538_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n539_), .B(KEYINPUT37), .C1(new_n521_), .C2(new_n527_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n534_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G57gat), .B(G64gat), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n542_), .A2(KEYINPUT11), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(KEYINPUT11), .ZN(new_n544_));
  XOR2_X1   g343(.A(G71gat), .B(G78gat), .Z(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n544_), .A2(new_n545_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n505_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT12), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT68), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n549_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n548_), .A2(KEYINPUT68), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n556_), .A2(new_n551_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(new_n505_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n486_), .B(new_n548_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT69), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G230gat), .A2(G233gat), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n559_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n560_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n552_), .B(new_n558_), .C1(new_n562_), .C2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n550_), .A2(KEYINPUT67), .A3(new_n559_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n561_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT67), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n505_), .A2(new_n567_), .A3(new_n549_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n565_), .A2(new_n566_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n564_), .A2(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(G120gat), .B(G148gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G176gat), .B(G204gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n570_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n564_), .A2(new_n569_), .A3(new_n575_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n579_), .A2(KEYINPUT13), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(KEYINPUT13), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(G127gat), .B(G155gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT16), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G183gat), .B(G211gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT17), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  AND2_X1   g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n444_), .B(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n588_), .B1(new_n591_), .B2(new_n548_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n592_), .B1(new_n548_), .B2(new_n591_), .ZN(new_n593_));
  AOI211_X1 g392(.A(new_n587_), .B(new_n586_), .C1(new_n590_), .C2(new_n556_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n594_), .B1(new_n556_), .B2(new_n590_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT78), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n541_), .A2(new_n582_), .A3(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n464_), .A2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT103), .ZN(new_n601_));
  INV_X1    g400(.A(new_n403_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(new_n432_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT38), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n528_), .A2(new_n533_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n420_), .A2(new_n606_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n582_), .A2(new_n463_), .A3(new_n596_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n609_), .B(KEYINPUT104), .Z(new_n610_));
  AOI21_X1  g409(.A(new_n432_), .B1(new_n610_), .B2(new_n602_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n605_), .A2(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n612_), .B1(new_n604_), .B2(new_n603_), .ZN(G1324gat));
  OAI21_X1  g412(.A(G8gat), .B1(new_n609_), .B2(new_n282_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT39), .ZN(new_n615_));
  INV_X1    g414(.A(new_n282_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n601_), .A2(new_n433_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g418(.A(new_n304_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n284_), .B1(new_n610_), .B2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT41), .ZN(new_n622_));
  INV_X1    g421(.A(new_n600_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n623_), .A2(new_n284_), .A3(new_n620_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(G1326gat));
  INV_X1    g424(.A(G22gat), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n626_), .B1(new_n610_), .B2(new_n402_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT42), .Z(new_n628_));
  NAND3_X1  g427(.A1(new_n623_), .A2(new_n626_), .A3(new_n402_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1327gat));
  NAND2_X1  g429(.A1(new_n606_), .A2(new_n598_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n631_), .A2(new_n582_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n464_), .A2(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(G29gat), .B1(new_n633_), .B2(new_n602_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n540_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n535_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(new_n526_), .ZN(new_n637_));
  AOI21_X1  g436(.A(KEYINPUT37), .B1(new_n637_), .B2(new_n539_), .ZN(new_n638_));
  OAI21_X1  g437(.A(KEYINPUT105), .B1(new_n635_), .B2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n635_), .A2(new_n638_), .ZN(new_n640_));
  OAI211_X1 g439(.A(KEYINPUT43), .B(new_n639_), .C1(new_n420_), .C2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n282_), .A2(new_n359_), .A3(new_n398_), .ZN(new_n642_));
  AOI22_X1  g441(.A1(new_n400_), .A2(new_n401_), .B1(new_n354_), .B2(new_n358_), .ZN(new_n643_));
  AOI22_X1  g442(.A1(new_n643_), .A2(new_n404_), .B1(new_n417_), .B2(new_n398_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n642_), .B1(new_n644_), .B2(new_n620_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT43), .ZN(new_n646_));
  OAI211_X1 g445(.A(new_n645_), .B(new_n541_), .C1(KEYINPUT105), .C2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n641_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n582_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n649_), .A2(new_n462_), .A3(new_n598_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(KEYINPUT44), .B1(new_n648_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT44), .ZN(new_n653_));
  AOI211_X1 g452(.A(new_n653_), .B(new_n650_), .C1(new_n641_), .C2(new_n647_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n602_), .A2(G29gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n634_), .B1(new_n655_), .B2(new_n656_), .ZN(G1328gat));
  INV_X1    g456(.A(KEYINPUT46), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n658_), .A2(KEYINPUT108), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT106), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n652_), .A2(new_n654_), .A3(new_n282_), .ZN(new_n662_));
  INV_X1    g461(.A(G36gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n661_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n648_), .A2(new_n651_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(new_n653_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n648_), .A2(KEYINPUT44), .A3(new_n651_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n666_), .A2(new_n616_), .A3(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n668_), .A2(KEYINPUT106), .A3(G36gat), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n664_), .A2(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n633_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n616_), .A2(new_n663_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n672_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n633_), .A2(new_n663_), .A3(new_n616_), .A4(new_n671_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n658_), .A2(KEYINPUT108), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n660_), .B1(new_n670_), .B2(new_n680_), .ZN(new_n681_));
  AOI211_X1 g480(.A(new_n659_), .B(new_n679_), .C1(new_n664_), .C2(new_n669_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1329gat));
  AOI21_X1  g482(.A(G43gat), .B1(new_n633_), .B2(new_n620_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n304_), .A2(new_n298_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n655_), .B2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(G1330gat));
  NAND2_X1  g487(.A1(new_n655_), .A2(new_n402_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n398_), .A2(G50gat), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT110), .Z(new_n691_));
  AOI22_X1  g490(.A1(new_n689_), .A2(G50gat), .B1(new_n633_), .B2(new_n691_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT111), .Z(G1331gat));
  NOR3_X1   g492(.A1(new_n420_), .A2(new_n649_), .A3(new_n462_), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n694_), .A2(new_n640_), .A3(new_n597_), .ZN(new_n695_));
  INV_X1    g494(.A(G57gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n695_), .A2(new_n696_), .A3(new_n602_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n607_), .A2(new_n463_), .A3(new_n582_), .A4(new_n597_), .ZN(new_n698_));
  OAI21_X1  g497(.A(G57gat), .B1(new_n698_), .B2(new_n403_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(G1332gat));
  OAI21_X1  g499(.A(G64gat), .B1(new_n698_), .B2(new_n282_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT48), .ZN(new_n702_));
  INV_X1    g501(.A(G64gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n695_), .A2(new_n703_), .A3(new_n616_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(G1333gat));
  OAI21_X1  g504(.A(G71gat), .B1(new_n698_), .B2(new_n304_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT49), .ZN(new_n707_));
  INV_X1    g506(.A(G71gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n695_), .A2(new_n708_), .A3(new_n620_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(G1334gat));
  OAI21_X1  g509(.A(G78gat), .B1(new_n698_), .B2(new_n398_), .ZN(new_n711_));
  XOR2_X1   g510(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n712_));
  XNOR2_X1  g511(.A(new_n711_), .B(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(G78gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n695_), .A2(new_n714_), .A3(new_n402_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1335gat));
  INV_X1    g515(.A(new_n631_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n694_), .A2(new_n717_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n718_), .A2(G85gat), .A3(new_n403_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n582_), .A2(new_n463_), .A3(new_n598_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n720_), .B1(new_n641_), .B2(new_n647_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(new_n602_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n719_), .B1(G85gat), .B2(new_n722_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT113), .Z(G1336gat));
  AND2_X1   g523(.A1(new_n721_), .A2(new_n616_), .ZN(new_n725_));
  INV_X1    g524(.A(G92gat), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n616_), .A2(new_n726_), .ZN(new_n727_));
  OAI22_X1  g526(.A1(new_n725_), .A2(new_n726_), .B1(new_n718_), .B2(new_n727_), .ZN(G1337gat));
  OR3_X1    g527(.A1(new_n718_), .A2(new_n304_), .A3(new_n475_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n721_), .A2(new_n620_), .ZN(new_n730_));
  INV_X1    g529(.A(G99gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n729_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n732_), .B(new_n733_), .Z(G1338gat));
  NAND2_X1  g533(.A1(new_n721_), .A2(new_n402_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(G106gat), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT116), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT116), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n735_), .A2(new_n738_), .A3(G106gat), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT52), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n737_), .A2(KEYINPUT52), .A3(new_n739_), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n718_), .A2(G106gat), .A3(new_n398_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT115), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n742_), .A2(new_n743_), .A3(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT53), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT53), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n742_), .A2(new_n748_), .A3(new_n743_), .A4(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1339gat));
  NAND3_X1  g549(.A1(new_n442_), .A2(new_n451_), .A3(new_n445_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n450_), .A2(new_n443_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(new_n752_), .A3(new_n457_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n459_), .A2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n579_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT120), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n579_), .A2(KEYINPUT120), .A3(new_n754_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT55), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n552_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n761_));
  AOI22_X1  g560(.A1(new_n564_), .A2(new_n760_), .B1(new_n761_), .B2(new_n566_), .ZN(new_n762_));
  AOI22_X1  g561(.A1(new_n550_), .A2(new_n551_), .B1(new_n557_), .B2(new_n505_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n763_), .B(KEYINPUT55), .C1(new_n563_), .C2(new_n562_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n575_), .B1(new_n762_), .B2(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(KEYINPUT118), .B1(new_n765_), .B2(KEYINPUT56), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n562_), .A2(new_n563_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n552_), .A2(new_n558_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n760_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n761_), .A2(new_n566_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n764_), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n576_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT118), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT56), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n772_), .A2(new_n773_), .A3(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n771_), .A2(KEYINPUT56), .A3(new_n576_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT119), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT119), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n765_), .A2(new_n778_), .A3(KEYINPUT56), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n766_), .A2(new_n775_), .A3(new_n777_), .A4(new_n779_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n462_), .A2(new_n578_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n759_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n606_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT57), .ZN(new_n784_));
  OR2_X1    g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT57), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n786_), .B1(new_n782_), .B2(new_n606_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n754_), .A2(new_n578_), .ZN(new_n788_));
  AOI211_X1 g587(.A(new_n774_), .B(new_n575_), .C1(new_n762_), .C2(new_n764_), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT56), .B1(new_n771_), .B2(new_n576_), .ZN(new_n790_));
  OAI211_X1 g589(.A(KEYINPUT58), .B(new_n788_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n791_), .A2(KEYINPUT121), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(KEYINPUT121), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n788_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT58), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n793_), .A2(new_n541_), .A3(new_n794_), .A4(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n785_), .A2(new_n787_), .A3(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n599_), .A2(new_n463_), .ZN(new_n800_));
  XOR2_X1   g599(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n599_), .B(new_n463_), .C1(KEYINPUT117), .C2(new_n803_), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n799_), .A2(new_n598_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n282_), .A2(new_n602_), .A3(new_n398_), .A4(new_n620_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(KEYINPUT123), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  OR2_X1    g607(.A1(new_n808_), .A2(KEYINPUT126), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT59), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(KEYINPUT126), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n809_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n805_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT125), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT122), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n780_), .A2(new_n781_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n759_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT57), .B1(new_n818_), .B2(new_n783_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n794_), .A2(new_n541_), .A3(new_n797_), .ZN(new_n820_));
  OAI22_X1  g619(.A1(new_n820_), .A2(new_n792_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n815_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n785_), .A2(new_n787_), .A3(new_n798_), .A4(KEYINPUT122), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n822_), .A2(new_n596_), .A3(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n802_), .A2(new_n804_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n808_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n814_), .B1(new_n826_), .B2(new_n810_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n802_), .A2(new_n804_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n596_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n829_), .B1(new_n799_), .B2(new_n815_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n828_), .B1(new_n830_), .B2(new_n823_), .ZN(new_n831_));
  OAI211_X1 g630(.A(KEYINPUT125), .B(KEYINPUT59), .C1(new_n831_), .C2(new_n808_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n813_), .B1(new_n827_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(G113gat), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n463_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT124), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n836_), .B1(new_n831_), .B2(new_n808_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n824_), .A2(new_n825_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n838_), .A2(KEYINPUT124), .A3(new_n807_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n837_), .A2(new_n462_), .A3(new_n839_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n833_), .A2(new_n835_), .B1(new_n834_), .B2(new_n840_), .ZN(G1340gat));
  INV_X1    g640(.A(KEYINPUT60), .ZN(new_n842_));
  AOI21_X1  g641(.A(G120gat), .B1(new_n582_), .B2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n843_), .B1(new_n842_), .B2(G120gat), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n837_), .A2(new_n839_), .A3(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n582_), .B1(new_n805_), .B2(new_n812_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n846_), .B1(new_n827_), .B2(new_n832_), .ZN(new_n847_));
  INV_X1    g646(.A(G120gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n845_), .B1(new_n847_), .B2(new_n848_), .ZN(G1341gat));
  INV_X1    g648(.A(G127gat), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n596_), .A2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n837_), .A2(new_n597_), .A3(new_n839_), .ZN(new_n852_));
  AOI22_X1  g651(.A1(new_n833_), .A2(new_n851_), .B1(new_n850_), .B2(new_n852_), .ZN(G1342gat));
  INV_X1    g652(.A(G134gat), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n640_), .A2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n837_), .A2(new_n606_), .A3(new_n839_), .ZN(new_n856_));
  AOI22_X1  g655(.A1(new_n833_), .A2(new_n855_), .B1(new_n854_), .B2(new_n856_), .ZN(G1343gat));
  NOR3_X1   g656(.A1(new_n616_), .A2(new_n403_), .A3(new_n398_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n838_), .A2(new_n462_), .A3(new_n304_), .A4(new_n858_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(G141gat), .ZN(G1344gat));
  NAND4_X1  g659(.A1(new_n838_), .A2(new_n304_), .A3(new_n582_), .A4(new_n858_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g661(.A1(new_n838_), .A2(new_n304_), .A3(new_n597_), .A4(new_n858_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(KEYINPUT61), .B(G155gat), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n863_), .B(new_n864_), .ZN(G1346gat));
  NAND2_X1  g664(.A1(new_n838_), .A2(new_n304_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n858_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(G162gat), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n868_), .A2(new_n869_), .A3(new_n606_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n866_), .A2(new_n640_), .A3(new_n867_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n869_), .B2(new_n871_), .ZN(G1347gat));
  NAND2_X1  g671(.A1(new_n616_), .A2(new_n359_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n398_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n805_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT22), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n876_), .A2(new_n877_), .A3(new_n462_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n878_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n805_), .A2(new_n875_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n880_), .A2(KEYINPUT62), .A3(new_n463_), .ZN(new_n881_));
  INV_X1    g680(.A(G169gat), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n878_), .A2(KEYINPUT62), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n879_), .B1(new_n883_), .B2(new_n884_), .ZN(G1348gat));
  AOI21_X1  g684(.A(G176gat), .B1(new_n876_), .B2(new_n582_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n831_), .A2(new_n402_), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n582_), .A2(G176gat), .A3(new_n874_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n886_), .B1(new_n887_), .B2(new_n888_), .ZN(G1349gat));
  NOR3_X1   g688(.A1(new_n880_), .A2(new_n222_), .A3(new_n596_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n887_), .A2(new_n597_), .A3(new_n874_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n214_), .ZN(G1350gat));
  OAI21_X1  g691(.A(G190gat), .B1(new_n880_), .B2(new_n640_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n876_), .A2(new_n223_), .A3(new_n606_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1351gat));
  NAND2_X1  g694(.A1(new_n616_), .A2(new_n643_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n831_), .A2(new_n620_), .A3(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT127), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n897_), .A2(new_n898_), .A3(G197gat), .A4(new_n462_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n896_), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n838_), .A2(new_n462_), .A3(new_n304_), .A4(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(G197gat), .ZN(new_n902_));
  OAI21_X1  g701(.A(KEYINPUT127), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n902_), .ZN(new_n904_));
  AND3_X1   g703(.A1(new_n899_), .A2(new_n903_), .A3(new_n904_), .ZN(G1352gat));
  NAND3_X1  g704(.A1(new_n838_), .A2(new_n304_), .A3(new_n900_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n906_), .A2(new_n649_), .ZN(new_n907_));
  INV_X1    g706(.A(G204gat), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n907_), .B(new_n908_), .ZN(G1353gat));
  OR2_X1    g708(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n910_), .B1(new_n897_), .B2(new_n829_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n906_), .A2(new_n596_), .ZN(new_n912_));
  XOR2_X1   g711(.A(KEYINPUT63), .B(G211gat), .Z(new_n913_));
  AOI21_X1  g712(.A(new_n911_), .B1(new_n912_), .B2(new_n913_), .ZN(G1354gat));
  OAI21_X1  g713(.A(G218gat), .B1(new_n906_), .B2(new_n640_), .ZN(new_n915_));
  OR2_X1    g714(.A1(new_n783_), .A2(G218gat), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n906_), .B2(new_n916_), .ZN(G1355gat));
endmodule


