//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 0 0 1 1 0 0 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n782_, new_n783_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n798_, new_n799_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n814_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n824_, new_n825_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G36gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT68), .B(G29gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT15), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT6), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n210_));
  OR3_X1    g009(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  XOR2_X1   g011(.A(G85gat), .B(G92gat), .Z(new_n213_));
  AND2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n214_), .A2(KEYINPUT8), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(KEYINPUT9), .ZN(new_n216_));
  XOR2_X1   g015(.A(KEYINPUT10), .B(G99gat), .Z(new_n217_));
  INV_X1    g016(.A(G106gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(G85gat), .ZN(new_n220_));
  INV_X1    g019(.A(G92gat), .ZN(new_n221_));
  OR3_X1    g020(.A1(new_n220_), .A2(new_n221_), .A3(KEYINPUT9), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n216_), .A2(new_n219_), .A3(new_n222_), .A4(new_n209_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n214_), .A2(KEYINPUT8), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n215_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n207_), .A2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n205_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G232gat), .A2(G233gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT34), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n226_), .B(new_n228_), .C1(KEYINPUT35), .C2(new_n230_), .ZN(new_n231_));
  OAI211_X1 g030(.A(KEYINPUT35), .B(new_n230_), .C1(new_n227_), .C2(KEYINPUT69), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G134gat), .B(G162gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(G190gat), .B(G218gat), .Z(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(new_n238_), .B(KEYINPUT36), .Z(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n233_), .A2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n238_), .A2(KEYINPUT36), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n233_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT72), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT72), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n233_), .A2(new_n245_), .A3(new_n242_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n241_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n247_), .A2(KEYINPUT37), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT37), .ZN(new_n249_));
  AOI211_X1 g048(.A(new_n249_), .B(new_n241_), .C1(new_n244_), .C2(new_n246_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n252_));
  XOR2_X1   g051(.A(G57gat), .B(G64gat), .Z(new_n253_));
  INV_X1    g052(.A(KEYINPUT11), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G71gat), .A2(G78gat), .ZN(new_n256_));
  INV_X1    g055(.A(G71gat), .ZN(new_n257_));
  INV_X1    g056(.A(G78gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n255_), .A2(new_n256_), .A3(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT64), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n261_), .B1(new_n254_), .B2(new_n253_), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n260_), .A2(KEYINPUT64), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n253_), .A2(new_n254_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n260_), .A2(KEYINPUT64), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n263_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n225_), .B1(new_n262_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(G230gat), .ZN(new_n268_));
  INV_X1    g067(.A(G233gat), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n252_), .B1(new_n267_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n270_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n261_), .B(new_n264_), .ZN(new_n273_));
  OAI211_X1 g072(.A(KEYINPUT66), .B(new_n272_), .C1(new_n273_), .C2(new_n225_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT65), .B(KEYINPUT12), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n273_), .A2(new_n225_), .A3(new_n276_), .ZN(new_n277_));
  AOI22_X1  g076(.A1(new_n273_), .A2(new_n225_), .B1(KEYINPUT65), .B2(KEYINPUT12), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n275_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n273_), .A2(new_n225_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n270_), .B1(new_n282_), .B2(new_n267_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G120gat), .B(G148gat), .ZN(new_n285_));
  INV_X1    g084(.A(G204gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G176gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n284_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n284_), .A2(new_n289_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(KEYINPUT67), .A2(KEYINPUT13), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(KEYINPUT67), .A2(KEYINPUT13), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n293_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n291_), .A2(new_n292_), .A3(new_n294_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G231gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n273_), .B(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G15gat), .B(G22gat), .ZN(new_n302_));
  INV_X1    g101(.A(G1gat), .ZN(new_n303_));
  INV_X1    g102(.A(G8gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT14), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G1gat), .B(G8gat), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n306_), .B(new_n307_), .Z(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT73), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n301_), .B(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT17), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n311_), .A2(KEYINPUT74), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  XOR2_X1   g112(.A(KEYINPUT75), .B(KEYINPUT16), .Z(new_n314_));
  XOR2_X1   g113(.A(new_n314_), .B(KEYINPUT76), .Z(new_n315_));
  XOR2_X1   g114(.A(G183gat), .B(G211gat), .Z(new_n316_));
  XNOR2_X1  g115(.A(G127gat), .B(G155gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n315_), .B(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n310_), .B1(new_n313_), .B2(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n313_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n322_), .B1(new_n311_), .B2(new_n320_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n321_), .B1(new_n310_), .B2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n251_), .A2(new_n299_), .A3(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT77), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT78), .ZN(new_n327_));
  INV_X1    g126(.A(new_n308_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n205_), .A2(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n329_), .B1(new_n207_), .B2(new_n328_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G229gat), .A2(G233gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n205_), .B(new_n328_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n331_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n327_), .B1(new_n332_), .B2(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(KEYINPUT78), .B1(new_n333_), .B2(new_n334_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G113gat), .B(G141gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G169gat), .B(G197gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(KEYINPUT79), .B1(new_n338_), .B2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n343_), .B1(new_n338_), .B2(new_n342_), .ZN(new_n344_));
  OR2_X1    g143(.A1(new_n336_), .A2(new_n337_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n345_), .A2(KEYINPUT79), .A3(new_n341_), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT99), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G8gat), .B(G36gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(G92gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT18), .B(G64gat), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n351_), .B(new_n352_), .Z(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G226gat), .A2(G233gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT19), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT21), .ZN(new_n358_));
  INV_X1    g157(.A(G197gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(G204gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n286_), .A2(G197gat), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n358_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  XOR2_X1   g161(.A(G211gat), .B(G218gat), .Z(new_n363_));
  NOR2_X1   g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n286_), .A2(G197gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT88), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT89), .B(KEYINPUT21), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT88), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n368_), .B1(G197gat), .B2(new_n286_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n366_), .B(new_n367_), .C1(new_n365_), .C2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n364_), .A2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n366_), .B1(new_n369_), .B2(new_n365_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n372_), .A2(KEYINPUT21), .A3(new_n363_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  NOR3_X1   g173(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G183gat), .A2(G190gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT23), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT23), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n378_), .A2(G183gat), .A3(G190gat), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n375_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G169gat), .A2(G176gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n380_), .A2(new_n384_), .ZN(new_n385_));
  XOR2_X1   g184(.A(KEYINPUT26), .B(G190gat), .Z(new_n386_));
  XOR2_X1   g185(.A(KEYINPUT25), .B(G183gat), .Z(new_n387_));
  NOR2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT22), .B(G169gat), .ZN(new_n389_));
  INV_X1    g188(.A(G176gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT81), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n383_), .B(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(G183gat), .A2(G190gat), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n395_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n396_));
  OAI22_X1  g195(.A1(new_n385_), .A2(new_n388_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT20), .B1(new_n374_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT97), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n393_), .A2(new_n382_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT80), .B(G183gat), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n401_), .B1(new_n402_), .B2(KEYINPUT25), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n400_), .B(new_n380_), .C1(new_n403_), .C2(new_n386_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n377_), .A2(new_n379_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n405_), .B1(new_n402_), .B2(G190gat), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n406_), .A2(new_n391_), .A3(new_n393_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n404_), .A2(new_n407_), .ZN(new_n408_));
  AOI22_X1  g207(.A1(new_n398_), .A2(new_n399_), .B1(new_n374_), .B2(new_n408_), .ZN(new_n409_));
  OAI211_X1 g208(.A(KEYINPUT97), .B(KEYINPUT20), .C1(new_n374_), .C2(new_n397_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n357_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT20), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n412_), .B1(new_n374_), .B2(new_n397_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n404_), .A2(new_n371_), .A3(new_n373_), .A4(new_n407_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n415_), .A2(new_n356_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n349_), .B(new_n354_), .C1(new_n411_), .C2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n408_), .A2(new_n374_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(new_n357_), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n419_), .A2(new_n398_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT93), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n421_), .B1(new_n415_), .B2(new_n356_), .ZN(new_n422_));
  AOI211_X1 g221(.A(KEYINPUT93), .B(new_n357_), .C1(new_n413_), .C2(new_n414_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n420_), .B(new_n353_), .C1(new_n422_), .C2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n417_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n416_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n398_), .A2(new_n399_), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n427_), .A2(new_n418_), .A3(new_n410_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n426_), .B1(new_n428_), .B2(new_n357_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n349_), .B1(new_n429_), .B2(new_n354_), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT27), .B1(new_n425_), .B2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n420_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n354_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT27), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(new_n434_), .A3(new_n424_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n431_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(G228gat), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n437_), .A2(new_n269_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n374_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT29), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G141gat), .A2(G148gat), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(G141gat), .A2(G148gat), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT85), .ZN(new_n445_));
  AND2_X1   g244(.A1(G155gat), .A2(G162gat), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT1), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n445_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G155gat), .A2(G162gat), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(KEYINPUT85), .A3(KEYINPUT1), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n446_), .A2(new_n447_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NOR3_X1   g253(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n452_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n444_), .B1(new_n451_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT84), .ZN(new_n458_));
  INV_X1    g257(.A(G155gat), .ZN(new_n459_));
  INV_X1    g258(.A(G162gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n446_), .B1(new_n461_), .B2(new_n453_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n443_), .A2(new_n463_), .ZN(new_n464_));
  OAI22_X1  g263(.A1(KEYINPUT86), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT2), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n441_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n469_));
  NAND3_X1  g268(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n468_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n462_), .B1(new_n466_), .B2(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n440_), .B1(new_n457_), .B2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n438_), .B1(new_n439_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT87), .ZN(new_n475_));
  INV_X1    g274(.A(new_n472_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n444_), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n449_), .A2(KEYINPUT85), .A3(KEYINPUT1), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT85), .B1(new_n449_), .B2(KEYINPUT1), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  AOI22_X1  g279(.A1(new_n461_), .A2(new_n453_), .B1(new_n447_), .B2(new_n446_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n477_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n475_), .B1(new_n476_), .B2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n457_), .A2(KEYINPUT87), .A3(new_n472_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n440_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n374_), .B1(new_n437_), .B2(new_n269_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n474_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT91), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G78gat), .B(G106gat), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT91), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n474_), .B(new_n490_), .C1(new_n485_), .C2(new_n486_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n488_), .A2(new_n489_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT92), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n483_), .A2(new_n484_), .ZN(new_n494_));
  OAI21_X1  g293(.A(G50gat), .B1(new_n494_), .B2(KEYINPUT29), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT28), .B(G22gat), .ZN(new_n496_));
  INV_X1    g295(.A(G50gat), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n483_), .A2(new_n440_), .A3(new_n497_), .A4(new_n484_), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n495_), .A2(new_n496_), .A3(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n496_), .B1(new_n495_), .B2(new_n498_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n487_), .A2(new_n489_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT92), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n488_), .A2(new_n503_), .A3(new_n489_), .A4(new_n491_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n493_), .A2(new_n501_), .A3(new_n502_), .A4(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT90), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n487_), .A2(new_n506_), .A3(new_n489_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n506_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n502_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n509_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n505_), .A2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n436_), .A2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G15gat), .B(G43gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G227gat), .A2(G233gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G71gat), .B(G99gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n408_), .B(KEYINPUT30), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT82), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n519_), .A2(KEYINPUT82), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n518_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n522_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n524_), .A2(new_n520_), .A3(new_n517_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(new_n525_), .A3(KEYINPUT83), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G127gat), .B(G134gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G113gat), .B(G120gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT31), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n526_), .B(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n529_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n457_), .A2(KEYINPUT87), .A3(new_n472_), .ZN(new_n534_));
  AOI21_X1  g333(.A(KEYINPUT87), .B1(new_n457_), .B2(new_n472_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n533_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G225gat), .A2(G233gat), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n457_), .A2(new_n529_), .A3(new_n472_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT94), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT94), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n536_), .A2(new_n541_), .A3(new_n537_), .A4(new_n538_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n537_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT4), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n545_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n546_));
  AOI21_X1  g345(.A(KEYINPUT4), .B1(new_n494_), .B2(new_n533_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n544_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G1gat), .B(G29gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(new_n220_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT0), .B(G57gat), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n550_), .B(new_n551_), .Z(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n543_), .A2(new_n548_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n553_), .B1(new_n543_), .B2(new_n548_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n532_), .A2(new_n557_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n512_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n511_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT33), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n554_), .A2(KEYINPUT95), .A3(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n561_), .B1(new_n554_), .B2(KEYINPUT95), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n537_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n536_), .A2(new_n544_), .A3(new_n538_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n564_), .A2(new_n552_), .A3(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n433_), .A2(new_n566_), .A3(new_n424_), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n562_), .A2(new_n563_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n556_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n411_), .A2(new_n416_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n420_), .B(KEYINPUT96), .C1(new_n422_), .C2(new_n423_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n353_), .A2(KEYINPUT32), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n570_), .A2(new_n571_), .A3(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n572_), .B1(new_n432_), .B2(KEYINPUT96), .ZN(new_n575_));
  AOI22_X1  g374(.A1(new_n569_), .A2(new_n554_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n560_), .B1(new_n568_), .B2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT98), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n431_), .A2(new_n435_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n579_), .A2(new_n557_), .A3(new_n511_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n554_), .A2(KEYINPUT95), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT33), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n433_), .A2(new_n424_), .A3(new_n566_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n554_), .A2(KEYINPUT95), .A3(new_n561_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n582_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n574_), .A2(new_n575_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n586_), .B1(new_n556_), .B2(new_n555_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n511_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT98), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n578_), .A2(new_n580_), .A3(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n532_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n559_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n326_), .A2(new_n348_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n557_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n594_), .A2(new_n303_), .A3(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT38), .ZN(new_n597_));
  INV_X1    g396(.A(new_n299_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n598_), .A2(new_n348_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n559_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n588_), .A2(new_n589_), .ZN(new_n601_));
  AOI211_X1 g400(.A(KEYINPUT98), .B(new_n511_), .C1(new_n585_), .C2(new_n587_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n580_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n601_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n600_), .B1(new_n604_), .B2(new_n532_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n247_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n599_), .A2(new_n605_), .A3(new_n606_), .A4(new_n324_), .ZN(new_n607_));
  OAI21_X1  g406(.A(G1gat), .B1(new_n607_), .B2(new_n557_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n597_), .A2(new_n608_), .ZN(G1324gat));
  OAI21_X1  g408(.A(G8gat), .B1(new_n607_), .B2(new_n579_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n610_), .A2(KEYINPUT101), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(KEYINPUT101), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT102), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n611_), .A2(KEYINPUT102), .A3(new_n612_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n615_), .A2(KEYINPUT39), .A3(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n594_), .A2(new_n304_), .A3(new_n436_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT100), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT39), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n613_), .A2(new_n614_), .A3(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n617_), .A2(new_n619_), .A3(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g422(.A(G15gat), .B1(new_n607_), .B2(new_n592_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT41), .Z(new_n625_));
  INV_X1    g424(.A(G15gat), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n594_), .A2(new_n626_), .A3(new_n532_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(G1326gat));
  OAI21_X1  g427(.A(G22gat), .B1(new_n607_), .B2(new_n560_), .ZN(new_n629_));
  XOR2_X1   g428(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(G22gat), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n594_), .A2(new_n632_), .A3(new_n511_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(G1327gat));
  NOR3_X1   g433(.A1(new_n598_), .A2(new_n348_), .A3(new_n324_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n635_), .A2(new_n605_), .A3(new_n247_), .ZN(new_n636_));
  AOI21_X1  g435(.A(G29gat), .B1(new_n636_), .B2(new_n595_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT43), .ZN(new_n638_));
  INV_X1    g437(.A(new_n251_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n605_), .B2(new_n639_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n593_), .A2(KEYINPUT43), .A3(new_n251_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n635_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT44), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  OAI211_X1 g443(.A(KEYINPUT44), .B(new_n635_), .C1(new_n640_), .C2(new_n641_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n595_), .A2(G29gat), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n637_), .B1(new_n647_), .B2(new_n648_), .ZN(G1328gat));
  NAND3_X1  g448(.A1(new_n644_), .A2(new_n436_), .A3(new_n645_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT104), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n644_), .A2(KEYINPUT104), .A3(new_n436_), .A4(new_n645_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(G36gat), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(G36gat), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n636_), .A2(new_n655_), .A3(new_n436_), .ZN(new_n656_));
  XOR2_X1   g455(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n654_), .A2(KEYINPUT106), .A3(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT107), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT46), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT108), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n654_), .A2(new_n658_), .ZN(new_n665_));
  OAI21_X1  g464(.A(KEYINPUT106), .B1(new_n662_), .B2(KEYINPUT107), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n663_), .A2(new_n664_), .A3(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(KEYINPUT46), .B1(new_n659_), .B2(new_n660_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n665_), .A2(new_n666_), .ZN(new_n670_));
  OAI21_X1  g469(.A(KEYINPUT108), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n668_), .A2(new_n671_), .ZN(G1329gat));
  OAI21_X1  g471(.A(G43gat), .B1(new_n646_), .B2(new_n592_), .ZN(new_n673_));
  INV_X1    g472(.A(G43gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n636_), .A2(new_n674_), .A3(new_n532_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g476(.A(G50gat), .B1(new_n646_), .B2(new_n560_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n636_), .A2(new_n497_), .A3(new_n511_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1331gat));
  NAND2_X1  g479(.A1(new_n598_), .A2(new_n348_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n324_), .ZN(new_n682_));
  NOR4_X1   g481(.A1(new_n681_), .A2(new_n639_), .A3(new_n593_), .A4(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(G57gat), .B1(new_n683_), .B2(new_n595_), .ZN(new_n684_));
  NOR4_X1   g483(.A1(new_n681_), .A2(new_n593_), .A3(new_n247_), .A4(new_n682_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n595_), .A2(G57gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n684_), .B1(new_n685_), .B2(new_n686_), .ZN(G1332gat));
  INV_X1    g486(.A(G64gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n685_), .B2(new_n436_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT48), .Z(new_n690_));
  NAND3_X1  g489(.A1(new_n683_), .A2(new_n688_), .A3(new_n436_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1333gat));
  AOI21_X1  g491(.A(new_n257_), .B1(new_n685_), .B2(new_n532_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT49), .Z(new_n694_));
  NAND3_X1  g493(.A1(new_n683_), .A2(new_n257_), .A3(new_n532_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT109), .ZN(G1334gat));
  AOI21_X1  g496(.A(new_n258_), .B1(new_n685_), .B2(new_n511_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n698_), .B(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n683_), .A2(new_n258_), .A3(new_n511_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1335gat));
  NOR4_X1   g501(.A1(new_n681_), .A2(new_n593_), .A3(new_n606_), .A4(new_n324_), .ZN(new_n703_));
  AOI21_X1  g502(.A(G85gat), .B1(new_n703_), .B2(new_n595_), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n640_), .A2(new_n641_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n681_), .A2(new_n324_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n557_), .A2(new_n220_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n704_), .B1(new_n707_), .B2(new_n708_), .ZN(G1336gat));
  AOI21_X1  g508(.A(G92gat), .B1(new_n703_), .B2(new_n436_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n579_), .A2(new_n221_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n707_), .B2(new_n711_), .ZN(G1337gat));
  INV_X1    g511(.A(new_n707_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G99gat), .B1(new_n713_), .B2(new_n592_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n703_), .A2(new_n217_), .A3(new_n532_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT111), .Z(new_n716_));
  NAND3_X1  g515(.A1(new_n714_), .A2(KEYINPUT112), .A3(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT51), .ZN(G1338gat));
  AOI21_X1  g517(.A(new_n218_), .B1(new_n707_), .B2(new_n511_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT52), .Z(new_n720_));
  NAND3_X1  g519(.A1(new_n703_), .A2(new_n218_), .A3(new_n511_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT113), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g523(.A1(new_n251_), .A2(new_n348_), .A3(new_n299_), .A4(new_n324_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT54), .Z(new_n726_));
  INV_X1    g525(.A(KEYINPUT55), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n280_), .A2(new_n727_), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n277_), .A2(new_n278_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n270_), .B1(new_n729_), .B2(new_n267_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n275_), .A2(new_n279_), .A3(KEYINPUT55), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n728_), .A2(new_n730_), .A3(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n289_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT56), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT114), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n732_), .A2(KEYINPUT56), .A3(new_n289_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n735_), .A2(new_n736_), .A3(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT56), .B1(new_n732_), .B2(new_n289_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n290_), .B1(new_n739_), .B2(KEYINPUT114), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n738_), .A2(new_n347_), .A3(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT115), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n333_), .A2(new_n331_), .ZN(new_n743_));
  AOI211_X1 g542(.A(new_n342_), .B(new_n743_), .C1(new_n334_), .C2(new_n330_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(new_n338_), .B2(new_n342_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n293_), .A2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT115), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n738_), .A2(new_n740_), .A3(new_n347_), .A4(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n742_), .A2(new_n746_), .A3(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(new_n606_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n735_), .A2(new_n737_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n753_), .A2(new_n291_), .A3(new_n745_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT58), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n755_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(new_n757_), .A3(new_n639_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n751_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n749_), .A2(new_n606_), .A3(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n752_), .A2(new_n758_), .A3(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n726_), .B1(new_n761_), .B2(new_n682_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n512_), .A2(new_n595_), .A3(new_n532_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT117), .Z(new_n764_));
  NOR2_X1   g563(.A1(new_n762_), .A2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(G113gat), .B1(new_n765_), .B2(new_n347_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT59), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT118), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n762_), .B2(new_n768_), .ZN(new_n769_));
  OR2_X1    g568(.A1(new_n769_), .A2(new_n765_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n765_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n348_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n766_), .B1(new_n772_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g572(.A(G120gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n774_), .B1(new_n299_), .B2(KEYINPUT60), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n765_), .B(new_n775_), .C1(KEYINPUT60), .C2(new_n774_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n299_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n777_), .B2(new_n774_), .ZN(G1341gat));
  AOI21_X1  g577(.A(G127gat), .B1(new_n765_), .B2(new_n324_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n682_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n780_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g580(.A(G134gat), .B1(new_n765_), .B2(new_n247_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n251_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n783_), .B2(G134gat), .ZN(G1343gat));
  NOR2_X1   g583(.A1(new_n532_), .A2(new_n560_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n785_), .A2(new_n595_), .A3(new_n579_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT119), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n762_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n347_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(KEYINPUT120), .B(G141gat), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n789_), .B(new_n790_), .ZN(G1344gat));
  NAND2_X1  g590(.A1(new_n788_), .A2(new_n598_), .ZN(new_n792_));
  XOR2_X1   g591(.A(KEYINPUT121), .B(G148gat), .Z(new_n793_));
  XNOR2_X1  g592(.A(new_n792_), .B(new_n793_), .ZN(G1345gat));
  NAND2_X1  g593(.A1(new_n788_), .A2(new_n324_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(KEYINPUT61), .B(G155gat), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n795_), .B(new_n796_), .ZN(G1346gat));
  AOI21_X1  g596(.A(G162gat), .B1(new_n788_), .B2(new_n247_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n251_), .A2(new_n460_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n788_), .B2(new_n799_), .ZN(G1347gat));
  INV_X1    g599(.A(G169gat), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n762_), .A2(new_n511_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n579_), .A2(new_n595_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n532_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT122), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n802_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n801_), .B1(new_n806_), .B2(new_n347_), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n807_), .A2(KEYINPUT62), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n802_), .A2(new_n805_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n389_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n809_), .A2(new_n348_), .A3(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(KEYINPUT62), .B1(new_n807_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n808_), .A2(new_n812_), .ZN(G1348gat));
  NOR2_X1   g612(.A1(new_n809_), .A2(new_n299_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(new_n390_), .ZN(G1349gat));
  OAI21_X1  g614(.A(new_n402_), .B1(new_n809_), .B2(new_n682_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n809_), .A2(new_n387_), .A3(new_n682_), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT123), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT123), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n806_), .A2(new_n324_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n820_), .B(new_n816_), .C1(new_n821_), .C2(new_n387_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n819_), .A2(new_n822_), .ZN(G1350gat));
  OAI21_X1  g622(.A(G190gat), .B1(new_n809_), .B2(new_n251_), .ZN(new_n824_));
  OR2_X1    g623(.A1(new_n809_), .A2(new_n386_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n825_), .B2(new_n606_), .ZN(G1351gat));
  INV_X1    g625(.A(new_n726_), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n749_), .A2(new_n606_), .A3(new_n759_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n759_), .B1(new_n749_), .B2(new_n606_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n758_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n828_), .A2(new_n829_), .A3(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n827_), .B1(new_n831_), .B2(new_n324_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(new_n785_), .A3(new_n803_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT124), .ZN(new_n834_));
  INV_X1    g633(.A(new_n785_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n761_), .A2(new_n682_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(new_n827_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT124), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(new_n838_), .A3(new_n803_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n834_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(G197gat), .B1(new_n841_), .B2(new_n348_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n840_), .A2(new_n359_), .A3(new_n347_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(G1352gat));
  XNOR2_X1  g643(.A(KEYINPUT125), .B(G204gat), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(new_n841_), .B2(new_n299_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n840_), .A2(new_n598_), .A3(new_n845_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1353gat));
  AOI21_X1  g648(.A(new_n838_), .B1(new_n837_), .B2(new_n803_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n803_), .ZN(new_n851_));
  NOR4_X1   g650(.A1(new_n762_), .A2(KEYINPUT124), .A3(new_n835_), .A4(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n324_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(KEYINPUT63), .B(G211gat), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT126), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n682_), .B1(new_n834_), .B2(new_n839_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n856_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n853_), .A2(KEYINPUT126), .A3(new_n858_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n855_), .B1(new_n860_), .B2(new_n861_), .ZN(G1354gat));
  XNOR2_X1  g661(.A(KEYINPUT127), .B(G218gat), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n863_), .B1(new_n840_), .B2(new_n247_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n639_), .A2(new_n863_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n840_), .B2(new_n865_), .ZN(G1355gat));
endmodule


