//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 1 1 0 1 1 0 1 1 1 0 0 1 1 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 1 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n873_, new_n874_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT69), .B(G71gat), .Z(new_n203_));
  INV_X1    g002(.A(G78gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT69), .B(G71gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G78gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT11), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G57gat), .B(G64gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n205_), .A2(KEYINPUT11), .A3(new_n207_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  OR3_X1    g012(.A1(new_n208_), .A2(new_n209_), .A3(new_n211_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT12), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT6), .ZN(new_n218_));
  AND3_X1   g017(.A1(KEYINPUT65), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT65), .B1(G99gat), .B2(G106gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n218_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G99gat), .A2(G106gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(KEYINPUT65), .A2(G99gat), .A3(G106gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(KEYINPUT6), .A3(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n221_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT10), .B(G99gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n228_), .A2(G106gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n227_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G85gat), .B(G92gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT9), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT9), .ZN(new_n233_));
  INV_X1    g032(.A(G85gat), .ZN(new_n234_));
  INV_X1    g033(.A(G92gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n233_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  AND3_X1   g035(.A1(new_n232_), .A2(KEYINPUT64), .A3(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(KEYINPUT64), .B1(new_n232_), .B2(new_n236_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n230_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n224_), .B(new_n225_), .C1(new_n242_), .C2(new_n243_), .ZN(new_n244_));
  OR2_X1    g043(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n245_), .B(new_n241_), .C1(new_n219_), .C2(new_n220_), .ZN(new_n246_));
  OR2_X1    g045(.A1(G99gat), .A2(G106gat), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT7), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n248_), .A2(KEYINPUT66), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n250_), .A2(KEYINPUT7), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n247_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(KEYINPUT7), .ZN(new_n253_));
  NOR2_X1   g052(.A1(G99gat), .A2(G106gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n244_), .A2(new_n246_), .A3(new_n252_), .A4(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n231_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT8), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT8), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n260_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n221_), .A2(new_n226_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n255_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n248_), .A2(KEYINPUT66), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n254_), .B1(new_n253_), .B2(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n261_), .B1(new_n262_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n259_), .A2(new_n268_), .A3(KEYINPUT70), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT70), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n260_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n270_), .B1(new_n271_), .B2(new_n267_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n240_), .B1(new_n269_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  AOI211_X1 g074(.A(KEYINPUT71), .B(new_n240_), .C1(new_n269_), .C2(new_n272_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n217_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  AND2_X1   g076(.A1(new_n213_), .A2(new_n214_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n239_), .B1(new_n271_), .B2(new_n267_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n239_), .B(KEYINPUT68), .C1(new_n271_), .C2(new_n267_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n278_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n281_), .A2(new_n282_), .A3(new_n278_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n283_), .B1(new_n216_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G230gat), .A2(G233gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n277_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n281_), .A2(new_n282_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n215_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(new_n284_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n286_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(G120gat), .B(G148gat), .Z(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XOR2_X1   g094(.A(G176gat), .B(G204gat), .Z(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT72), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n287_), .A2(new_n292_), .A3(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n298_), .B1(new_n287_), .B2(new_n292_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n202_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n301_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n303_), .A2(KEYINPUT13), .A3(new_n299_), .ZN(new_n304_));
  AND3_X1   g103(.A1(new_n302_), .A2(new_n304_), .A3(KEYINPUT74), .ZN(new_n305_));
  AOI21_X1  g104(.A(KEYINPUT74), .B1(new_n302_), .B2(new_n304_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  AND2_X1   g106(.A1(G231gat), .A2(G233gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n278_), .B(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(G15gat), .B(G22gat), .Z(new_n310_));
  XOR2_X1   g109(.A(KEYINPUT80), .B(G1gat), .Z(new_n311_));
  XOR2_X1   g110(.A(KEYINPUT81), .B(G8gat), .Z(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n310_), .B1(new_n313_), .B2(KEYINPUT14), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G1gat), .B(G8gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n314_), .B(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n309_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G127gat), .B(G155gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G183gat), .B(G211gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n323_), .A2(KEYINPUT17), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n215_), .B(new_n308_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n314_), .B(new_n315_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n318_), .A2(new_n324_), .A3(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n323_), .B(KEYINPUT17), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n329_), .B1(new_n318_), .B2(new_n327_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT83), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT37), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G232gat), .A2(G233gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT34), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT35), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G29gat), .B(G36gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT75), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G43gat), .B(G50gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n342_), .A2(KEYINPUT15), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n342_), .A2(KEYINPUT15), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(KEYINPUT70), .B1(new_n259_), .B2(new_n268_), .ZN(new_n346_));
  NOR3_X1   g145(.A1(new_n271_), .A2(new_n267_), .A3(new_n270_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n239_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT71), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n273_), .A2(new_n274_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n345_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  AOI22_X1  g150(.A1(new_n288_), .A2(new_n342_), .B1(new_n337_), .B2(new_n336_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n338_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n354_));
  OAI22_X1  g153(.A1(new_n275_), .A2(new_n276_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n338_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n355_), .A2(new_n356_), .A3(new_n352_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G190gat), .B(G218gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT76), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G134gat), .B(G162gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT36), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(KEYINPUT77), .B(KEYINPUT78), .Z(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n354_), .A2(new_n357_), .A3(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n361_), .B(new_n362_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT79), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n368_), .B1(new_n354_), .B2(new_n357_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n333_), .B1(new_n366_), .B2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n354_), .A2(new_n357_), .A3(new_n365_), .ZN(new_n371_));
  NOR3_X1   g170(.A1(new_n351_), .A2(new_n353_), .A3(new_n338_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n356_), .B1(new_n355_), .B2(new_n352_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  OAI211_X1 g173(.A(KEYINPUT37), .B(new_n371_), .C1(new_n374_), .C2(new_n368_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n332_), .A2(new_n370_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT104), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G127gat), .B(G134gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G113gat), .B(G120gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  OR2_X1    g180(.A1(new_n381_), .A2(KEYINPUT101), .ZN(new_n382_));
  NOR2_X1   g181(.A1(KEYINPUT91), .A2(KEYINPUT3), .ZN(new_n383_));
  INV_X1    g182(.A(G141gat), .ZN(new_n384_));
  INV_X1    g183(.A(G148gat), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n383_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G141gat), .A2(G148gat), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT2), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n390_));
  OAI22_X1  g189(.A1(KEYINPUT91), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n386_), .A2(new_n389_), .A3(new_n390_), .A4(new_n391_), .ZN(new_n392_));
  OR2_X1    g191(.A1(G155gat), .A2(G162gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G155gat), .A2(G162gat), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n392_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  OR2_X1    g194(.A1(new_n394_), .A2(KEYINPUT1), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(KEYINPUT1), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n396_), .A2(new_n393_), .A3(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n384_), .A2(new_n385_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(new_n387_), .A3(new_n399_), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n395_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n381_), .A2(KEYINPUT101), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n382_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n380_), .A2(KEYINPUT89), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n378_), .A2(new_n379_), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n405_), .A2(KEYINPUT89), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  OR2_X1    g206(.A1(new_n407_), .A2(new_n401_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n403_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G225gat), .A2(G233gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G1gat), .B(G29gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(G85gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT0), .B(G57gat), .ZN(new_n414_));
  XOR2_X1   g213(.A(new_n413_), .B(new_n414_), .Z(new_n415_));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n408_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n403_), .A2(new_n408_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n417_), .B1(KEYINPUT4), .B2(new_n418_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n411_), .B(new_n415_), .C1(new_n419_), .C2(new_n410_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT102), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n410_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n409_), .A2(new_n416_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n423_), .B1(new_n424_), .B2(new_n417_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n425_), .A2(KEYINPUT102), .A3(new_n411_), .A4(new_n415_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n411_), .B1(new_n419_), .B2(new_n410_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n415_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n422_), .A2(new_n426_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G228gat), .A2(G233gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(new_n204_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  XOR2_X1   g232(.A(G197gat), .B(G204gat), .Z(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT21), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT93), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G211gat), .B(G218gat), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT94), .ZN(new_n438_));
  OR3_X1    g237(.A1(new_n434_), .A2(new_n438_), .A3(KEYINPUT21), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n438_), .B1(new_n434_), .B2(KEYINPUT21), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n436_), .A2(new_n437_), .A3(new_n439_), .A4(new_n440_), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n437_), .A2(KEYINPUT95), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n437_), .A2(KEYINPUT95), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n442_), .A2(KEYINPUT21), .A3(new_n443_), .A4(new_n434_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n441_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(G106gat), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT29), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n401_), .A2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n445_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n446_), .B1(new_n445_), .B2(new_n448_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n433_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n451_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n453_), .A2(new_n432_), .A3(new_n449_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT92), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n452_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT96), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT96), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n452_), .A2(new_n454_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n401_), .A2(new_n447_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT28), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G22gat), .B(G50gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n457_), .A2(new_n459_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n463_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n456_), .A2(KEYINPUT96), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G183gat), .A2(G190gat), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n469_), .A2(KEYINPUT23), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n468_), .B(KEYINPUT87), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n470_), .B1(new_n471_), .B2(KEYINPUT23), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n472_), .B1(G183gat), .B2(G190gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT22), .B(G169gat), .ZN(new_n474_));
  INV_X1    g273(.A(G176gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G169gat), .A2(G176gat), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n473_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(KEYINPUT24), .ZN(new_n479_));
  NOR2_X1   g278(.A1(G169gat), .A2(G176gat), .ZN(new_n480_));
  MUX2_X1   g279(.A(new_n479_), .B(KEYINPUT24), .S(new_n480_), .Z(new_n481_));
  XNOR2_X1  g280(.A(KEYINPUT26), .B(G190gat), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT86), .ZN(new_n483_));
  INV_X1    g282(.A(G183gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT25), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n484_), .A2(KEYINPUT25), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n482_), .B(new_n485_), .C1(new_n486_), .C2(new_n483_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n481_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT23), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n469_), .A2(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n490_), .B1(new_n471_), .B2(new_n489_), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(G71gat), .B(G99gat), .Z(new_n493_));
  XNOR2_X1  g292(.A(G15gat), .B(G43gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n478_), .A2(new_n492_), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n495_), .B1(new_n478_), .B2(new_n492_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n404_), .B(new_n406_), .C1(new_n497_), .C2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G227gat), .A2(G233gat), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n500_), .B(KEYINPUT88), .Z(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT30), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT31), .ZN(new_n503_));
  INV_X1    g302(.A(new_n498_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n504_), .A2(new_n407_), .A3(new_n496_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n499_), .A2(new_n503_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n503_), .B1(new_n499_), .B2(new_n505_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n467_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT90), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n512_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n508_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(KEYINPUT90), .A3(new_n506_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n464_), .A2(new_n466_), .A3(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n430_), .B1(new_n511_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT99), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n441_), .A2(new_n444_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(G183gat), .A2(G190gat), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT98), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n474_), .B(new_n522_), .ZN(new_n523_));
  OAI221_X1 g322(.A(new_n477_), .B1(new_n491_), .B2(new_n521_), .C1(G176gat), .C2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT25), .B(G183gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n482_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n472_), .A2(new_n481_), .A3(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n519_), .B1(new_n520_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT20), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n478_), .A2(new_n492_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n531_), .B1(new_n520_), .B2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n445_), .A2(KEYINPUT99), .A3(new_n528_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n530_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G226gat), .A2(G233gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT19), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n538_), .B(KEYINPUT97), .Z(new_n539_));
  NAND2_X1  g338(.A1(new_n536_), .A2(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n531_), .B1(new_n520_), .B2(new_n529_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n538_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n445_), .A2(new_n532_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT100), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT100), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n541_), .A2(new_n546_), .A3(new_n542_), .A4(new_n543_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n540_), .A2(new_n545_), .A3(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G8gat), .B(G36gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT18), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G64gat), .B(G92gat), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n550_), .B(new_n551_), .Z(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n548_), .A2(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n540_), .A2(new_n545_), .A3(new_n552_), .A4(new_n547_), .ZN(new_n555_));
  AOI21_X1  g354(.A(KEYINPUT27), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n541_), .A2(new_n543_), .ZN(new_n557_));
  OAI22_X1  g356(.A1(new_n557_), .A2(new_n542_), .B1(new_n536_), .B2(new_n539_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n553_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n559_), .A2(new_n555_), .A3(KEYINPUT103), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n540_), .A2(new_n545_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT103), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n561_), .A2(new_n562_), .A3(new_n552_), .A4(new_n547_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n560_), .A2(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n556_), .B1(new_n564_), .B2(KEYINPUT27), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n552_), .A2(KEYINPUT32), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n558_), .A2(new_n566_), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n430_), .B(new_n567_), .C1(new_n548_), .C2(new_n566_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT33), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n420_), .A2(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n410_), .B1(new_n424_), .B2(new_n417_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n415_), .B1(new_n409_), .B2(new_n423_), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n420_), .A2(new_n569_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n570_), .A2(new_n554_), .A3(new_n573_), .A4(new_n555_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n568_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n516_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n576_), .B1(new_n464_), .B2(new_n466_), .ZN(new_n577_));
  AOI22_X1  g376(.A1(new_n518_), .A2(new_n565_), .B1(new_n575_), .B2(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n317_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G229gat), .A2(G233gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n326_), .A2(new_n342_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n341_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n340_), .B(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n317_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT84), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(new_n581_), .A3(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n317_), .A2(KEYINPUT84), .A3(new_n584_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n580_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n587_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G113gat), .B(G141gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G169gat), .B(G197gat), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n591_), .B(new_n592_), .Z(new_n593_));
  NAND3_X1  g392(.A1(new_n582_), .A2(new_n590_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT85), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n582_), .A2(new_n590_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n593_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n596_), .B(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n377_), .B1(new_n578_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n575_), .A2(new_n577_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n564_), .A2(KEYINPUT27), .ZN(new_n604_));
  INV_X1    g403(.A(new_n556_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n430_), .ZN(new_n607_));
  AND3_X1   g406(.A1(new_n464_), .A2(new_n466_), .A3(new_n516_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n509_), .B1(new_n464_), .B2(new_n466_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n607_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n603_), .B1(new_n606_), .B2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n611_), .A2(KEYINPUT104), .A3(new_n600_), .ZN(new_n612_));
  AOI211_X1 g411(.A(new_n307_), .B(new_n376_), .C1(new_n602_), .C2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n311_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n430_), .B(KEYINPUT105), .Z(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n613_), .A2(new_n614_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT107), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n617_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n618_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n621_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n366_), .A2(new_n369_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n611_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n331_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n307_), .A2(new_n601_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(new_n430_), .ZN(new_n631_));
  AOI22_X1  g430(.A1(new_n617_), .A2(new_n623_), .B1(new_n631_), .B2(G1gat), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n622_), .A2(new_n632_), .ZN(G1324gat));
  NAND3_X1  g432(.A1(new_n628_), .A2(new_n606_), .A3(new_n629_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(G8gat), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT39), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n635_), .A2(KEYINPUT108), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n312_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n613_), .A2(new_n638_), .A3(new_n606_), .ZN(new_n639_));
  XOR2_X1   g438(.A(KEYINPUT108), .B(KEYINPUT39), .Z(new_n640_));
  OAI211_X1 g439(.A(new_n637_), .B(new_n639_), .C1(new_n635_), .C2(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(G1325gat));
  INV_X1    g442(.A(G15gat), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n613_), .A2(new_n644_), .A3(new_n576_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n628_), .A2(new_n576_), .A3(new_n629_), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n646_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT41), .B1(new_n646_), .B2(G15gat), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n645_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT110), .Z(G1326gat));
  INV_X1    g449(.A(G22gat), .ZN(new_n651_));
  INV_X1    g450(.A(new_n467_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n651_), .B1(new_n630_), .B2(new_n652_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT42), .Z(new_n654_));
  NAND3_X1  g453(.A1(new_n613_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1327gat));
  INV_X1    g455(.A(KEYINPUT83), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n331_), .B(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(new_n624_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT112), .ZN(new_n660_));
  INV_X1    g459(.A(new_n307_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n662_), .B1(new_n602_), .B2(new_n612_), .ZN(new_n663_));
  AOI21_X1  g462(.A(G29gat), .B1(new_n663_), .B2(new_n430_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n370_), .A2(new_n375_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n611_), .A2(new_n665_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n370_), .A2(new_n375_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT111), .ZN(new_n668_));
  OAI21_X1  g467(.A(KEYINPUT43), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n666_), .A2(new_n669_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n611_), .A2(new_n668_), .A3(KEYINPUT43), .A4(new_n665_), .ZN(new_n671_));
  AND4_X1   g470(.A1(new_n658_), .A2(new_n670_), .A3(new_n629_), .A4(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT44), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n673_), .A2(G29gat), .A3(new_n616_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n332_), .B1(new_n666_), .B2(new_n669_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n675_), .A2(new_n629_), .A3(new_n671_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n664_), .B1(new_n674_), .B2(new_n678_), .ZN(G1328gat));
  INV_X1    g478(.A(KEYINPUT46), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT45), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT113), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n565_), .A2(G36gat), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n663_), .A2(new_n682_), .A3(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n682_), .B1(new_n663_), .B2(new_n683_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n681_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n663_), .A2(new_n683_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT113), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n663_), .A2(new_n682_), .A3(new_n683_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n688_), .A2(KEYINPUT45), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n686_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(G36gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n565_), .B1(new_n672_), .B2(KEYINPUT44), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n693_), .B2(new_n678_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n680_), .B1(new_n691_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n678_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n606_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n697_));
  OAI21_X1  g496(.A(G36gat), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n698_), .A2(KEYINPUT46), .A3(new_n690_), .A4(new_n686_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n695_), .A2(new_n699_), .ZN(G1329gat));
  INV_X1    g499(.A(G43gat), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n509_), .A2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n673_), .A2(new_n678_), .A3(new_n702_), .ZN(new_n703_));
  AOI211_X1 g502(.A(KEYINPUT114), .B(G43gat), .C1(new_n663_), .C2(new_n576_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT114), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n663_), .A2(new_n576_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n706_), .B2(new_n701_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n703_), .B1(new_n704_), .B2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(KEYINPUT47), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT47), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n703_), .B(new_n710_), .C1(new_n704_), .C2(new_n707_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n711_), .ZN(G1330gat));
  AOI21_X1  g511(.A(G50gat), .B1(new_n663_), .B2(new_n652_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n673_), .A2(G50gat), .A3(new_n652_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n714_), .B2(new_n678_), .ZN(G1331gat));
  INV_X1    g514(.A(KEYINPUT115), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n661_), .A2(new_n716_), .A3(new_n376_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n376_), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT115), .B1(new_n307_), .B2(new_n718_), .ZN(new_n719_));
  NOR4_X1   g518(.A1(new_n717_), .A2(new_n600_), .A3(new_n719_), .A4(new_n578_), .ZN(new_n720_));
  INV_X1    g519(.A(G57gat), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n720_), .A2(new_n721_), .A3(new_n616_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n307_), .A2(new_n601_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n626_), .A2(new_n658_), .A3(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(G57gat), .B1(new_n725_), .B2(new_n607_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n722_), .A2(new_n726_), .ZN(G1332gat));
  INV_X1    g526(.A(G64gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n724_), .B2(new_n606_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT48), .Z(new_n730_));
  NAND3_X1  g529(.A1(new_n720_), .A2(new_n728_), .A3(new_n606_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1333gat));
  INV_X1    g531(.A(G71gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n724_), .B2(new_n576_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT49), .Z(new_n735_));
  NAND3_X1  g534(.A1(new_n720_), .A2(new_n733_), .A3(new_n576_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1334gat));
  AOI21_X1  g536(.A(new_n204_), .B1(new_n724_), .B2(new_n652_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT50), .Z(new_n739_));
  NAND3_X1  g538(.A1(new_n720_), .A2(new_n204_), .A3(new_n652_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1335gat));
  INV_X1    g540(.A(new_n723_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n675_), .A2(new_n671_), .A3(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(G85gat), .B1(new_n743_), .B2(new_n607_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n660_), .A2(new_n611_), .ZN(new_n745_));
  OR3_X1    g544(.A1(new_n745_), .A2(KEYINPUT116), .A3(new_n723_), .ZN(new_n746_));
  OAI21_X1  g545(.A(KEYINPUT116), .B1(new_n745_), .B2(new_n723_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n616_), .A2(new_n234_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n744_), .B1(new_n749_), .B2(new_n750_), .ZN(G1336gat));
  OAI21_X1  g550(.A(G92gat), .B1(new_n743_), .B2(new_n565_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n606_), .A2(new_n235_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n752_), .B1(new_n749_), .B2(new_n753_), .ZN(G1337gat));
  OAI21_X1  g553(.A(G99gat), .B1(new_n743_), .B2(new_n516_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT117), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n509_), .A2(new_n228_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n748_), .B2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n757_), .ZN(new_n759_));
  AOI211_X1 g558(.A(KEYINPUT117), .B(new_n759_), .C1(new_n746_), .C2(new_n747_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n755_), .B1(new_n758_), .B2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(KEYINPUT118), .A3(KEYINPUT51), .ZN(new_n762_));
  NAND2_X1  g561(.A1(KEYINPUT118), .A2(KEYINPUT51), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n763_), .B(new_n755_), .C1(new_n758_), .C2(new_n760_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(G1338gat));
  NAND3_X1  g564(.A1(new_n748_), .A2(new_n446_), .A3(new_n652_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n675_), .A2(new_n652_), .A3(new_n671_), .A4(new_n742_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n767_), .A2(new_n768_), .A3(G106gat), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(new_n767_), .B2(G106gat), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n766_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g571(.A1(new_n616_), .A2(new_n565_), .A3(new_n609_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n287_), .A2(new_n292_), .ZN(new_n774_));
  OR2_X1    g573(.A1(new_n774_), .A2(new_n297_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n587_), .A2(new_n580_), .A3(new_n588_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n580_), .B1(new_n326_), .B2(new_n342_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n579_), .A2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n776_), .A2(new_n598_), .A3(new_n778_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n594_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n775_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n217_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n782_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n284_), .A2(new_n216_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n289_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n291_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT121), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n287_), .A2(new_n788_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n277_), .A2(new_n285_), .A3(KEYINPUT55), .A4(new_n286_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT121), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n791_), .B(new_n291_), .C1(new_n783_), .C2(new_n785_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n787_), .A2(new_n789_), .A3(new_n790_), .A4(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n297_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT56), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n793_), .A2(KEYINPUT56), .A3(new_n297_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n781_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT123), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n799_), .A2(KEYINPUT58), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n665_), .B1(new_n798_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n781_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n793_), .A2(KEYINPUT56), .A3(new_n297_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT56), .B1(new_n793_), .B2(new_n297_), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n801_), .B(new_n803_), .C1(new_n804_), .C2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n600_), .A2(new_n775_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n809_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n780_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n624_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(KEYINPUT122), .A2(KEYINPUT57), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  OAI22_X1  g613(.A1(new_n802_), .A2(new_n807_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n808_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n811_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n625_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n818_), .A2(new_n813_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n627_), .B1(new_n815_), .B2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n601_), .A2(new_n302_), .A3(new_n304_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT54), .B1(new_n376_), .B2(new_n821_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(KEYINPUT120), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n601_), .A2(new_n302_), .A3(new_n304_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n824_), .A2(new_n667_), .A3(new_n825_), .A4(new_n332_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT119), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n718_), .A2(new_n824_), .A3(KEYINPUT119), .A4(new_n825_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n823_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n773_), .B1(new_n820_), .B2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(G113gat), .B1(new_n831_), .B2(new_n600_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n773_), .A2(KEYINPUT59), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n803_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n667_), .B1(new_n834_), .B2(new_n800_), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n818_), .A2(new_n813_), .B1(new_n835_), .B2(new_n806_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n812_), .A2(new_n814_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n332_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n828_), .A2(new_n829_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n822_), .A2(KEYINPUT120), .ZN(new_n840_));
  OR2_X1    g639(.A1(new_n822_), .A2(KEYINPUT120), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n839_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n833_), .B1(new_n838_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n831_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT124), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT124), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n843_), .B(new_n847_), .C1(new_n831_), .C2(new_n844_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n600_), .A2(G113gat), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n832_), .B1(new_n849_), .B2(new_n850_), .ZN(G1340gat));
  OAI21_X1  g650(.A(G120gat), .B1(new_n845_), .B2(new_n661_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n831_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT60), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n307_), .A2(new_n854_), .ZN(new_n855_));
  MUX2_X1   g654(.A(new_n855_), .B(new_n854_), .S(G120gat), .Z(new_n856_));
  OAI21_X1  g655(.A(new_n852_), .B1(new_n853_), .B2(new_n856_), .ZN(G1341gat));
  AOI21_X1  g656(.A(G127gat), .B1(new_n831_), .B2(new_n332_), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n331_), .A2(G127gat), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n858_), .B1(new_n849_), .B2(new_n859_), .ZN(G1342gat));
  AOI21_X1  g659(.A(G134gat), .B1(new_n831_), .B2(new_n624_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(KEYINPUT125), .B(G134gat), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n667_), .A2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n861_), .B1(new_n849_), .B2(new_n863_), .ZN(G1343gat));
  NAND2_X1  g663(.A1(new_n820_), .A2(new_n830_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n606_), .A2(new_n615_), .A3(new_n517_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(KEYINPUT126), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n601_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(new_n384_), .ZN(G1344gat));
  NOR2_X1   g669(.A1(new_n868_), .A2(new_n661_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(new_n385_), .ZN(G1345gat));
  NOR2_X1   g671(.A1(new_n868_), .A2(new_n658_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT61), .B(G155gat), .ZN(new_n874_));
  XOR2_X1   g673(.A(new_n873_), .B(new_n874_), .Z(G1346gat));
  OAI21_X1  g674(.A(G162gat), .B1(new_n868_), .B2(new_n667_), .ZN(new_n876_));
  OR2_X1    g675(.A1(new_n625_), .A2(G162gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n868_), .B2(new_n877_), .ZN(G1347gat));
  OAI21_X1  g677(.A(new_n658_), .B1(new_n815_), .B2(new_n819_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n830_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n616_), .A2(new_n565_), .A3(new_n516_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n652_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n880_), .A2(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(G169gat), .B1(new_n884_), .B2(new_n601_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n886_), .ZN(new_n888_));
  OAI211_X1 g687(.A(G169gat), .B(new_n888_), .C1(new_n884_), .C2(new_n601_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n884_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n600_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n887_), .B(new_n889_), .C1(new_n523_), .C2(new_n891_), .ZN(G1348gat));
  AOI21_X1  g691(.A(G176gat), .B1(new_n890_), .B2(new_n307_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n820_), .A2(new_n830_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n894_), .A2(new_n652_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n882_), .A2(new_n475_), .A3(new_n661_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n893_), .B1(new_n895_), .B2(new_n896_), .ZN(G1349gat));
  NOR3_X1   g696(.A1(new_n884_), .A2(new_n525_), .A3(new_n627_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n895_), .A2(new_n332_), .A3(new_n881_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n484_), .ZN(G1350gat));
  OAI21_X1  g699(.A(G190gat), .B1(new_n884_), .B2(new_n667_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n624_), .A2(new_n482_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n884_), .B2(new_n902_), .ZN(G1351gat));
  NOR3_X1   g702(.A1(new_n565_), .A2(new_n517_), .A3(new_n430_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n894_), .A2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n600_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n307_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G204gat), .ZN(G1353gat));
  XNOR2_X1  g709(.A(KEYINPUT63), .B(G211gat), .ZN(new_n911_));
  NOR4_X1   g710(.A1(new_n894_), .A2(new_n627_), .A3(new_n905_), .A4(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n906_), .A2(new_n331_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n912_), .B1(new_n913_), .B2(new_n914_), .ZN(G1354gat));
  INV_X1    g714(.A(G218gat), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n906_), .A2(new_n916_), .A3(new_n624_), .ZN(new_n917_));
  NOR3_X1   g716(.A1(new_n894_), .A2(new_n667_), .A3(new_n905_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n918_), .B2(new_n916_), .ZN(G1355gat));
endmodule


