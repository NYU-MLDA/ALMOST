//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 1 0 1 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n889_, new_n891_, new_n892_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_;
  XNOR2_X1  g000(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G232gat), .A2(G233gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  INV_X1    g003(.A(KEYINPUT65), .ZN(new_n205_));
  AND3_X1   g004(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n206_));
  AOI21_X1  g005(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n205_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT6), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n211_), .A2(KEYINPUT65), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n208_), .A2(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(KEYINPUT10), .B(G99gat), .Z(new_n215_));
  INV_X1    g014(.A(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(G85gat), .A2(G92gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G85gat), .A2(G92gat), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .A4(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n222_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(new_n218_), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n214_), .A2(new_n217_), .A3(new_n223_), .A4(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT66), .ZN(new_n227_));
  AOI22_X1  g026(.A1(new_n208_), .A2(new_n213_), .B1(new_n218_), .B2(new_n224_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n228_), .A2(new_n229_), .A3(new_n223_), .A4(new_n217_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n227_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT7), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n233_), .B(new_n234_), .C1(G99gat), .C2(G106gat), .ZN(new_n235_));
  INV_X1    g034(.A(G99gat), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n236_), .B(new_n216_), .C1(KEYINPUT67), .C2(KEYINPUT7), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n206_), .A2(new_n207_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n220_), .A2(new_n222_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n242_), .A2(new_n243_), .A3(KEYINPUT8), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n220_), .A2(new_n222_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n245_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT8), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT68), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n244_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n241_), .A2(new_n247_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n250_), .B1(new_n214_), .B2(new_n238_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(KEYINPUT72), .B1(new_n249_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT72), .ZN(new_n254_));
  AOI211_X1 g053(.A(new_n254_), .B(new_n251_), .C1(new_n244_), .C2(new_n248_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n232_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G29gat), .B(G36gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G43gat), .B(G50gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n259_), .B(KEYINPUT15), .Z(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n251_), .B1(new_n244_), .B2(new_n248_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n262_), .A2(new_n231_), .ZN(new_n263_));
  AOI22_X1  g062(.A1(new_n256_), .A2(new_n261_), .B1(new_n259_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT35), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n204_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n263_), .A2(new_n259_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n243_), .B1(new_n242_), .B2(KEYINPUT8), .ZN(new_n268_));
  NOR3_X1   g067(.A1(new_n246_), .A2(KEYINPUT68), .A3(new_n247_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n252_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(new_n254_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n262_), .A2(KEYINPUT72), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n231_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n267_), .B1(new_n273_), .B2(new_n260_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT75), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n204_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n277_), .A2(KEYINPUT35), .ZN(new_n278_));
  NOR3_X1   g077(.A1(new_n266_), .A2(new_n276_), .A3(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n264_), .A2(KEYINPUT75), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n277_), .B1(new_n274_), .B2(KEYINPUT35), .ZN(new_n281_));
  INV_X1    g080(.A(new_n278_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n280_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT77), .B1(new_n279_), .B2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G134gat), .B(G162gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(G218gat), .ZN(new_n286_));
  XOR2_X1   g085(.A(KEYINPUT76), .B(G190gat), .Z(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT36), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n276_), .B1(new_n266_), .B2(new_n278_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT77), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n281_), .A2(new_n280_), .A3(new_n282_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n284_), .A2(new_n289_), .A3(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT36), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n290_), .A2(new_n292_), .A3(new_n295_), .A4(new_n288_), .ZN(new_n296_));
  AOI21_X1  g095(.A(KEYINPUT37), .B1(new_n294_), .B2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G1gat), .B(G8gat), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n298_), .A2(KEYINPUT78), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(KEYINPUT78), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G15gat), .B(G22gat), .ZN(new_n302_));
  INV_X1    g101(.A(G1gat), .ZN(new_n303_));
  INV_X1    g102(.A(G8gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT14), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n301_), .A2(new_n306_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n299_), .A2(new_n305_), .A3(new_n302_), .A4(new_n300_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G231gat), .A2(G233gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(G57gat), .B(G64gat), .Z(new_n312_));
  INV_X1    g111(.A(KEYINPUT11), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(KEYINPUT69), .B(G71gat), .Z(new_n315_));
  INV_X1    g114(.A(G78gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT69), .B(G71gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(G78gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n314_), .A2(new_n317_), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT70), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n318_), .B(new_n316_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT70), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n322_), .A2(new_n323_), .A3(new_n314_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n312_), .A2(new_n313_), .ZN(new_n325_));
  AND3_X1   g124(.A1(new_n321_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n325_), .B1(new_n321_), .B2(new_n324_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n311_), .B(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT17), .ZN(new_n330_));
  XOR2_X1   g129(.A(G183gat), .B(G211gat), .Z(new_n331_));
  XNOR2_X1  g130(.A(G127gat), .B(G155gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  NOR3_X1   g134(.A1(new_n329_), .A2(new_n330_), .A3(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(KEYINPUT17), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n329_), .A2(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n289_), .B1(new_n279_), .B2(new_n283_), .ZN(new_n341_));
  AND3_X1   g140(.A1(new_n341_), .A2(KEYINPUT37), .A3(new_n296_), .ZN(new_n342_));
  NOR3_X1   g141(.A1(new_n297_), .A2(new_n340_), .A3(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n343_), .B(KEYINPUT80), .Z(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT5), .B(G176gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(G204gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G120gat), .B(G148gat), .ZN(new_n347_));
  XOR2_X1   g146(.A(new_n346_), .B(new_n347_), .Z(new_n348_));
  INV_X1    g147(.A(KEYINPUT71), .ZN(new_n349_));
  INV_X1    g148(.A(new_n325_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n323_), .B1(new_n322_), .B2(new_n314_), .ZN(new_n351_));
  AND4_X1   g150(.A1(new_n323_), .A2(new_n314_), .A3(new_n317_), .A4(new_n319_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n350_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n321_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT12), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n256_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G230gat), .A2(G233gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n263_), .A2(new_n355_), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n354_), .B(new_n353_), .C1(new_n262_), .C2(new_n231_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n356_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n358_), .A2(new_n359_), .A3(new_n360_), .A4(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n360_), .A2(new_n361_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n359_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n349_), .B1(new_n363_), .B2(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(KEYINPUT71), .B1(new_n364_), .B2(new_n365_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n348_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT73), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n328_), .A2(KEYINPUT12), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n360_), .B(new_n362_), .C1(new_n273_), .C2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n366_), .B1(new_n372_), .B2(new_n365_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n368_), .B1(new_n373_), .B2(KEYINPUT71), .ZN(new_n374_));
  INV_X1    g173(.A(new_n348_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n370_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  NOR4_X1   g175(.A1(new_n367_), .A2(KEYINPUT73), .A3(new_n368_), .A4(new_n348_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n369_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n378_), .A2(KEYINPUT13), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(KEYINPUT13), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n309_), .A2(new_n259_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT81), .ZN(new_n383_));
  INV_X1    g182(.A(new_n309_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n383_), .B1(new_n384_), .B2(new_n261_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G229gat), .A2(G233gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n309_), .A2(new_n259_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n383_), .A2(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n387_), .B1(new_n386_), .B2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G113gat), .B(G141gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G169gat), .B(G197gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n390_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n393_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n387_), .B(new_n395_), .C1(new_n386_), .C2(new_n389_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n381_), .A2(new_n397_), .ZN(new_n398_));
  XOR2_X1   g197(.A(G15gat), .B(G43gat), .Z(new_n399_));
  XNOR2_X1  g198(.A(G71gat), .B(G99gat), .ZN(new_n400_));
  XOR2_X1   g199(.A(new_n399_), .B(new_n400_), .Z(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(G169gat), .ZN(new_n403_));
  INV_X1    g202(.A(G176gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G169gat), .A2(G176gat), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n405_), .A2(KEYINPUT24), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G183gat), .A2(G190gat), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT23), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n405_), .A2(KEYINPUT24), .ZN(new_n413_));
  NOR3_X1   g212(.A1(new_n407_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT25), .B(G183gat), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT26), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(G190gat), .ZN(new_n417_));
  OR2_X1    g216(.A1(KEYINPUT82), .A2(G190gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(KEYINPUT82), .A2(G190gat), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n416_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n415_), .B(new_n417_), .C1(new_n420_), .C2(KEYINPUT83), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n418_), .A2(new_n419_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n422_), .A2(KEYINPUT83), .A3(KEYINPUT26), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n414_), .B1(new_n421_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT22), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n426_), .A2(KEYINPUT84), .ZN(new_n427_));
  OAI21_X1  g226(.A(G169gat), .B1(new_n427_), .B2(G176gat), .ZN(new_n428_));
  AOI21_X1  g227(.A(G183gat), .B1(new_n418_), .B2(new_n419_), .ZN(new_n429_));
  OAI221_X1 g228(.A(new_n428_), .B1(new_n405_), .B2(new_n427_), .C1(new_n429_), .C2(new_n412_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n425_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT30), .ZN(new_n432_));
  XOR2_X1   g231(.A(G113gat), .B(G120gat), .Z(new_n433_));
  XNOR2_X1  g232(.A(G127gat), .B(G134gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  OR2_X1    g234(.A1(new_n432_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n432_), .A2(new_n435_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G227gat), .A2(G233gat), .ZN(new_n438_));
  XOR2_X1   g237(.A(new_n438_), .B(KEYINPUT31), .Z(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n436_), .A2(new_n437_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n440_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n402_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n443_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(new_n401_), .A3(new_n441_), .ZN(new_n446_));
  XOR2_X1   g245(.A(G78gat), .B(G106gat), .Z(new_n447_));
  INV_X1    g246(.A(KEYINPUT21), .ZN(new_n448_));
  INV_X1    g247(.A(G204gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(G197gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT85), .B(G197gat), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n448_), .B(new_n450_), .C1(new_n451_), .C2(new_n449_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT87), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(G197gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT85), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT85), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(G197gat), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n456_), .A2(new_n458_), .A3(new_n449_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT86), .B1(new_n449_), .B2(G197gat), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT86), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(new_n455_), .A3(G204gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT21), .B1(new_n459_), .B2(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n457_), .A2(G197gat), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n455_), .A2(KEYINPUT85), .ZN(new_n466_));
  OAI21_X1  g265(.A(G204gat), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n467_), .A2(KEYINPUT87), .A3(new_n448_), .A4(new_n450_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G211gat), .B(G218gat), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n454_), .A2(new_n464_), .A3(new_n468_), .A4(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n469_), .B1(new_n467_), .B2(new_n450_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT21), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  AND3_X1   g272(.A1(KEYINPUT88), .A2(G228gat), .A3(G233gat), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT3), .ZN(new_n475_));
  INV_X1    g274(.A(G141gat), .ZN(new_n476_));
  INV_X1    g275(.A(G148gat), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G141gat), .A2(G148gat), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT2), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n478_), .A2(new_n481_), .A3(new_n482_), .A4(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G155gat), .A2(G162gat), .ZN(new_n485_));
  OR2_X1    g284(.A1(G155gat), .A2(G162gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n484_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n476_), .A2(new_n477_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n485_), .A2(KEYINPUT1), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(new_n486_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n485_), .A2(KEYINPUT1), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n488_), .B(new_n479_), .C1(new_n490_), .C2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n487_), .A2(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n474_), .B1(new_n493_), .B2(KEYINPUT29), .ZN(new_n494_));
  AOI21_X1  g293(.A(KEYINPUT88), .B1(G228gat), .B2(G233gat), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n473_), .A2(new_n494_), .A3(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n496_), .B1(new_n473_), .B2(new_n494_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n447_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT90), .ZN(new_n500_));
  OR3_X1    g299(.A1(new_n493_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT28), .B1(new_n493_), .B2(KEYINPUT29), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G22gat), .B(G50gat), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n501_), .A2(new_n502_), .A3(new_n504_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n500_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n499_), .A2(new_n508_), .A3(KEYINPUT89), .ZN(new_n511_));
  INV_X1    g310(.A(new_n498_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n473_), .A2(new_n494_), .A3(new_n496_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n447_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n512_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT91), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT91), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n512_), .A2(new_n517_), .A3(new_n513_), .A4(new_n514_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n510_), .A2(new_n511_), .A3(new_n516_), .A4(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n516_), .A2(new_n518_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n511_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n508_), .B1(KEYINPUT90), .B2(new_n499_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n520_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  AOI22_X1  g322(.A1(new_n444_), .A2(new_n446_), .B1(new_n519_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n493_), .A2(new_n435_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G113gat), .B(G120gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n434_), .B(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n528_), .A2(new_n492_), .A3(new_n487_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n526_), .A2(new_n529_), .A3(KEYINPUT4), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT94), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G225gat), .A2(G233gat), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n526_), .A2(KEYINPUT4), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT94), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n526_), .A2(new_n529_), .A3(new_n535_), .A4(KEYINPUT4), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n531_), .A2(new_n533_), .A3(new_n534_), .A4(new_n536_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n526_), .A2(new_n529_), .A3(KEYINPUT95), .A4(new_n532_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT95), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n526_), .A2(new_n529_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n539_), .B1(new_n540_), .B2(new_n533_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n537_), .A2(new_n538_), .A3(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G1gat), .B(G29gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(G85gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT0), .B(G57gat), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n544_), .B(new_n545_), .Z(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n542_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT99), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n537_), .A2(new_n546_), .A3(new_n538_), .A4(new_n541_), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n548_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n549_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT27), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G8gat), .B(G36gat), .ZN(new_n555_));
  INV_X1    g354(.A(G92gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT18), .B(G64gat), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n557_), .B(new_n558_), .Z(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT20), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n470_), .A2(new_n472_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(KEYINPUT26), .B(G190gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(new_n415_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n414_), .A2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(G183gat), .A2(G190gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT22), .B(G169gat), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  OAI221_X1 g367(.A(new_n406_), .B1(new_n412_), .B2(new_n566_), .C1(new_n568_), .C2(G176gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n565_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n561_), .B1(new_n562_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n473_), .A2(new_n431_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT93), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G226gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT19), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n473_), .A2(KEYINPUT93), .A3(new_n431_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n572_), .A2(new_n575_), .A3(new_n578_), .A4(new_n579_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n470_), .A2(new_n472_), .A3(new_n425_), .A4(new_n430_), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n581_), .A2(KEYINPUT92), .A3(KEYINPUT20), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT92), .B1(new_n581_), .B2(KEYINPUT20), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n473_), .A2(new_n570_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n582_), .A2(new_n583_), .A3(new_n585_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n560_), .B(new_n580_), .C1(new_n586_), .C2(new_n578_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n581_), .A2(KEYINPUT20), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT92), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n581_), .A2(KEYINPUT92), .A3(KEYINPUT20), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n591_), .A2(new_n584_), .A3(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(new_n577_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n560_), .B1(new_n594_), .B2(new_n580_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n554_), .B1(new_n588_), .B2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n572_), .A2(new_n575_), .A3(new_n579_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(new_n577_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n591_), .A2(new_n578_), .A3(new_n584_), .A4(new_n592_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  OAI211_X1 g399(.A(KEYINPUT27), .B(new_n587_), .C1(new_n600_), .C2(new_n560_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n596_), .A2(new_n601_), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n525_), .A2(new_n553_), .A3(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n596_), .A2(new_n601_), .ZN(new_n604_));
  OAI211_X1 g403(.A(new_n519_), .B(new_n523_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n604_), .A2(new_n606_), .A3(KEYINPUT100), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT100), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n608_), .B1(new_n602_), .B2(new_n605_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n523_), .A2(new_n519_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n580_), .B1(new_n586_), .B2(new_n578_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(new_n559_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n531_), .A2(new_n532_), .A3(new_n534_), .A4(new_n536_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n540_), .B(KEYINPUT97), .Z(new_n614_));
  OAI211_X1 g413(.A(new_n547_), .B(new_n613_), .C1(new_n614_), .C2(new_n532_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n612_), .A2(new_n587_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT96), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n550_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT33), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT33), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n550_), .A2(new_n617_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n616_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n560_), .A2(KEYINPUT32), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT98), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n626_), .B(new_n580_), .C1(new_n586_), .C2(new_n578_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n600_), .A2(new_n625_), .A3(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n624_), .B1(new_n611_), .B2(new_n626_), .ZN(new_n629_));
  AOI22_X1  g428(.A1(new_n628_), .A2(new_n629_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n610_), .B1(new_n623_), .B2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n607_), .A2(new_n609_), .A3(new_n631_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n444_), .A2(new_n446_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n603_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n398_), .A2(new_n634_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n344_), .A2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n636_), .A2(new_n303_), .A3(new_n553_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT38), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n294_), .A2(new_n296_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n634_), .A2(new_n641_), .A3(new_n340_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n642_), .A2(new_n397_), .A3(new_n381_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n553_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G1gat), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n636_), .A2(KEYINPUT38), .A3(new_n303_), .A4(new_n553_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n639_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT101), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(G1324gat));
  OAI21_X1  g448(.A(G8gat), .B1(new_n643_), .B2(new_n604_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n651_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(KEYINPUT39), .A3(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n636_), .A2(new_n304_), .A3(new_n602_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT39), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n650_), .A2(new_n651_), .A3(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n654_), .A2(new_n655_), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT40), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n654_), .A2(new_n655_), .A3(KEYINPUT40), .A4(new_n657_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1325gat));
  INV_X1    g461(.A(G15gat), .ZN(new_n663_));
  INV_X1    g462(.A(new_n633_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n636_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT103), .ZN(new_n666_));
  OAI21_X1  g465(.A(G15gat), .B1(new_n643_), .B2(new_n633_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT41), .Z(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(G1326gat));
  INV_X1    g468(.A(G22gat), .ZN(new_n670_));
  INV_X1    g469(.A(new_n610_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n636_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(G22gat), .B1(new_n643_), .B2(new_n610_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n673_), .A2(KEYINPUT42), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(KEYINPUT42), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n672_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT104), .ZN(G1327gat));
  NOR4_X1   g476(.A1(new_n398_), .A2(new_n640_), .A3(new_n634_), .A4(new_n339_), .ZN(new_n678_));
  AOI21_X1  g477(.A(G29gat), .B1(new_n678_), .B2(new_n553_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n297_), .A2(new_n342_), .ZN(new_n680_));
  OAI21_X1  g479(.A(KEYINPUT105), .B1(new_n634_), .B2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT43), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n683_));
  OAI211_X1 g482(.A(KEYINPUT105), .B(new_n683_), .C1(new_n634_), .C2(new_n680_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n398_), .A2(new_n339_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n682_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n682_), .A2(KEYINPUT44), .A3(new_n685_), .A4(new_n684_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT106), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n689_), .A2(new_n690_), .ZN(new_n692_));
  OAI211_X1 g491(.A(G29gat), .B(new_n688_), .C1(new_n691_), .C2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n679_), .B1(new_n694_), .B2(new_n553_), .ZN(G1328gat));
  XNOR2_X1  g494(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n602_), .B(new_n688_), .C1(new_n691_), .C2(new_n692_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(G36gat), .ZN(new_n698_));
  INV_X1    g497(.A(G36gat), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n640_), .A2(new_n339_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n635_), .A2(new_n699_), .A3(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(KEYINPUT45), .B1(new_n701_), .B2(new_n604_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT45), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n678_), .A2(new_n703_), .A3(new_n699_), .A4(new_n602_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n696_), .B1(new_n698_), .B2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n696_), .ZN(new_n708_));
  AOI211_X1 g507(.A(new_n705_), .B(new_n708_), .C1(new_n697_), .C2(G36gat), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n707_), .A2(new_n709_), .ZN(G1329gat));
  INV_X1    g509(.A(G43gat), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n633_), .A2(new_n711_), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n688_), .B(new_n712_), .C1(new_n691_), .C2(new_n692_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n678_), .A2(new_n664_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g516(.A(G50gat), .B1(new_n678_), .B2(new_n671_), .ZN(new_n718_));
  OAI211_X1 g517(.A(G50gat), .B(new_n688_), .C1(new_n691_), .C2(new_n692_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n718_), .B1(new_n720_), .B2(new_n671_), .ZN(G1331gat));
  INV_X1    g520(.A(G57gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(new_n553_), .B2(KEYINPUT110), .ZN(new_n723_));
  INV_X1    g522(.A(new_n397_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n381_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n642_), .A2(new_n724_), .A3(new_n725_), .ZN(new_n726_));
  AOI211_X1 g525(.A(new_n723_), .B(new_n726_), .C1(KEYINPUT110), .C2(new_n722_), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n634_), .A2(new_n397_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT109), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT108), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n344_), .A2(new_n731_), .A3(new_n725_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n731_), .B1(new_n344_), .B2(new_n725_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n730_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n735_), .A2(new_n644_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n727_), .B1(new_n736_), .B2(new_n722_), .ZN(G1332gat));
  OAI21_X1  g536(.A(G64gat), .B1(new_n726_), .B2(new_n604_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT48), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n604_), .A2(G64gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n735_), .B2(new_n740_), .ZN(G1333gat));
  OAI21_X1  g540(.A(G71gat), .B1(new_n726_), .B2(new_n633_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT49), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n633_), .A2(G71gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n735_), .B2(new_n744_), .ZN(G1334gat));
  OAI21_X1  g544(.A(G78gat), .B1(new_n726_), .B2(new_n610_), .ZN(new_n746_));
  XOR2_X1   g545(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n747_));
  XNOR2_X1  g546(.A(new_n746_), .B(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n671_), .A2(new_n316_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n735_), .B2(new_n749_), .ZN(G1335gat));
  NOR2_X1   g549(.A1(new_n729_), .A2(new_n381_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n751_), .A2(new_n700_), .ZN(new_n752_));
  AOI21_X1  g551(.A(G85gat), .B1(new_n752_), .B2(new_n553_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n381_), .A2(new_n397_), .A3(new_n339_), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n682_), .A2(new_n684_), .A3(new_n754_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n755_), .A2(G85gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n753_), .B1(new_n553_), .B2(new_n756_), .ZN(G1336gat));
  AOI21_X1  g556(.A(G92gat), .B1(new_n752_), .B2(new_n602_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n604_), .A2(new_n556_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n755_), .B2(new_n759_), .ZN(G1337gat));
  AND2_X1   g559(.A1(new_n664_), .A2(new_n215_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n751_), .A2(new_n700_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n682_), .A2(new_n664_), .A3(new_n684_), .A4(new_n754_), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT112), .B1(new_n764_), .B2(G99gat), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n764_), .A2(KEYINPUT112), .A3(G99gat), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n762_), .B(new_n763_), .C1(new_n765_), .C2(new_n766_), .ZN(new_n767_));
  OR2_X1    g566(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n767_), .B(new_n768_), .ZN(G1338gat));
  NAND4_X1  g568(.A1(new_n682_), .A2(new_n671_), .A3(new_n684_), .A4(new_n754_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(G106gat), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT114), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n770_), .A2(new_n773_), .A3(G106gat), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n772_), .A2(KEYINPUT52), .A3(new_n774_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n751_), .A2(new_n216_), .A3(new_n671_), .A4(new_n700_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n771_), .A2(KEYINPUT114), .A3(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n775_), .A2(new_n776_), .A3(new_n778_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g579(.A(new_n386_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n393_), .B1(new_n389_), .B2(new_n781_), .ZN(new_n782_));
  OR2_X1    g581(.A1(new_n782_), .A2(KEYINPUT117), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n385_), .A2(new_n781_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(KEYINPUT117), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n783_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n396_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n378_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n372_), .B2(new_n365_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n372_), .A2(new_n365_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n372_), .A2(new_n790_), .A3(new_n365_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n348_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n795_), .A2(new_n798_), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n799_), .B(new_n397_), .C1(new_n376_), .C2(new_n377_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n797_), .B(new_n348_), .C1(new_n793_), .C2(new_n794_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT56), .B1(new_n801_), .B2(KEYINPUT116), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n789_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n803_), .A2(KEYINPUT57), .A3(new_n640_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT118), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n803_), .A2(new_n640_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  OR2_X1    g608(.A1(new_n297_), .A2(new_n342_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT58), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n788_), .B1(KEYINPUT56), .B2(new_n795_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n795_), .A2(KEYINPUT56), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n811_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n795_), .A2(KEYINPUT56), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n816_), .A2(new_n787_), .ZN(new_n817_));
  OR2_X1    g616(.A1(new_n376_), .A2(new_n377_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n817_), .A2(new_n818_), .A3(KEYINPUT58), .A4(new_n813_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n810_), .A2(new_n815_), .A3(new_n819_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n803_), .A2(KEYINPUT118), .A3(KEYINPUT57), .A4(new_n640_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n806_), .A2(new_n809_), .A3(new_n820_), .A4(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n343_), .A2(new_n381_), .A3(new_n724_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT54), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n343_), .A2(new_n381_), .A3(new_n825_), .A4(new_n724_), .ZN(new_n826_));
  AOI22_X1  g625(.A1(new_n822_), .A2(new_n340_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n602_), .A2(new_n644_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n829_), .A2(new_n525_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  OR3_X1    g630(.A1(new_n827_), .A2(KEYINPUT59), .A3(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT59), .B1(new_n827_), .B2(new_n831_), .ZN(new_n833_));
  AND4_X1   g632(.A1(G113gat), .A2(new_n832_), .A3(new_n397_), .A4(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n822_), .A2(new_n340_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n824_), .A2(new_n826_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT119), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(new_n838_), .A3(new_n830_), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT119), .B1(new_n827_), .B2(new_n831_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(G113gat), .B1(new_n841_), .B2(new_n397_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n834_), .A2(new_n842_), .ZN(G1340gat));
  NAND3_X1  g642(.A1(new_n832_), .A2(new_n725_), .A3(new_n833_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(KEYINPUT120), .B(G120gat), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n845_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n381_), .B2(KEYINPUT60), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n841_), .B(new_n848_), .C1(KEYINPUT60), .C2(new_n847_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n846_), .A2(new_n849_), .ZN(G1341gat));
  AOI21_X1  g649(.A(G127gat), .B1(new_n841_), .B2(new_n339_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n832_), .A2(new_n833_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n339_), .A2(G127gat), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n851_), .B1(new_n852_), .B2(new_n853_), .ZN(G1342gat));
  AOI21_X1  g653(.A(G134gat), .B1(new_n841_), .B2(new_n641_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n810_), .A2(G134gat), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n855_), .B1(new_n852_), .B2(new_n856_), .ZN(G1343gat));
  NOR2_X1   g656(.A1(new_n827_), .A2(new_n829_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n664_), .A2(new_n610_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(new_n724_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(new_n476_), .ZN(G1344gat));
  NOR2_X1   g661(.A1(new_n860_), .A2(new_n381_), .ZN(new_n863_));
  XOR2_X1   g662(.A(KEYINPUT121), .B(G148gat), .Z(new_n864_));
  XNOR2_X1  g663(.A(new_n863_), .B(new_n864_), .ZN(G1345gat));
  NAND4_X1  g664(.A1(new_n837_), .A2(new_n339_), .A3(new_n828_), .A4(new_n859_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(KEYINPUT122), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n858_), .A2(new_n868_), .A3(new_n339_), .A4(new_n859_), .ZN(new_n869_));
  XOR2_X1   g668(.A(KEYINPUT61), .B(G155gat), .Z(new_n870_));
  AND3_X1   g669(.A1(new_n867_), .A2(new_n869_), .A3(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n867_), .B2(new_n869_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1346gat));
  INV_X1    g672(.A(G162gat), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n860_), .A2(new_n874_), .A3(new_n680_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n858_), .A2(new_n641_), .A3(new_n859_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n874_), .B2(new_n876_), .ZN(G1347gat));
  NOR3_X1   g676(.A1(new_n525_), .A2(new_n604_), .A3(new_n553_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n837_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n397_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n881_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT62), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n879_), .A2(new_n724_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n884_), .B2(new_n403_), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n882_), .B(new_n885_), .C1(new_n568_), .C2(new_n881_), .ZN(G1348gat));
  NOR2_X1   g685(.A1(new_n879_), .A2(new_n381_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(new_n404_), .ZN(G1349gat));
  NOR2_X1   g687(.A1(new_n879_), .A2(new_n340_), .ZN(new_n889_));
  MUX2_X1   g688(.A(G183gat), .B(new_n415_), .S(new_n889_), .Z(G1350gat));
  OAI21_X1  g689(.A(G190gat), .B1(new_n879_), .B2(new_n680_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n641_), .A2(new_n563_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n879_), .B2(new_n892_), .ZN(G1351gat));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n664_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n837_), .A2(new_n894_), .A3(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n895_), .ZN(new_n897_));
  OAI21_X1  g696(.A(KEYINPUT123), .B1(new_n827_), .B2(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n724_), .B1(new_n896_), .B2(new_n898_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n455_), .ZN(G1352gat));
  AOI21_X1  g699(.A(new_n381_), .B1(new_n896_), .B2(new_n898_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n449_), .A2(KEYINPUT124), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(KEYINPUT125), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n901_), .B(new_n903_), .ZN(G1353gat));
  AOI21_X1  g703(.A(new_n340_), .B1(new_n896_), .B2(new_n898_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT126), .ZN(new_n906_));
  XOR2_X1   g705(.A(KEYINPUT63), .B(G211gat), .Z(new_n907_));
  NAND3_X1  g706(.A1(new_n905_), .A2(new_n906_), .A3(new_n907_), .ZN(new_n908_));
  OR2_X1    g707(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n909_));
  OAI21_X1  g708(.A(KEYINPUT126), .B1(new_n905_), .B2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n907_), .ZN(new_n911_));
  AOI211_X1 g710(.A(new_n340_), .B(new_n911_), .C1(new_n896_), .C2(new_n898_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n908_), .B1(new_n910_), .B2(new_n912_), .ZN(G1354gat));
  NAND2_X1  g712(.A1(new_n896_), .A2(new_n898_), .ZN(new_n914_));
  AOI21_X1  g713(.A(G218gat), .B1(new_n914_), .B2(new_n641_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n680_), .B1(new_n896_), .B2(new_n898_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n915_), .B1(G218gat), .B2(new_n916_), .ZN(G1355gat));
endmodule


