//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 1 0 1 1 1 0 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0 1 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n906_, new_n907_, new_n909_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_;
  XOR2_X1   g000(.A(G29gat), .B(G36gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G29gat), .B(G36gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G43gat), .B(G50gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT74), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G15gat), .B(G22gat), .ZN(new_n211_));
  INV_X1    g010(.A(G1gat), .ZN(new_n212_));
  INV_X1    g011(.A(G8gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT14), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G1gat), .B(G8gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n210_), .B(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G229gat), .A2(G233gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n210_), .A2(new_n217_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n208_), .B(KEYINPUT15), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(new_n217_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n224_), .A3(new_n219_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n221_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G113gat), .B(G141gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT75), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G169gat), .B(G197gat), .ZN(new_n229_));
  XOR2_X1   g028(.A(new_n228_), .B(new_n229_), .Z(new_n230_));
  NAND2_X1  g029(.A1(new_n226_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n230_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n221_), .A2(new_n225_), .A3(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT26), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(G190gat), .ZN(new_n237_));
  INV_X1    g036(.A(G190gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT26), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT76), .ZN(new_n241_));
  INV_X1    g040(.A(G183gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT25), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT25), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(G183gat), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n237_), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n241_), .B(new_n246_), .C1(KEYINPUT76), .C2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G183gat), .A2(G190gat), .ZN(new_n249_));
  AND2_X1   g048(.A1(KEYINPUT77), .A2(KEYINPUT23), .ZN(new_n250_));
  NOR2_X1   g049(.A1(KEYINPUT77), .A2(KEYINPUT23), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n249_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n249_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT23), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n252_), .A2(new_n255_), .ZN(new_n256_));
  OR2_X1    g055(.A1(G169gat), .A2(G176gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G169gat), .A2(G176gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(KEYINPUT24), .A3(new_n258_), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n257_), .A2(KEYINPUT24), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n248_), .A2(new_n256_), .A3(new_n259_), .A4(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n262_));
  INV_X1    g061(.A(G169gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n253_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n249_), .A2(new_n254_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(G183gat), .A2(G190gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n265_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n261_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G227gat), .A2(G233gat), .ZN(new_n272_));
  INV_X1    g071(.A(G15gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT30), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n271_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G71gat), .B(G99gat), .ZN(new_n277_));
  INV_X1    g076(.A(G43gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n276_), .B(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(G134gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(G127gat), .ZN(new_n282_));
  INV_X1    g081(.A(G127gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(G134gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(G120gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(G113gat), .ZN(new_n287_));
  INV_X1    g086(.A(G113gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(G120gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(KEYINPUT78), .B1(new_n285_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n285_), .A2(new_n290_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n282_), .A2(new_n284_), .A3(new_n287_), .A4(new_n289_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n291_), .B1(new_n294_), .B2(KEYINPUT78), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT31), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT79), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n280_), .A2(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n296_), .A2(new_n297_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n280_), .B1(new_n300_), .B2(new_n298_), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(G233gat), .ZN(new_n303_));
  NOR2_X1   g102(.A1(KEYINPUT81), .A2(G228gat), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(KEYINPUT81), .A2(G228gat), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n303_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT3), .ZN(new_n308_));
  INV_X1    g107(.A(G141gat), .ZN(new_n309_));
  INV_X1    g108(.A(G148gat), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n308_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G141gat), .A2(G148gat), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT2), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n311_), .A2(new_n314_), .A3(new_n315_), .A4(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(G155gat), .B(G162gat), .Z(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  AND2_X1   g118(.A1(G141gat), .A2(G148gat), .ZN(new_n320_));
  NOR2_X1   g119(.A1(G141gat), .A2(G148gat), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G155gat), .B(G162gat), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n322_), .B(new_n323_), .C1(new_n324_), .C2(KEYINPUT1), .ZN(new_n325_));
  AND3_X1   g124(.A1(new_n319_), .A2(KEYINPUT80), .A3(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(KEYINPUT80), .B1(new_n319_), .B2(new_n325_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n307_), .B1(new_n328_), .B2(KEYINPUT29), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT85), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT21), .ZN(new_n331_));
  INV_X1    g130(.A(G197gat), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n332_), .A2(G204gat), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n331_), .B1(new_n333_), .B2(KEYINPUT82), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT83), .ZN(new_n335_));
  INV_X1    g134(.A(G204gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(G197gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n332_), .A2(G204gat), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT82), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n334_), .A2(new_n335_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(G218gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(G211gat), .ZN(new_n343_));
  INV_X1    g142(.A(G211gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(G218gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G197gat), .B(G204gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT84), .B(KEYINPUT21), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n346_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n341_), .A2(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n335_), .B1(new_n334_), .B2(new_n340_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n330_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n334_), .A2(new_n340_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT83), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n354_), .A2(KEYINPUT85), .A3(new_n341_), .A4(new_n349_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n352_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n346_), .ZN(new_n357_));
  NOR3_X1   g156(.A1(new_n357_), .A2(new_n331_), .A3(new_n347_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n356_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n329_), .A2(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n358_), .B1(new_n352_), .B2(new_n355_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n316_), .ZN(new_n363_));
  NOR3_X1   g162(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n315_), .ZN(new_n366_));
  AOI21_X1  g165(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n324_), .B1(new_n365_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n309_), .A2(new_n310_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(new_n323_), .A3(new_n312_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT1), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n371_), .B1(new_n318_), .B2(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n369_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT29), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n307_), .B1(new_n362_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n361_), .A2(new_n377_), .ZN(new_n378_));
  XOR2_X1   g177(.A(G78gat), .B(G106gat), .Z(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n379_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n361_), .A2(new_n377_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n328_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT28), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT80), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n386_), .B1(new_n369_), .B2(new_n373_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n319_), .A2(KEYINPUT80), .A3(new_n325_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n385_), .B1(new_n389_), .B2(new_n375_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G22gat), .B(G50gat), .ZN(new_n391_));
  OR3_X1    g190(.A1(new_n384_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n391_), .B1(new_n384_), .B2(new_n390_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n383_), .A2(new_n394_), .ZN(new_n395_));
  AOI22_X1  g194(.A1(new_n380_), .A2(new_n382_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G8gat), .B(G36gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT18), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G64gat), .B(G92gat), .ZN(new_n401_));
  XOR2_X1   g200(.A(new_n400_), .B(new_n401_), .Z(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G226gat), .A2(G233gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT19), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT20), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n243_), .A2(new_n245_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n266_), .B(new_n267_), .C1(new_n240_), .C2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n260_), .A2(new_n259_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n269_), .B1(new_n252_), .B2(new_n255_), .ZN(new_n411_));
  OAI22_X1  g210(.A1(new_n409_), .A2(new_n410_), .B1(new_n411_), .B2(new_n264_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n407_), .B1(new_n360_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n271_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(new_n362_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n406_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n412_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n356_), .A2(new_n359_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT20), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n406_), .B1(new_n414_), .B2(new_n362_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n403_), .B1(new_n416_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n360_), .A2(new_n271_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n423_), .A2(KEYINPUT20), .A3(new_n406_), .A4(new_n418_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n415_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT20), .B1(new_n362_), .B2(new_n417_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n402_), .B(new_n424_), .C1(new_n427_), .C2(new_n406_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n422_), .A2(new_n428_), .A3(KEYINPUT86), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n424_), .B1(new_n427_), .B2(new_n406_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT86), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n430_), .A2(new_n431_), .A3(new_n403_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n429_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G1gat), .B(G29gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(G85gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT0), .B(G57gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G225gat), .A2(G233gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n294_), .A2(KEYINPUT88), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT88), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n292_), .A2(new_n441_), .A3(new_n293_), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n374_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT87), .B1(new_n328_), .B2(new_n295_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n387_), .A2(new_n295_), .A3(KEYINPUT87), .A4(new_n388_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  OAI211_X1 g246(.A(KEYINPUT4), .B(new_n444_), .C1(new_n445_), .C2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n387_), .A2(new_n388_), .A3(new_n295_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(KEYINPUT89), .A2(KEYINPUT4), .ZN(new_n450_));
  AND2_X1   g249(.A1(KEYINPUT89), .A2(KEYINPUT4), .ZN(new_n451_));
  NOR3_X1   g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n439_), .B1(new_n448_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT87), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n449_), .A2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n443_), .B1(new_n456_), .B2(new_n446_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n439_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  OAI211_X1 g258(.A(KEYINPUT33), .B(new_n438_), .C1(new_n454_), .C2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT92), .ZN(new_n461_));
  AOI211_X1 g260(.A(new_n439_), .B(new_n443_), .C1(new_n456_), .C2(new_n446_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n461_), .B1(new_n462_), .B2(new_n438_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n457_), .A2(new_n458_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n464_), .A2(KEYINPUT92), .A3(new_n437_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n448_), .A2(new_n439_), .A3(new_n453_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n463_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n460_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT91), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT4), .ZN(new_n470_));
  AOI211_X1 g269(.A(new_n470_), .B(new_n443_), .C1(new_n456_), .C2(new_n446_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n458_), .B1(new_n471_), .B2(new_n452_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n459_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n437_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT90), .B(KEYINPUT33), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n469_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n438_), .B1(new_n454_), .B2(new_n459_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n475_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(KEYINPUT91), .A3(new_n478_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n433_), .A2(new_n468_), .A3(new_n476_), .A4(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n472_), .A2(new_n437_), .A3(new_n473_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(new_n477_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n430_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n402_), .A2(KEYINPUT32), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  AOI211_X1 g284(.A(new_n358_), .B(new_n412_), .C1(new_n352_), .C2(new_n355_), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT93), .B1(new_n486_), .B2(new_n407_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT93), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n418_), .A2(new_n488_), .A3(KEYINPUT20), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n489_), .A3(new_n423_), .ZN(new_n490_));
  AND3_X1   g289(.A1(new_n490_), .A2(KEYINPUT94), .A3(new_n405_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n360_), .A2(new_n412_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n492_), .A2(KEYINPUT20), .A3(new_n406_), .A4(new_n415_), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n490_), .A2(new_n405_), .B1(KEYINPUT94), .B2(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n491_), .A2(new_n494_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n482_), .B(new_n485_), .C1(new_n495_), .C2(new_n484_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n398_), .B1(new_n480_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT27), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n429_), .A2(new_n498_), .A3(new_n432_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n428_), .A2(KEYINPUT27), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n490_), .A2(KEYINPUT94), .A3(new_n405_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n414_), .A2(new_n362_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n502_), .B1(new_n419_), .B2(KEYINPUT93), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n406_), .B1(new_n503_), .B2(new_n489_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n493_), .A2(KEYINPUT94), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n501_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n500_), .B1(new_n506_), .B2(new_n403_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n477_), .B(new_n481_), .C1(new_n395_), .C2(new_n396_), .ZN(new_n508_));
  NOR3_X1   g307(.A1(new_n499_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n302_), .B1(new_n497_), .B2(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n302_), .A2(new_n482_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n403_), .B1(new_n491_), .B2(new_n494_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n500_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n429_), .A2(new_n498_), .A3(new_n432_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n514_), .A2(KEYINPUT95), .A3(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT95), .B1(new_n514_), .B2(new_n515_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n397_), .B(new_n511_), .C1(new_n516_), .C2(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n235_), .B1(new_n510_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT64), .ZN(new_n520_));
  OR2_X1    g319(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n521_));
  INV_X1    g320(.A(G106gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(G85gat), .ZN(new_n525_));
  INV_X1    g324(.A(G92gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G85gat), .A2(G92gat), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n527_), .A2(KEYINPUT9), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n524_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT6), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n531_), .B1(G99gat), .B2(G106gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G99gat), .A2(G106gat), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n533_), .A2(KEYINPUT6), .ZN(new_n534_));
  OAI22_X1  g333(.A1(new_n532_), .A2(new_n534_), .B1(KEYINPUT9), .B2(new_n528_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n520_), .B1(new_n530_), .B2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n528_), .A2(KEYINPUT9), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n533_), .A2(KEYINPUT6), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n531_), .A2(G99gat), .A3(G106gat), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n537_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n540_), .A2(KEYINPUT64), .A3(new_n524_), .A4(new_n529_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n536_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G57gat), .B(G64gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G71gat), .B(G78gat), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(new_n544_), .A3(KEYINPUT11), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(KEYINPUT11), .ZN(new_n546_));
  INV_X1    g345(.A(new_n544_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n543_), .A2(KEYINPUT11), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n545_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n527_), .A2(new_n528_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n532_), .A2(new_n534_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT7), .ZN(new_n553_));
  INV_X1    g352(.A(G99gat), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(new_n554_), .A3(new_n522_), .ZN(new_n555_));
  OAI21_X1  g354(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n551_), .B1(new_n552_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT8), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  OAI211_X1 g359(.A(KEYINPUT8), .B(new_n551_), .C1(new_n552_), .C2(new_n557_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n542_), .A2(new_n550_), .A3(new_n560_), .A4(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(KEYINPUT67), .B(KEYINPUT12), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n543_), .A2(KEYINPUT11), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n565_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n536_), .A2(new_n541_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n560_), .A2(new_n561_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n545_), .B(new_n566_), .C1(new_n567_), .C2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n564_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT65), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n571_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n542_), .A2(KEYINPUT65), .A3(new_n560_), .A4(new_n561_), .ZN(new_n573_));
  OAI211_X1 g372(.A(KEYINPUT66), .B(new_n545_), .C1(new_n548_), .C2(new_n549_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(KEYINPUT12), .ZN(new_n575_));
  AOI21_X1  g374(.A(KEYINPUT66), .B1(new_n566_), .B2(new_n545_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n572_), .A2(new_n573_), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G230gat), .A2(G233gat), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n570_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n569_), .A2(new_n562_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n581_), .A2(G230gat), .A3(G233gat), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(G120gat), .B(G148gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G176gat), .B(G204gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n583_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n580_), .A2(new_n582_), .A3(new_n588_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT13), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT13), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n590_), .A2(new_n594_), .A3(new_n591_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(KEYINPUT71), .B(KEYINPUT37), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n572_), .A2(new_n223_), .A3(new_n573_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT70), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n542_), .A2(new_n208_), .A3(new_n560_), .A4(new_n561_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G232gat), .A2(G233gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT34), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n604_), .A2(KEYINPUT35), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n599_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n604_), .A2(KEYINPUT35), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT69), .Z(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n601_), .A2(new_n607_), .A3(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G190gat), .B(G218gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G134gat), .B(G162gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n614_), .A2(KEYINPUT36), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n599_), .B(new_n606_), .C1(new_n600_), .C2(new_n609_), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n611_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n614_), .B(KEYINPUT36), .Z(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n619_), .B1(new_n611_), .B2(new_n616_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n598_), .B1(new_n617_), .B2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n611_), .A2(new_n616_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(new_n618_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n611_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n623_), .A2(new_n624_), .A3(new_n597_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n621_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G231gat), .A2(G233gat), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n550_), .B(new_n628_), .Z(new_n629_));
  XNOR2_X1  g428(.A(new_n217_), .B(KEYINPUT72), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  XOR2_X1   g431(.A(G127gat), .B(G155gat), .Z(new_n633_));
  XNOR2_X1  g432(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G183gat), .B(G211gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT17), .ZN(new_n638_));
  OR3_X1    g437(.A1(new_n637_), .A2(KEYINPUT66), .A3(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n637_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n639_), .B1(KEYINPUT17), .B2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n632_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n631_), .A2(new_n639_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n627_), .A2(new_n645_), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n519_), .A2(new_n596_), .A3(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n647_), .A2(new_n212_), .A3(new_n482_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT38), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n617_), .A2(new_n620_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n510_), .B2(new_n518_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n596_), .A2(new_n234_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n653_), .A2(new_n645_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT96), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n652_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n482_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G1gat), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n648_), .A2(new_n649_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n650_), .A2(new_n658_), .A3(new_n659_), .ZN(G1324gat));
  NOR2_X1   g459(.A1(new_n516_), .A2(new_n517_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n647_), .A2(new_n213_), .A3(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n652_), .A2(new_n661_), .A3(new_n655_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT97), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n652_), .A2(KEYINPUT97), .A3(new_n661_), .A4(new_n655_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n665_), .A2(G8gat), .A3(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT98), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT39), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT98), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n665_), .A2(new_n670_), .A3(G8gat), .A4(new_n666_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n668_), .A2(new_n669_), .A3(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n669_), .B1(new_n668_), .B2(new_n671_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n662_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n662_), .B(new_n675_), .C1(new_n672_), .C2(new_n673_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1325gat));
  INV_X1    g478(.A(new_n302_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n647_), .A2(new_n273_), .A3(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT100), .ZN(new_n682_));
  OAI21_X1  g481(.A(G15gat), .B1(new_n656_), .B2(new_n302_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT41), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n683_), .A2(KEYINPUT41), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n682_), .A2(new_n684_), .A3(new_n685_), .ZN(G1326gat));
  OAI21_X1  g485(.A(G22gat), .B1(new_n656_), .B2(new_n397_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT42), .ZN(new_n688_));
  INV_X1    g487(.A(G22gat), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n647_), .A2(new_n689_), .A3(new_n398_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(G1327gat));
  NOR2_X1   g490(.A1(new_n653_), .A2(new_n644_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n510_), .A2(new_n518_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n694_), .B2(new_n627_), .ZN(new_n695_));
  AOI211_X1 g494(.A(KEYINPUT43), .B(new_n626_), .C1(new_n510_), .C2(new_n518_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n692_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  OAI211_X1 g498(.A(KEYINPUT44), .B(new_n692_), .C1(new_n695_), .C2(new_n696_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(G29gat), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n701_), .A2(new_n702_), .A3(new_n657_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n596_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n651_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n704_), .A2(new_n644_), .A3(new_n705_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n519_), .A2(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(G29gat), .B1(new_n707_), .B2(new_n482_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n703_), .A2(new_n708_), .ZN(G1328gat));
  INV_X1    g508(.A(G36gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n707_), .A2(new_n710_), .A3(new_n661_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT45), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n699_), .A2(new_n661_), .A3(new_n700_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT101), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n713_), .A2(new_n714_), .A3(G36gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n713_), .B2(G36gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT46), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  OAI211_X1 g518(.A(KEYINPUT46), .B(new_n712_), .C1(new_n715_), .C2(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1329gat));
  INV_X1    g520(.A(new_n707_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n278_), .B1(new_n722_), .B2(new_n302_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n680_), .A2(G43gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n723_), .B1(new_n701_), .B2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g525(.A(G50gat), .B1(new_n701_), .B2(new_n397_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n397_), .A2(G50gat), .ZN(new_n728_));
  XOR2_X1   g527(.A(new_n728_), .B(KEYINPUT102), .Z(new_n729_));
  OAI21_X1  g528(.A(new_n727_), .B1(new_n722_), .B2(new_n729_), .ZN(G1331gat));
  NOR2_X1   g529(.A1(new_n596_), .A2(new_n234_), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n652_), .A2(new_n644_), .A3(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(G57gat), .B1(new_n733_), .B2(new_n657_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n731_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n735_), .B1(new_n510_), .B2(new_n518_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n736_), .A2(new_n646_), .ZN(new_n737_));
  INV_X1    g536(.A(G57gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n737_), .A2(new_n738_), .A3(new_n482_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n734_), .A2(new_n739_), .ZN(G1332gat));
  INV_X1    g539(.A(G64gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n732_), .B2(new_n661_), .ZN(new_n742_));
  XOR2_X1   g541(.A(KEYINPUT103), .B(KEYINPUT48), .Z(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n737_), .A2(new_n741_), .A3(new_n661_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1333gat));
  INV_X1    g545(.A(G71gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n732_), .B2(new_n680_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT49), .Z(new_n749_));
  NAND3_X1  g548(.A1(new_n737_), .A2(new_n747_), .A3(new_n680_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1334gat));
  INV_X1    g550(.A(G78gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(new_n732_), .B2(new_n398_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT50), .Z(new_n754_));
  NAND2_X1  g553(.A1(new_n398_), .A2(new_n752_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT104), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n737_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n754_), .A2(new_n757_), .ZN(G1335gat));
  OR2_X1    g557(.A1(new_n695_), .A2(new_n696_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n735_), .A2(new_n644_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(G85gat), .B1(new_n761_), .B2(new_n657_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n736_), .A2(new_n645_), .A3(new_n651_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n763_), .A2(new_n525_), .A3(new_n482_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT105), .ZN(G1336gat));
  NAND3_X1  g565(.A1(new_n763_), .A2(new_n526_), .A3(new_n661_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n759_), .A2(new_n661_), .A3(new_n760_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n767_), .B1(new_n769_), .B2(new_n526_), .ZN(G1337gat));
  OAI21_X1  g569(.A(G99gat), .B1(new_n761_), .B2(new_n302_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n763_), .A2(new_n680_), .A3(new_n521_), .A4(new_n523_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g573(.A(KEYINPUT108), .B(KEYINPUT53), .ZN(new_n775_));
  XNOR2_X1  g574(.A(KEYINPUT106), .B(KEYINPUT52), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n777_), .A2(KEYINPUT107), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n759_), .A2(new_n398_), .A3(new_n760_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n522_), .B1(new_n777_), .B2(KEYINPUT107), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n778_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n779_), .A2(new_n778_), .A3(new_n780_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n763_), .A2(new_n522_), .A3(new_n398_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n775_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n783_), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n785_), .B(new_n775_), .C1(new_n787_), .C2(new_n781_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n786_), .A2(new_n789_), .ZN(G1339gat));
  NAND2_X1  g589(.A1(new_n218_), .A2(new_n219_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n222_), .A2(new_n224_), .A3(new_n220_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n230_), .A3(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n791_), .A2(KEYINPUT112), .A3(new_n230_), .A4(new_n792_), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n795_), .A2(new_n233_), .A3(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n591_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n570_), .A2(new_n578_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n799_), .A2(KEYINPUT111), .A3(KEYINPUT55), .A4(new_n579_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n579_), .B1(new_n570_), .B2(new_n578_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n580_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n580_), .B2(new_n802_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n800_), .A2(new_n803_), .A3(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n589_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT56), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n806_), .A2(KEYINPUT56), .A3(new_n589_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n798_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n627_), .B1(new_n811_), .B2(KEYINPUT58), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n797_), .A2(new_n591_), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n806_), .A2(KEYINPUT56), .A3(new_n589_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT56), .B1(new_n806_), .B2(new_n589_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n813_), .B(KEYINPUT58), .C1(new_n814_), .C2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n234_), .A2(new_n591_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n818_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n797_), .A2(new_n592_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n651_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  OAI22_X1  g620(.A1(new_n812_), .A2(new_n817_), .B1(new_n821_), .B2(KEYINPUT57), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n821_), .A2(KEYINPUT57), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n645_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT110), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n626_), .A2(new_n596_), .A3(new_n235_), .A4(new_n644_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT109), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n825_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  AOI211_X1 g628(.A(KEYINPUT110), .B(KEYINPUT54), .C1(new_n826_), .C2(KEYINPUT109), .ZN(new_n830_));
  OAI22_X1  g629(.A1(new_n829_), .A2(new_n830_), .B1(KEYINPUT109), .B2(new_n826_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n827_), .A2(new_n828_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT110), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n826_), .A2(KEYINPUT109), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n827_), .A2(new_n825_), .A3(new_n828_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n833_), .A2(new_n834_), .A3(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n824_), .A2(new_n831_), .A3(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n661_), .A2(new_n398_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n302_), .A2(new_n657_), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n838_), .A2(KEYINPUT113), .A3(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT113), .B1(new_n838_), .B2(new_n839_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n837_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(G113gat), .B1(new_n844_), .B2(new_n234_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT114), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n837_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n843_), .A2(new_n847_), .A3(new_n848_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n837_), .B(new_n842_), .C1(new_n846_), .C2(KEYINPUT59), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n234_), .A2(G113gat), .ZN(new_n852_));
  XOR2_X1   g651(.A(new_n852_), .B(KEYINPUT115), .Z(new_n853_));
  AOI21_X1  g652(.A(new_n845_), .B1(new_n851_), .B2(new_n853_), .ZN(G1340gat));
  NOR2_X1   g653(.A1(new_n596_), .A2(G120gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n844_), .B1(KEYINPUT60), .B2(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n596_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(KEYINPUT116), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT116), .ZN(new_n859_));
  AOI211_X1 g658(.A(new_n859_), .B(new_n596_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n860_));
  OAI21_X1  g659(.A(G120gat), .B1(new_n858_), .B2(new_n860_), .ZN(new_n861_));
  OR2_X1    g660(.A1(new_n856_), .A2(KEYINPUT60), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1341gat));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n283_), .B1(new_n843_), .B2(new_n645_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(KEYINPUT117), .ZN(new_n866_));
  AOI211_X1 g665(.A(new_n283_), .B(new_n645_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n864_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT117), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n865_), .B(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n851_), .A2(G127gat), .A3(new_n644_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n870_), .A2(KEYINPUT118), .A3(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n868_), .A2(new_n872_), .ZN(G1342gat));
  OAI21_X1  g672(.A(new_n281_), .B1(new_n843_), .B2(new_n705_), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n874_), .A2(KEYINPUT119), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(KEYINPUT119), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n626_), .A2(new_n281_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(KEYINPUT120), .ZN(new_n878_));
  AOI22_X1  g677(.A1(new_n875_), .A2(new_n876_), .B1(new_n851_), .B2(new_n878_), .ZN(G1343gat));
  AND2_X1   g678(.A1(new_n837_), .A2(new_n302_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n661_), .A2(new_n397_), .A3(new_n657_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n235_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(new_n309_), .ZN(G1344gat));
  NOR2_X1   g683(.A1(new_n882_), .A2(new_n596_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(new_n310_), .ZN(G1345gat));
  NOR2_X1   g685(.A1(new_n882_), .A2(new_n645_), .ZN(new_n887_));
  XOR2_X1   g686(.A(KEYINPUT61), .B(G155gat), .Z(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1346gat));
  OAI21_X1  g688(.A(G162gat), .B1(new_n882_), .B2(new_n626_), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n705_), .A2(G162gat), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n882_), .B2(new_n891_), .ZN(G1347gat));
  AND3_X1   g691(.A1(new_n661_), .A2(new_n397_), .A3(new_n511_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n837_), .A2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n234_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(KEYINPUT62), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n263_), .B1(new_n896_), .B2(KEYINPUT62), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n895_), .A2(new_n897_), .A3(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n897_), .B1(new_n895_), .B2(new_n898_), .ZN(new_n900_));
  XOR2_X1   g699(.A(KEYINPUT22), .B(G169gat), .Z(new_n901_));
  OAI22_X1  g700(.A1(new_n899_), .A2(new_n900_), .B1(new_n895_), .B2(new_n901_), .ZN(G1348gat));
  NAND2_X1  g701(.A1(new_n894_), .A2(new_n704_), .ZN(new_n903_));
  XOR2_X1   g702(.A(KEYINPUT122), .B(G176gat), .Z(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1349gat));
  NAND2_X1  g704(.A1(new_n894_), .A2(new_n644_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n906_), .A2(new_n246_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n907_), .B1(new_n242_), .B2(new_n906_), .ZN(G1350gat));
  INV_X1    g707(.A(new_n894_), .ZN(new_n909_));
  OAI21_X1  g708(.A(G190gat), .B1(new_n909_), .B2(new_n626_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n651_), .A2(new_n237_), .A3(new_n239_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n909_), .B2(new_n911_), .ZN(G1351gat));
  XOR2_X1   g711(.A(KEYINPUT124), .B(G197gat), .Z(new_n913_));
  INV_X1    g712(.A(new_n508_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n880_), .A2(new_n914_), .A3(new_n661_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT123), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n880_), .A2(KEYINPUT123), .A3(new_n914_), .A4(new_n661_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n913_), .B1(new_n919_), .B2(new_n234_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(KEYINPUT124), .A2(G197gat), .ZN(new_n921_));
  AOI211_X1 g720(.A(new_n235_), .B(new_n921_), .C1(new_n917_), .C2(new_n918_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n920_), .A2(new_n922_), .ZN(G1352gat));
  AOI21_X1  g722(.A(new_n596_), .B1(new_n917_), .B2(new_n918_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n925_));
  XOR2_X1   g724(.A(new_n925_), .B(KEYINPUT126), .Z(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n924_), .B(new_n927_), .ZN(G1353gat));
  OR2_X1    g727(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n929_), .B1(new_n919_), .B2(new_n644_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(KEYINPUT63), .B(G211gat), .ZN(new_n931_));
  AOI211_X1 g730(.A(new_n645_), .B(new_n931_), .C1(new_n917_), .C2(new_n918_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n930_), .A2(new_n932_), .ZN(G1354gat));
  NAND3_X1  g732(.A1(new_n919_), .A2(new_n342_), .A3(new_n651_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n626_), .B1(new_n917_), .B2(new_n918_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n342_), .B2(new_n935_), .ZN(G1355gat));
endmodule


