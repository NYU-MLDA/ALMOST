//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 1 0 1 0 0 1 0 0 0 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n861_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n899_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_;
  XNOR2_X1  g000(.A(G22gat), .B(G50gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G78gat), .B(G106gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT88), .ZN(new_n206_));
  INV_X1    g005(.A(G155gat), .ZN(new_n207_));
  INV_X1    g006(.A(G162gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT1), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(G155gat), .A3(G162gat), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n209_), .B(new_n211_), .C1(G155gat), .C2(G162gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G141gat), .A2(G148gat), .ZN(new_n213_));
  INV_X1    g012(.A(G141gat), .ZN(new_n214_));
  INV_X1    g013(.A(G148gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n212_), .A2(new_n213_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n214_), .A2(new_n215_), .A3(KEYINPUT3), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT3), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n220_), .B1(G141gat), .B2(G148gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT2), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT82), .B1(new_n213_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n213_), .A2(new_n223_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT82), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n226_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n222_), .A2(new_n224_), .A3(new_n225_), .A4(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(G155gat), .B(G162gat), .Z(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT83), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n228_), .A2(KEYINPUT83), .A3(new_n229_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n218_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT29), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n206_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT21), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT85), .ZN(new_n238_));
  INV_X1    g037(.A(G204gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(new_n239_), .A3(G197gat), .ZN(new_n240_));
  INV_X1    g039(.A(G197gat), .ZN(new_n241_));
  AOI21_X1  g040(.A(KEYINPUT85), .B1(new_n241_), .B2(G204gat), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(G204gat), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n237_), .B(new_n240_), .C1(new_n242_), .C2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT86), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n239_), .A2(G197gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n239_), .A2(G197gat), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n247_), .B1(new_n248_), .B2(KEYINPUT85), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n249_), .A2(KEYINPUT86), .A3(new_n237_), .A4(new_n240_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n241_), .A2(G204gat), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n237_), .B1(new_n247_), .B2(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(G211gat), .B(G218gat), .Z(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n246_), .A2(new_n250_), .A3(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT89), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n249_), .A2(new_n240_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(KEYINPUT21), .A3(new_n253_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n255_), .A2(new_n256_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n256_), .B1(new_n255_), .B2(new_n258_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  AND3_X1   g061(.A1(new_n228_), .A2(KEYINPUT83), .A3(new_n229_), .ZN(new_n263_));
  AOI21_X1  g062(.A(KEYINPUT83), .B1(new_n228_), .B2(new_n229_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n217_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(KEYINPUT88), .A3(KEYINPUT29), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n236_), .A2(new_n262_), .A3(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT84), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(G233gat), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n268_), .A2(G233gat), .ZN(new_n271_));
  OAI21_X1  g070(.A(G228gat), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n267_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n255_), .A2(new_n258_), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n275_), .B(new_n272_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT87), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n273_), .B1(new_n265_), .B2(KEYINPUT29), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT87), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(new_n279_), .A3(new_n275_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n277_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n234_), .A2(new_n235_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT28), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  AND3_X1   g083(.A1(new_n274_), .A2(new_n281_), .A3(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n284_), .B1(new_n274_), .B2(new_n281_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n205_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n274_), .A2(new_n281_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n284_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n274_), .A2(new_n281_), .A3(new_n284_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n290_), .A2(new_n291_), .A3(new_n204_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n287_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G8gat), .B(G36gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT18), .ZN(new_n295_));
  INV_X1    g094(.A(G64gat), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n296_), .ZN(new_n298_));
  AND3_X1   g097(.A1(new_n297_), .A2(G92gat), .A3(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(G92gat), .B1(new_n297_), .B2(new_n298_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n301_), .A2(KEYINPUT32), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT90), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT25), .B(G183gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT26), .B(G190gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G183gat), .A2(G190gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT23), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  OR2_X1    g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n312_), .A2(KEYINPUT24), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n312_), .A2(KEYINPUT24), .A3(new_n314_), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n306_), .A2(new_n311_), .A3(new_n313_), .A4(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(G169gat), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n309_), .B(new_n310_), .C1(G183gat), .C2(G190gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n316_), .A2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n303_), .B1(new_n275_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT20), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT78), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT26), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n324_), .B1(new_n325_), .B2(G190gat), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n304_), .B(new_n326_), .C1(new_n305_), .C2(new_n324_), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n327_), .A2(new_n311_), .A3(new_n313_), .A4(new_n315_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(new_n320_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n323_), .B1(new_n275_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G226gat), .A2(G233gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT19), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n316_), .A2(new_n320_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n334_), .A2(KEYINPUT90), .A3(new_n255_), .A4(new_n258_), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n322_), .A2(new_n330_), .A3(new_n333_), .A4(new_n335_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n255_), .A2(new_n320_), .A3(new_n328_), .A4(new_n258_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT20), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n334_), .B1(new_n255_), .B2(new_n258_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n332_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n336_), .A2(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n302_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n275_), .A2(new_n321_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n343_), .A2(KEYINPUT20), .A3(new_n333_), .A4(new_n337_), .ZN(new_n344_));
  OR2_X1    g143(.A1(new_n344_), .A2(KEYINPUT95), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(KEYINPUT95), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT94), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n334_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(new_n330_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n348_), .B1(new_n350_), .B2(new_n332_), .ZN(new_n351_));
  AOI211_X1 g150(.A(KEYINPUT94), .B(new_n333_), .C1(new_n349_), .C2(new_n330_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n347_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G127gat), .B(G134gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G113gat), .B(G120gat), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n354_), .B(new_n355_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n358_), .B1(new_n359_), .B2(new_n357_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT91), .B1(new_n234_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G225gat), .A2(G233gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n234_), .A2(new_n359_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT91), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n265_), .A2(new_n365_), .A3(new_n360_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n362_), .A2(new_n363_), .A3(new_n364_), .A4(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT93), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n367_), .A2(new_n368_), .ZN(new_n370_));
  AOI21_X1  g169(.A(KEYINPUT4), .B1(new_n265_), .B2(new_n360_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n362_), .A2(new_n364_), .A3(new_n366_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n371_), .B1(new_n372_), .B2(KEYINPUT4), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n363_), .B(KEYINPUT92), .ZN(new_n374_));
  OAI22_X1  g173(.A1(new_n369_), .A2(new_n370_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G1gat), .B(G29gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(G85gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT0), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(G57gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n375_), .A2(new_n379_), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n265_), .A2(new_n365_), .A3(new_n360_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n365_), .B1(new_n265_), .B2(new_n360_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n383_), .A2(KEYINPUT93), .A3(new_n363_), .A4(new_n364_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n367_), .A2(new_n368_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n379_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n386_), .B(new_n387_), .C1(new_n374_), .C2(new_n373_), .ZN(new_n388_));
  AOI221_X4 g187(.A(new_n342_), .B1(new_n353_), .B2(new_n302_), .C1(new_n380_), .C2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT33), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n390_), .B1(new_n375_), .B2(new_n379_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n374_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n383_), .A2(new_n392_), .A3(new_n364_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n363_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n379_), .B(new_n393_), .C1(new_n373_), .C2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n301_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n341_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n336_), .A2(new_n340_), .A3(new_n301_), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  AND2_X1   g198(.A1(new_n395_), .A2(new_n399_), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n373_), .A2(new_n374_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n401_), .A2(KEYINPUT33), .A3(new_n387_), .A4(new_n386_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n391_), .A2(new_n400_), .A3(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n293_), .B1(new_n389_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT27), .ZN(new_n405_));
  AND3_X1   g204(.A1(new_n397_), .A2(new_n405_), .A3(new_n398_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT96), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n398_), .A2(new_n407_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n336_), .A2(new_n340_), .A3(new_n301_), .A4(KEYINPUT96), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n275_), .A2(KEYINPUT89), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n321_), .B1(new_n410_), .B2(new_n259_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n330_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n332_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT94), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n350_), .A2(new_n348_), .A3(new_n332_), .ZN(new_n415_));
  AOI22_X1  g214(.A1(new_n414_), .A2(new_n415_), .B1(new_n346_), .B2(new_n345_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n408_), .B(new_n409_), .C1(new_n416_), .C2(new_n301_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n406_), .B1(new_n417_), .B2(KEYINPUT27), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n380_), .A2(new_n287_), .A3(new_n292_), .A4(new_n388_), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT97), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n406_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n408_), .A2(new_n409_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n422_), .B1(new_n396_), .B2(new_n353_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n421_), .B1(new_n423_), .B2(new_n405_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n287_), .A2(new_n292_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n380_), .A2(new_n388_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT97), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .A4(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n404_), .A2(new_n420_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(G43gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n329_), .B(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G71gat), .B(G99gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT30), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G227gat), .A2(G233gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(G15gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n433_), .B(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n431_), .B(new_n436_), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n437_), .A2(KEYINPUT80), .ZN(new_n438_));
  XOR2_X1   g237(.A(new_n360_), .B(KEYINPUT31), .Z(new_n439_));
  OR2_X1    g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n437_), .A2(KEYINPUT80), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n439_), .B1(new_n438_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  XOR2_X1   g242(.A(new_n443_), .B(KEYINPUT81), .Z(new_n444_));
  INV_X1    g243(.A(new_n443_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT98), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n446_), .B1(new_n418_), .B2(new_n425_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n424_), .A2(KEYINPUT98), .A3(new_n293_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n445_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  AOI22_X1  g248(.A1(new_n429_), .A2(new_n444_), .B1(new_n449_), .B2(new_n426_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT69), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G85gat), .B(G92gat), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT8), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(G99gat), .ZN(new_n457_));
  INV_X1    g256(.A(G106gat), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT7), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n457_), .A2(new_n458_), .B1(new_n459_), .B2(KEYINPUT66), .ZN(new_n460_));
  NOR2_X1   g259(.A1(G99gat), .A2(G106gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(KEYINPUT66), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT66), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT7), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n460_), .B1(new_n461_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G99gat), .A2(G106gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT6), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT6), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n469_), .A2(G99gat), .A3(G106gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n456_), .B1(new_n466_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT67), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n469_), .B1(G99gat), .B2(G106gat), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n467_), .A2(KEYINPUT6), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n473_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n465_), .A2(new_n461_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n460_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n468_), .A2(new_n470_), .A3(KEYINPUT67), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .A4(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n454_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n472_), .B1(new_n481_), .B2(KEYINPUT8), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT9), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n453_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(G85gat), .A3(G92gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n471_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT10), .B(G99gat), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT65), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  AOI211_X1 g288(.A(new_n484_), .B(new_n486_), .C1(new_n489_), .C2(new_n458_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n452_), .B(KEYINPUT12), .C1(new_n482_), .C2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n466_), .A2(new_n471_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n492_), .A2(new_n455_), .A3(new_n454_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n468_), .A2(new_n470_), .A3(KEYINPUT67), .ZN(new_n494_));
  AOI21_X1  g293(.A(KEYINPUT67), .B1(new_n468_), .B2(new_n470_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n453_), .B1(new_n496_), .B2(new_n466_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n493_), .B1(new_n497_), .B2(new_n455_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT12), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n486_), .B1(new_n489_), .B2(new_n458_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n454_), .A2(KEYINPUT9), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n498_), .A2(new_n499_), .A3(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n491_), .A2(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(G57gat), .B(G64gat), .Z(new_n505_));
  INV_X1    g304(.A(KEYINPUT11), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  AOI22_X1  g307(.A1(new_n505_), .A2(new_n506_), .B1(G71gat), .B2(G78gat), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT68), .ZN(new_n510_));
  INV_X1    g309(.A(G71gat), .ZN(new_n511_));
  INV_X1    g310(.A(G78gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n509_), .A2(new_n510_), .A3(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n510_), .B1(new_n509_), .B2(new_n513_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n508_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n505_), .A2(new_n506_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G71gat), .A2(G78gat), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(new_n513_), .A3(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT68), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n509_), .A2(new_n510_), .A3(new_n513_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n521_), .A3(new_n507_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n516_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n504_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G230gat), .A2(G233gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT64), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n516_), .A2(new_n522_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(new_n491_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n524_), .A2(new_n527_), .A3(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(G120gat), .B(G148gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(G176gat), .B(G204gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n482_), .A2(new_n490_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(new_n528_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n523_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n538_), .A2(new_n526_), .A3(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n530_), .A2(new_n535_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n535_), .B(KEYINPUT71), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n543_), .B1(new_n530_), .B2(new_n540_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(KEYINPUT72), .B(KEYINPUT13), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT72), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n545_), .B1(new_n548_), .B2(KEYINPUT13), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G229gat), .A2(G233gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G29gat), .B(G36gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(new_n430_), .ZN(new_n554_));
  INV_X1    g353(.A(G50gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G15gat), .B(G22gat), .ZN(new_n557_));
  INV_X1    g356(.A(G1gat), .ZN(new_n558_));
  INV_X1    g357(.A(G8gat), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT14), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n557_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G1gat), .B(G8gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n556_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT15), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n556_), .B(new_n566_), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n552_), .B(new_n565_), .C1(new_n567_), .C2(new_n564_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n556_), .B(new_n564_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n569_), .A2(G229gat), .A3(G233gat), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G113gat), .B(G141gat), .ZN(new_n572_));
  INV_X1    g371(.A(G169gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(new_n241_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n571_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n575_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n568_), .A2(new_n570_), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n551_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n451_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n563_), .B(new_n583_), .Z(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(new_n523_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G127gat), .B(G155gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G183gat), .B(G211gat), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n588_), .B(new_n589_), .Z(new_n590_));
  AND3_X1   g389(.A1(new_n590_), .A2(new_n452_), .A3(KEYINPUT17), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n585_), .A2(new_n592_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n585_), .B(new_n592_), .C1(KEYINPUT17), .C2(new_n590_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n556_), .B(KEYINPUT15), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(new_n537_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n536_), .A2(new_n556_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G232gat), .A2(G233gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT34), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT35), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n599_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT73), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT73), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n599_), .A2(new_n607_), .A3(new_n604_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G190gat), .B(G218gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT74), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(G134gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(new_n208_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n613_), .A2(KEYINPUT36), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n599_), .B1(new_n603_), .B2(new_n602_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n604_), .B(KEYINPUT75), .Z(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n609_), .A2(new_n614_), .A3(new_n617_), .ZN(new_n618_));
  AOI22_X1  g417(.A1(new_n606_), .A2(new_n608_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n613_), .B(KEYINPUT36), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n618_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT76), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n622_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n621_), .A2(new_n623_), .A3(KEYINPUT37), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT37), .ZN(new_n625_));
  OAI221_X1 g424(.A(new_n618_), .B1(new_n622_), .B2(new_n625_), .C1(new_n619_), .C2(new_n620_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n595_), .B1(new_n624_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n582_), .A2(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n426_), .B(KEYINPUT99), .Z(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(new_n558_), .A3(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n632_));
  XOR2_X1   g431(.A(new_n631_), .B(new_n632_), .Z(new_n633_));
  INV_X1    g432(.A(new_n621_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n582_), .A2(new_n634_), .A3(new_n595_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n426_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n558_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n633_), .A2(new_n637_), .ZN(G1324gat));
  AOI21_X1  g437(.A(new_n559_), .B1(new_n635_), .B2(new_n418_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT39), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n629_), .A2(new_n559_), .A3(new_n418_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT101), .Z(new_n642_));
  NOR2_X1   g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT40), .ZN(G1325gat));
  INV_X1    g443(.A(G15gat), .ZN(new_n645_));
  INV_X1    g444(.A(new_n444_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n635_), .B2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT41), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n629_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(G1326gat));
  INV_X1    g449(.A(G22gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n293_), .B(KEYINPUT102), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n651_), .B1(new_n635_), .B2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT103), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT42), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n629_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1327gat));
  NAND2_X1  g456(.A1(new_n634_), .A2(new_n595_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n582_), .A2(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(G29gat), .B1(new_n659_), .B2(new_n636_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n630_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n624_), .A2(new_n626_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n420_), .A2(new_n428_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n353_), .A2(new_n302_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n342_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n380_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n388_), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n665_), .B(new_n666_), .C1(new_n667_), .C2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n391_), .A2(new_n400_), .A3(new_n402_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n425_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n444_), .B1(new_n664_), .B2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n447_), .A2(new_n448_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n673_), .A2(new_n426_), .A3(new_n443_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n663_), .B1(new_n672_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n662_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  OAI211_X1 g476(.A(KEYINPUT104), .B(KEYINPUT43), .C1(new_n450_), .C2(new_n663_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n675_), .A2(new_n676_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n677_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT105), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT44), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n581_), .B1(new_n681_), .B2(KEYINPUT44), .ZN(new_n683_));
  INV_X1    g482(.A(new_n595_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n680_), .A2(new_n682_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n682_), .B1(new_n680_), .B2(new_n685_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n661_), .B1(new_n687_), .B2(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n660_), .B1(new_n690_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g490(.A(new_n659_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n692_), .A2(G36gat), .A3(new_n424_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n418_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n696_), .A2(KEYINPUT106), .A3(G36gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT106), .B1(new_n696_), .B2(G36gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n695_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT46), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  OAI211_X1 g500(.A(KEYINPUT46), .B(new_n695_), .C1(new_n697_), .C2(new_n698_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1329gat));
  NOR3_X1   g502(.A1(new_n692_), .A2(G43gat), .A3(new_n444_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n443_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(G43gat), .ZN(new_n706_));
  XNOR2_X1  g505(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n706_), .B(new_n707_), .ZN(G1330gat));
  NAND3_X1  g507(.A1(new_n659_), .A2(new_n555_), .A3(new_n652_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n293_), .B1(new_n687_), .B2(new_n689_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(new_n710_), .B2(new_n555_), .ZN(G1331gat));
  NOR2_X1   g510(.A1(new_n550_), .A2(new_n579_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n451_), .A2(new_n712_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n713_), .A2(new_n628_), .ZN(new_n714_));
  AOI21_X1  g513(.A(G57gat), .B1(new_n714_), .B2(new_n630_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n713_), .A2(new_n634_), .A3(new_n595_), .ZN(new_n716_));
  XOR2_X1   g515(.A(KEYINPUT109), .B(G57gat), .Z(new_n717_));
  NOR2_X1   g516(.A1(new_n426_), .A2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n715_), .B1(new_n716_), .B2(new_n718_), .ZN(G1332gat));
  AOI21_X1  g518(.A(new_n296_), .B1(new_n716_), .B2(new_n418_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT48), .Z(new_n721_));
  NAND3_X1  g520(.A1(new_n714_), .A2(new_n296_), .A3(new_n418_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1333gat));
  AOI21_X1  g522(.A(new_n511_), .B1(new_n716_), .B2(new_n646_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT49), .Z(new_n725_));
  NAND3_X1  g524(.A1(new_n714_), .A2(new_n511_), .A3(new_n646_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1334gat));
  AOI21_X1  g526(.A(new_n512_), .B1(new_n716_), .B2(new_n652_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT110), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT50), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n714_), .A2(new_n512_), .A3(new_n652_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1335gat));
  NAND3_X1  g531(.A1(new_n680_), .A2(new_n595_), .A3(new_n712_), .ZN(new_n733_));
  OAI21_X1  g532(.A(G85gat), .B1(new_n733_), .B2(new_n426_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n713_), .A2(new_n658_), .ZN(new_n735_));
  INV_X1    g534(.A(G85gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(new_n736_), .A3(new_n630_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n734_), .A2(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT111), .ZN(G1336gat));
  AOI21_X1  g538(.A(G92gat), .B1(new_n735_), .B2(new_n418_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n733_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n418_), .A2(G92gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n740_), .B1(new_n741_), .B2(new_n742_), .ZN(G1337gat));
  OAI21_X1  g542(.A(G99gat), .B1(new_n733_), .B2(new_n444_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n735_), .A2(new_n489_), .A3(new_n443_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n746_), .A2(KEYINPUT112), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(KEYINPUT112), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n747_), .A2(KEYINPUT51), .A3(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(KEYINPUT51), .B1(new_n747_), .B2(new_n748_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1338gat));
  NAND3_X1  g550(.A1(new_n735_), .A2(new_n458_), .A3(new_n425_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n680_), .A2(new_n425_), .A3(new_n595_), .A4(new_n712_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n753_), .A2(G106gat), .A3(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n753_), .B2(G106gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n752_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g557(.A1(new_n449_), .A2(new_n630_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n543_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n528_), .B1(new_n491_), .B2(new_n503_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n499_), .B1(new_n498_), .B2(new_n502_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n523_), .B1(new_n762_), .B2(new_n452_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n761_), .A2(new_n763_), .A3(new_n526_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n526_), .B1(new_n761_), .B2(new_n763_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(KEYINPUT55), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT55), .ZN(new_n767_));
  NOR4_X1   g566(.A1(new_n761_), .A2(new_n763_), .A3(new_n767_), .A4(new_n526_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n760_), .B1(new_n766_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT56), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n527_), .B1(new_n524_), .B2(new_n529_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n530_), .B1(new_n772_), .B2(new_n767_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n768_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(KEYINPUT56), .A3(new_n760_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n771_), .A2(KEYINPUT115), .A3(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n579_), .A2(new_n541_), .ZN(new_n778_));
  AOI211_X1 g577(.A(new_n770_), .B(new_n543_), .C1(new_n773_), .C2(new_n774_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT115), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n778_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n777_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n569_), .A2(new_n552_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n565_), .B1(new_n567_), .B2(new_n564_), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n783_), .B(new_n575_), .C1(new_n784_), .C2(new_n552_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n785_), .A2(new_n578_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n786_), .B1(new_n542_), .B2(new_n544_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT116), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT116), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n786_), .B(new_n789_), .C1(new_n542_), .C2(new_n544_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n634_), .B1(new_n782_), .B2(new_n792_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT118), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT118), .ZN(new_n796_));
  INV_X1    g595(.A(new_n794_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n791_), .B1(new_n777_), .B2(new_n781_), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n796_), .B(new_n797_), .C1(new_n798_), .C2(new_n634_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n795_), .A2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT56), .B1(new_n775_), .B2(new_n760_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n541_), .B(new_n786_), .C1(new_n801_), .C2(new_n779_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT58), .ZN(new_n803_));
  INV_X1    g602(.A(new_n663_), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n803_), .A2(new_n804_), .B1(new_n793_), .B2(KEYINPUT57), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n800_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT119), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT119), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n800_), .A2(new_n808_), .A3(new_n805_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n807_), .A2(new_n595_), .A3(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n627_), .A2(new_n811_), .A3(new_n580_), .A4(new_n550_), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n812_), .A2(KEYINPUT114), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n627_), .A2(new_n580_), .A3(new_n550_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT54), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n812_), .A2(KEYINPUT114), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n813_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n759_), .B1(new_n810_), .B2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(G113gat), .B1(new_n818_), .B2(new_n579_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT59), .ZN(new_n820_));
  OR2_X1    g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n803_), .A2(new_n804_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n793_), .A2(KEYINPUT57), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n797_), .B1(new_n798_), .B2(new_n634_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n822_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n595_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT120), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n825_), .A2(KEYINPUT120), .A3(new_n595_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n817_), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n759_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n830_), .A2(new_n820_), .A3(new_n831_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n821_), .A2(new_n832_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n579_), .A2(G113gat), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n819_), .B1(new_n833_), .B2(new_n834_), .ZN(G1340gat));
  OAI211_X1 g634(.A(new_n551_), .B(new_n832_), .C1(new_n818_), .C2(new_n820_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(G120gat), .ZN(new_n837_));
  INV_X1    g636(.A(G120gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n550_), .B2(KEYINPUT60), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n818_), .B(new_n839_), .C1(KEYINPUT60), .C2(new_n838_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n837_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT121), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n837_), .A2(KEYINPUT121), .A3(new_n840_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(G1341gat));
  AOI21_X1  g644(.A(G127gat), .B1(new_n818_), .B2(new_n684_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n684_), .A2(G127gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n833_), .B2(new_n847_), .ZN(G1342gat));
  AOI21_X1  g647(.A(G134gat), .B1(new_n818_), .B2(new_n634_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n804_), .A2(G134gat), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n849_), .B1(new_n833_), .B2(new_n850_), .ZN(G1343gat));
  INV_X1    g650(.A(KEYINPUT122), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n810_), .A2(new_n817_), .ZN(new_n853_));
  NOR4_X1   g652(.A1(new_n661_), .A2(new_n646_), .A3(new_n418_), .A4(new_n293_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n852_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n854_), .ZN(new_n856_));
  AOI211_X1 g655(.A(KEYINPUT122), .B(new_n856_), .C1(new_n810_), .C2(new_n817_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n579_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(KEYINPUT123), .B(G141gat), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1344gat));
  OAI21_X1  g659(.A(new_n551_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(G148gat), .ZN(G1345gat));
  OAI21_X1  g661(.A(new_n684_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(KEYINPUT61), .B(G155gat), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n863_), .B(new_n864_), .ZN(G1346gat));
  OAI211_X1 g664(.A(G162gat), .B(new_n804_), .C1(new_n855_), .C2(new_n857_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  AND3_X1   g666(.A1(new_n800_), .A2(new_n808_), .A3(new_n805_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n808_), .B1(new_n800_), .B2(new_n805_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n868_), .A2(new_n869_), .A3(new_n684_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n817_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n854_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(KEYINPUT122), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n853_), .A2(new_n852_), .A3(new_n854_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n621_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(KEYINPUT124), .B1(new_n875_), .B2(G162gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n634_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT124), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n877_), .A2(new_n878_), .A3(new_n208_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n867_), .B1(new_n876_), .B2(new_n879_), .ZN(G1347gat));
  INV_X1    g679(.A(new_n652_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n661_), .A2(new_n646_), .A3(new_n418_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n830_), .A2(new_n579_), .A3(new_n881_), .A4(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(G169gat), .B1(new_n884_), .B2(KEYINPUT62), .ZN(new_n885_));
  OAI21_X1  g684(.A(KEYINPUT62), .B1(new_n884_), .B2(KEYINPUT22), .ZN(new_n886_));
  MUX2_X1   g685(.A(G169gat), .B(new_n885_), .S(new_n886_), .Z(G1348gat));
  NAND3_X1  g686(.A1(new_n830_), .A2(new_n881_), .A3(new_n883_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(G176gat), .B1(new_n889_), .B2(new_n551_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n425_), .B1(new_n810_), .B2(new_n817_), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n891_), .A2(G176gat), .A3(new_n883_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n890_), .B1(new_n551_), .B2(new_n892_), .ZN(G1349gat));
  NOR3_X1   g692(.A1(new_n888_), .A2(new_n304_), .A3(new_n595_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n891_), .A2(new_n684_), .A3(new_n883_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(KEYINPUT125), .ZN(new_n896_));
  INV_X1    g695(.A(G183gat), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n894_), .B1(new_n896_), .B2(new_n897_), .ZN(G1350gat));
  OAI21_X1  g697(.A(G190gat), .B1(new_n888_), .B2(new_n663_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n634_), .A2(new_n305_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(KEYINPUT126), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n899_), .B1(new_n888_), .B2(new_n901_), .ZN(G1351gat));
  AOI21_X1  g701(.A(new_n424_), .B1(new_n810_), .B2(new_n817_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n646_), .A2(new_n419_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n905_), .A2(new_n580_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT127), .B(G197gat), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n906_), .B(new_n907_), .ZN(G1352gat));
  NOR2_X1   g707(.A1(new_n905_), .A2(new_n550_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(new_n239_), .ZN(G1353gat));
  NOR2_X1   g709(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n911_));
  AND2_X1   g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  NOR4_X1   g711(.A1(new_n905_), .A2(new_n595_), .A3(new_n911_), .A4(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n905_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(new_n684_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n913_), .B1(new_n915_), .B2(new_n911_), .ZN(G1354gat));
  AND3_X1   g715(.A1(new_n914_), .A2(G218gat), .A3(new_n804_), .ZN(new_n917_));
  AOI21_X1  g716(.A(G218gat), .B1(new_n914_), .B2(new_n634_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1355gat));
endmodule


