//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n642_,
    new_n643_, new_n644_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n853_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n895_, new_n897_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_;
  XNOR2_X1  g000(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT23), .ZN(new_n207_));
  INV_X1    g006(.A(G169gat), .ZN(new_n208_));
  INV_X1    g007(.A(G176gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n210_), .A2(KEYINPUT24), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(KEYINPUT24), .A3(new_n212_), .ZN(new_n213_));
  AND3_X1   g012(.A1(new_n207_), .A2(new_n211_), .A3(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT25), .B(G183gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT94), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT26), .B(G190gat), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n214_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT22), .B(G169gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(new_n209_), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n222_), .A2(new_n212_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n207_), .B1(G183gat), .B2(G190gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n220_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT88), .B(G197gat), .ZN(new_n227_));
  MUX2_X1   g026(.A(G197gat), .B(new_n227_), .S(G204gat), .Z(new_n228_));
  INV_X1    g027(.A(KEYINPUT21), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G211gat), .B(G218gat), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n229_), .B1(new_n230_), .B2(KEYINPUT90), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n228_), .B(new_n231_), .C1(KEYINPUT90), .C2(new_n230_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n230_), .ZN(new_n233_));
  INV_X1    g032(.A(G204gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n227_), .A2(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n229_), .B1(G197gat), .B2(G204gat), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n233_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT89), .B(KEYINPUT21), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n237_), .B1(new_n228_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n232_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n226_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT20), .ZN(new_n242_));
  NOR2_X1   g041(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT80), .B(G183gat), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n243_), .B1(new_n244_), .B2(KEYINPUT25), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n214_), .B1(new_n219_), .B2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n207_), .B1(G190gat), .B2(new_n244_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n222_), .A2(KEYINPUT81), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT81), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n221_), .A2(new_n249_), .A3(new_n209_), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n247_), .A2(new_n248_), .A3(new_n212_), .A4(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n246_), .A2(new_n251_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n252_), .A2(new_n240_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n205_), .B1(new_n242_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT20), .ZN(new_n255_));
  AND2_X1   g054(.A1(new_n220_), .A2(new_n225_), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n232_), .A2(new_n239_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n255_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n252_), .A2(new_n240_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(new_n204_), .A3(new_n259_), .ZN(new_n260_));
  XOR2_X1   g059(.A(G8gat), .B(G36gat), .Z(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G64gat), .B(G92gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n254_), .A2(new_n260_), .A3(new_n265_), .ZN(new_n266_));
  NOR3_X1   g065(.A1(new_n242_), .A2(new_n205_), .A3(new_n253_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n204_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n265_), .B(KEYINPUT98), .ZN(new_n270_));
  OAI211_X1 g069(.A(KEYINPUT27), .B(new_n266_), .C1(new_n269_), .C2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT27), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT20), .B1(new_n226_), .B2(new_n240_), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n252_), .A2(new_n240_), .ZN(new_n274_));
  NOR3_X1   g073(.A1(new_n273_), .A2(new_n274_), .A3(new_n205_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n257_), .A2(new_n246_), .A3(new_n251_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n255_), .B1(new_n226_), .B2(new_n240_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n204_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n265_), .ZN(new_n279_));
  NOR3_X1   g078(.A1(new_n275_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n265_), .B1(new_n254_), .B2(new_n260_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n272_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n271_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G141gat), .A2(G148gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT2), .ZN(new_n285_));
  NOR2_X1   g084(.A1(G141gat), .A2(G148gat), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT84), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n287_), .B1(new_n288_), .B2(KEYINPUT3), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT3), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n286_), .A2(KEYINPUT84), .A3(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n285_), .A2(new_n289_), .A3(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT85), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT85), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n285_), .A2(new_n289_), .A3(new_n294_), .A4(new_n291_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n296_), .A2(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(G127gat), .B(G134gat), .Z(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT82), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G127gat), .B(G134gat), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT82), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G113gat), .B(G120gat), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n304_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n308_), .B1(new_n304_), .B2(new_n307_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n299_), .B1(KEYINPUT1), .B2(new_n297_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n313_), .B1(KEYINPUT1), .B2(new_n297_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(new_n284_), .A3(new_n287_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n302_), .A2(new_n312_), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n311_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n309_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n300_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n315_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n318_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n316_), .A2(KEYINPUT4), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT96), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT96), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n316_), .A2(new_n321_), .A3(new_n324_), .A4(KEYINPUT4), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT4), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n327_), .B(new_n318_), .C1(new_n319_), .C2(new_n320_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G225gat), .A2(G233gat), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n326_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n316_), .A2(new_n321_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n334_), .A2(new_n330_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G1gat), .B(G29gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(G85gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT0), .B(G57gat), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n338_), .B(new_n339_), .Z(new_n340_));
  NAND3_X1  g139(.A1(new_n333_), .A2(new_n336_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT83), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n318_), .A2(KEYINPUT31), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT31), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n344_), .B1(new_n317_), .B2(new_n309_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G227gat), .A2(G233gat), .ZN(new_n347_));
  XOR2_X1   g146(.A(new_n347_), .B(G15gat), .Z(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT30), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G71gat), .B(G99gat), .ZN(new_n351_));
  INV_X1    g150(.A(G43gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n246_), .A2(new_n251_), .A3(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n354_), .B1(new_n246_), .B2(new_n251_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n350_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n252_), .A2(new_n353_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n246_), .A2(new_n251_), .A3(new_n354_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n358_), .A2(new_n349_), .A3(new_n359_), .ZN(new_n360_));
  AOI211_X1 g159(.A(new_n342_), .B(new_n346_), .C1(new_n357_), .C2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n357_), .A2(new_n360_), .A3(new_n342_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n362_), .A2(new_n346_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n357_), .A2(new_n360_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT83), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n361_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n340_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n331_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n367_), .B1(new_n368_), .B2(new_n335_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n341_), .A2(new_n366_), .A3(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n319_), .A2(new_n320_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n240_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G78gat), .B(G106gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT91), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n373_), .A2(new_n376_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n240_), .B(new_n375_), .C1(new_n371_), .C2(new_n372_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(G233gat), .ZN(new_n380_));
  NOR2_X1   g179(.A1(KEYINPUT87), .A2(G228gat), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(KEYINPUT87), .A2(G228gat), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n380_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n379_), .B(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT28), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n387_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n388_));
  NOR4_X1   g187(.A1(new_n319_), .A2(KEYINPUT28), .A3(new_n320_), .A4(KEYINPUT29), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT86), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n302_), .A2(new_n372_), .A3(new_n315_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT28), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT86), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n371_), .A2(new_n387_), .A3(new_n372_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n392_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  XOR2_X1   g194(.A(G22gat), .B(G50gat), .Z(new_n396_));
  NAND3_X1  g195(.A1(new_n390_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n390_), .A2(new_n395_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n396_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n386_), .A2(KEYINPUT92), .A3(new_n397_), .A4(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT92), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n390_), .A2(new_n396_), .A3(new_n395_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n396_), .B1(new_n390_), .B2(new_n395_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n402_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n400_), .A2(KEYINPUT92), .A3(new_n397_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n379_), .B(new_n384_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n405_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  AOI211_X1 g207(.A(new_n283_), .B(new_n370_), .C1(new_n401_), .C2(new_n408_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n271_), .A2(new_n341_), .A3(new_n282_), .A4(new_n369_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n410_), .A2(new_n408_), .A3(new_n401_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n366_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NOR3_X1   g212(.A1(new_n368_), .A2(new_n335_), .A3(new_n367_), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT33), .B1(new_n414_), .B2(KEYINPUT97), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT97), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT33), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n341_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n279_), .B1(new_n275_), .B2(new_n278_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n266_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n326_), .A2(new_n329_), .A3(new_n328_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n334_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n340_), .B1(new_n422_), .B2(new_n330_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n420_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n415_), .A2(new_n418_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n408_), .A2(new_n401_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n265_), .A2(KEYINPUT32), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n254_), .A2(new_n260_), .A3(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n340_), .B1(new_n333_), .B2(new_n336_), .ZN(new_n429_));
  OAI221_X1 g228(.A(new_n428_), .B1(new_n269_), .B2(new_n427_), .C1(new_n429_), .C2(new_n414_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n425_), .A2(new_n426_), .A3(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n409_), .B1(new_n413_), .B2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G15gat), .B(G22gat), .ZN(new_n433_));
  INV_X1    g232(.A(G1gat), .ZN(new_n434_));
  INV_X1    g233(.A(G8gat), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT14), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n433_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G1gat), .B(G8gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G29gat), .B(G36gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G43gat), .B(G50gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(new_n439_), .B(new_n442_), .Z(new_n443_));
  NAND2_X1  g242(.A1(G229gat), .A2(G233gat), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n442_), .B(KEYINPUT15), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n439_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n439_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(new_n442_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n446_), .B1(new_n451_), .B2(new_n445_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G113gat), .B(G141gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G169gat), .B(G197gat), .ZN(new_n454_));
  XOR2_X1   g253(.A(new_n453_), .B(new_n454_), .Z(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n452_), .A2(new_n456_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n446_), .B(new_n455_), .C1(new_n445_), .C2(new_n451_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n432_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G85gat), .B(G92gat), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT9), .ZN(new_n464_));
  XOR2_X1   g263(.A(KEYINPUT10), .B(G99gat), .Z(new_n465_));
  INV_X1    g264(.A(G106gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G99gat), .A2(G106gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT6), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT6), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n470_), .A2(G99gat), .A3(G106gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT9), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(G85gat), .A3(G92gat), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n464_), .A2(new_n467_), .A3(new_n472_), .A4(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT8), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NOR3_X1   g278(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n462_), .B1(new_n481_), .B2(new_n472_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT65), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n477_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT7), .ZN(new_n485_));
  INV_X1    g284(.A(G99gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n486_), .A3(new_n466_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n472_), .A2(new_n478_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n463_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT65), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n484_), .A2(new_n490_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n469_), .A2(new_n471_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n487_), .A2(new_n478_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT64), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT64), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n472_), .A2(new_n495_), .A3(new_n478_), .A4(new_n487_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n462_), .A2(KEYINPUT8), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n494_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n476_), .B1(new_n491_), .B2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT72), .B1(new_n499_), .B2(new_n442_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n483_), .B(new_n463_), .C1(new_n492_), .C2(new_n493_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT8), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n483_), .B1(new_n488_), .B2(new_n463_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n498_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n504_), .A2(KEYINPUT72), .A3(new_n442_), .A4(new_n475_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G232gat), .A2(G233gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT34), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n507_), .A2(KEYINPUT35), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n505_), .A2(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n500_), .A2(new_n509_), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n496_), .A2(new_n497_), .ZN(new_n511_));
  AOI22_X1  g310(.A1(new_n484_), .A2(new_n490_), .B1(new_n511_), .B2(new_n494_), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT67), .B1(new_n512_), .B2(new_n476_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT67), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n504_), .A2(new_n514_), .A3(new_n475_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n513_), .A2(new_n447_), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT71), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n507_), .A2(KEYINPUT35), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT70), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n510_), .B(new_n516_), .C1(new_n517_), .C2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n504_), .A2(new_n442_), .A3(new_n475_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT72), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n523_), .A2(new_n517_), .A3(new_n508_), .A4(new_n505_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n519_), .ZN(new_n525_));
  AND3_X1   g324(.A1(new_n513_), .A2(new_n447_), .A3(new_n515_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n523_), .A2(new_n508_), .A3(new_n505_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n524_), .B(new_n525_), .C1(new_n526_), .C2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n520_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT73), .ZN(new_n530_));
  XOR2_X1   g329(.A(G190gat), .B(G218gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(G134gat), .B(G162gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT36), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n529_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n533_), .A2(new_n534_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n530_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n537_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n529_), .B(KEYINPUT73), .C1(new_n539_), .C2(new_n535_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n538_), .A2(KEYINPUT37), .A3(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(KEYINPUT37), .B1(new_n538_), .B2(new_n540_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G231gat), .A2(G233gat), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n439_), .B(new_n544_), .Z(new_n545_));
  XOR2_X1   g344(.A(new_n545_), .B(KEYINPUT74), .Z(new_n546_));
  XNOR2_X1  g345(.A(G57gat), .B(G64gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT11), .ZN(new_n548_));
  XOR2_X1   g347(.A(G71gat), .B(G78gat), .Z(new_n549_));
  OR2_X1    g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n547_), .A2(KEYINPUT11), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n548_), .A2(new_n549_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n550_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n546_), .B(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(G183gat), .B(G211gat), .Z(new_n555_));
  XNOR2_X1  g354(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G127gat), .B(G155gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT17), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT78), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n554_), .A2(new_n563_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n561_), .A2(KEYINPUT17), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n553_), .A2(KEYINPUT66), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT66), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n550_), .B(new_n567_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(new_n545_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n565_), .A2(new_n571_), .A3(new_n562_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n564_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT79), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n543_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT12), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n553_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n513_), .A2(new_n515_), .A3(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n576_), .B1(new_n499_), .B2(new_n569_), .ZN(new_n580_));
  AND2_X1   g379(.A1(G230gat), .A2(G233gat), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n581_), .B1(new_n499_), .B2(new_n569_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n579_), .A2(new_n580_), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT68), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n499_), .A2(new_n569_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n499_), .A2(new_n569_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n581_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n579_), .A2(KEYINPUT68), .A3(new_n580_), .A4(new_n582_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n585_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G120gat), .B(G148gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT5), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G176gat), .B(G204gat), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n593_), .B(new_n594_), .Z(new_n595_));
  NAND2_X1  g394(.A1(new_n591_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n595_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n585_), .A2(new_n589_), .A3(new_n590_), .A4(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT13), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n600_), .A2(KEYINPUT69), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT69), .B(KEYINPUT13), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n603_), .B1(new_n596_), .B2(new_n598_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n461_), .A2(new_n575_), .A3(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT99), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n429_), .A2(new_n414_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n608_), .A2(new_n434_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT38), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n283_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n426_), .A2(new_n614_), .A3(new_n609_), .A4(new_n366_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n425_), .A2(new_n426_), .A3(new_n430_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n411_), .A2(new_n412_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n615_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n538_), .A2(new_n540_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT100), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n605_), .A2(new_n460_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n622_), .A2(new_n572_), .A3(new_n564_), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(G1gat), .B1(new_n624_), .B2(new_n609_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n611_), .A2(new_n612_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n626_), .A2(KEYINPUT101), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(KEYINPUT101), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n613_), .B(new_n625_), .C1(new_n627_), .C2(new_n628_), .ZN(G1324gat));
  OAI21_X1  g428(.A(G8gat), .B1(new_n624_), .B2(new_n614_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT39), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n608_), .A2(new_n435_), .A3(new_n283_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT40), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(G1325gat));
  OAI21_X1  g434(.A(G15gat), .B1(new_n624_), .B2(new_n412_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(KEYINPUT102), .B(KEYINPUT41), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n637_), .ZN(new_n639_));
  OR3_X1    g438(.A1(new_n607_), .A2(G15gat), .A3(new_n412_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n638_), .A2(new_n639_), .A3(new_n640_), .ZN(G1326gat));
  OAI21_X1  g440(.A(G22gat), .B1(new_n624_), .B2(new_n426_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT42), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n426_), .A2(G22gat), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n643_), .B1(new_n607_), .B2(new_n644_), .ZN(G1327gat));
  NAND2_X1  g444(.A1(new_n574_), .A2(new_n619_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n646_), .A2(new_n605_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(new_n461_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(G29gat), .B1(new_n649_), .B2(new_n610_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n541_), .A2(new_n542_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n651_), .B1(new_n432_), .B2(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n618_), .A2(KEYINPUT43), .A3(new_n543_), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n653_), .A2(new_n654_), .A3(new_n574_), .A4(new_n622_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT44), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n573_), .B(KEYINPUT79), .Z(new_n658_));
  NAND2_X1  g457(.A1(new_n618_), .A2(new_n543_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n659_), .B2(new_n651_), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n660_), .A2(KEYINPUT44), .A3(new_n622_), .A4(new_n654_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n657_), .A2(new_n661_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n610_), .A2(G29gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n650_), .B1(new_n662_), .B2(new_n663_), .ZN(G1328gat));
  NOR3_X1   g463(.A1(new_n648_), .A2(G36gat), .A3(new_n614_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT45), .Z(new_n666_));
  NAND3_X1  g465(.A1(new_n657_), .A2(new_n661_), .A3(new_n283_), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n667_), .A2(KEYINPUT103), .A3(G36gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(KEYINPUT103), .B1(new_n667_), .B2(G36gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n666_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT46), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OAI211_X1 g471(.A(KEYINPUT46), .B(new_n666_), .C1(new_n668_), .C2(new_n669_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1329gat));
  NAND4_X1  g473(.A1(new_n657_), .A2(new_n661_), .A3(G43gat), .A4(new_n366_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n352_), .B1(new_n648_), .B2(new_n412_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT105), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT105), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n675_), .A2(new_n679_), .A3(new_n676_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n678_), .A2(new_n680_), .A3(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n678_), .B2(new_n680_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1330gat));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n685_));
  INV_X1    g484(.A(new_n426_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n662_), .A2(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n685_), .B1(new_n687_), .B2(G50gat), .ZN(new_n688_));
  INV_X1    g487(.A(G50gat), .ZN(new_n689_));
  AOI211_X1 g488(.A(KEYINPUT106), .B(new_n689_), .C1(new_n662_), .C2(new_n686_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n426_), .A2(G50gat), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT107), .ZN(new_n692_));
  OAI22_X1  g491(.A1(new_n688_), .A2(new_n690_), .B1(new_n648_), .B2(new_n692_), .ZN(G1331gat));
  INV_X1    g492(.A(new_n621_), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n574_), .A2(new_n606_), .A3(new_n459_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(G57gat), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n696_), .A2(new_n697_), .A3(new_n609_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n432_), .A2(new_n459_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n699_), .A2(new_n575_), .A3(new_n605_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n701_), .A2(KEYINPUT108), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(KEYINPUT108), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n702_), .A2(new_n610_), .A3(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n698_), .B1(new_n704_), .B2(new_n697_), .ZN(G1332gat));
  OAI21_X1  g504(.A(G64gat), .B1(new_n696_), .B2(new_n614_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT48), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n614_), .A2(G64gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n707_), .B1(new_n700_), .B2(new_n708_), .ZN(G1333gat));
  OAI21_X1  g508(.A(G71gat), .B1(new_n696_), .B2(new_n412_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT49), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n412_), .A2(G71gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n711_), .B1(new_n700_), .B2(new_n712_), .ZN(G1334gat));
  NAND3_X1  g512(.A1(new_n694_), .A2(new_n686_), .A3(new_n695_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(G78gat), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT110), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n715_), .B(new_n716_), .ZN(new_n717_));
  XOR2_X1   g516(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n718_));
  AND2_X1   g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n717_), .A2(new_n718_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n426_), .A2(G78gat), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT111), .Z(new_n722_));
  OAI22_X1  g521(.A1(new_n719_), .A2(new_n720_), .B1(new_n700_), .B2(new_n722_), .ZN(G1335gat));
  NOR4_X1   g522(.A1(new_n646_), .A2(new_n432_), .A3(new_n459_), .A4(new_n606_), .ZN(new_n724_));
  AOI21_X1  g523(.A(G85gat), .B1(new_n724_), .B2(new_n610_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n606_), .A2(new_n459_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n653_), .A2(new_n654_), .A3(new_n574_), .A4(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n610_), .A2(G85gat), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT112), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n725_), .B1(new_n728_), .B2(new_n730_), .ZN(G1336gat));
  AOI21_X1  g530(.A(G92gat), .B1(new_n724_), .B2(new_n283_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT113), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n283_), .A2(G92gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n728_), .B2(new_n734_), .ZN(G1337gat));
  OAI21_X1  g534(.A(G99gat), .B1(new_n727_), .B2(new_n412_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n724_), .A2(new_n366_), .A3(new_n465_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g538(.A1(new_n724_), .A2(new_n466_), .A3(new_n686_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT52), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n727_), .A2(new_n426_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n466_), .B1(new_n742_), .B2(KEYINPUT114), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT114), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n744_), .B1(new_n727_), .B2(new_n426_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n741_), .B1(new_n743_), .B2(new_n745_), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n653_), .A2(new_n574_), .A3(new_n654_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n747_), .A2(KEYINPUT114), .A3(new_n686_), .A4(new_n726_), .ZN(new_n748_));
  AND4_X1   g547(.A1(new_n741_), .A2(new_n748_), .A3(G106gat), .A4(new_n745_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n740_), .B1(new_n746_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT53), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT53), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n752_), .B(new_n740_), .C1(new_n746_), .C2(new_n749_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(G1339gat));
  NOR2_X1   g553(.A1(new_n686_), .A2(new_n283_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n609_), .A2(new_n412_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT117), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n443_), .A2(new_n444_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(new_n456_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n444_), .B1(new_n451_), .B2(KEYINPUT116), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT116), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n448_), .A2(new_n762_), .A3(new_n450_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n760_), .B1(new_n761_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n458_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n758_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n451_), .A2(KEYINPUT116), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n767_), .A2(new_n445_), .A3(new_n763_), .ZN(new_n768_));
  OAI211_X1 g567(.A(KEYINPUT117), .B(new_n458_), .C1(new_n768_), .C2(new_n760_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n766_), .A2(new_n769_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n770_), .A2(new_n598_), .ZN(new_n771_));
  XOR2_X1   g570(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n772_));
  NAND3_X1  g571(.A1(new_n585_), .A2(new_n590_), .A3(new_n772_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n579_), .A2(new_n580_), .A3(new_n582_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n579_), .A2(new_n586_), .A3(new_n580_), .ZN(new_n775_));
  AOI22_X1  g574(.A1(new_n774_), .A2(KEYINPUT55), .B1(new_n775_), .B2(new_n581_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n773_), .A2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT56), .B1(new_n777_), .B2(new_n595_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT56), .ZN(new_n779_));
  AOI211_X1 g578(.A(new_n779_), .B(new_n597_), .C1(new_n773_), .C2(new_n776_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n771_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT58), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n771_), .B(KEYINPUT58), .C1(new_n778_), .C2(new_n780_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n543_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT119), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT119), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n543_), .A2(new_n783_), .A3(new_n787_), .A4(new_n784_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT57), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n599_), .A2(new_n770_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n597_), .B1(new_n773_), .B2(new_n776_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(KEYINPUT56), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n598_), .A2(new_n459_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n791_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  OAI211_X1 g594(.A(KEYINPUT118), .B(new_n789_), .C1(new_n795_), .C2(new_n619_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n786_), .A2(new_n788_), .A3(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n794_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n790_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n619_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(KEYINPUT57), .A3(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT57), .B1(new_n799_), .B2(new_n800_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(KEYINPUT118), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n573_), .B1(new_n797_), .B2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n652_), .A2(new_n658_), .A3(new_n606_), .ZN(new_n805_));
  OAI21_X1  g604(.A(KEYINPUT54), .B1(new_n805_), .B2(new_n459_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n575_), .A2(new_n807_), .A3(new_n460_), .A4(new_n606_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n757_), .B1(new_n804_), .B2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(G113gat), .B1(new_n810_), .B2(new_n459_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n757_), .A2(KEYINPUT59), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n806_), .A2(new_n808_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n801_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n814_), .A2(new_n802_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n658_), .B1(new_n815_), .B2(new_n785_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n812_), .B1(new_n813_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT59), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n810_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n459_), .A2(G113gat), .ZN(new_n821_));
  XOR2_X1   g620(.A(new_n821_), .B(KEYINPUT120), .Z(new_n822_));
  AOI21_X1  g621(.A(new_n811_), .B1(new_n820_), .B2(new_n822_), .ZN(G1340gat));
  NAND2_X1  g622(.A1(new_n804_), .A2(new_n809_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n757_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(KEYINPUT121), .B(G120gat), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT60), .B1(new_n605_), .B2(new_n827_), .ZN(new_n828_));
  OR3_X1    g627(.A1(new_n826_), .A2(KEYINPUT60), .A3(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n605_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n830_), .A2(new_n819_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n829_), .B1(new_n831_), .B2(new_n827_), .ZN(G1341gat));
  INV_X1    g631(.A(G127gat), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n833_), .B1(new_n826_), .B2(new_n574_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n573_), .A2(new_n833_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n817_), .B(new_n835_), .C1(new_n810_), .C2(new_n818_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT122), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT122), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n834_), .A2(new_n839_), .A3(new_n836_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(G1342gat));
  OAI21_X1  g640(.A(G134gat), .B1(new_n819_), .B2(new_n652_), .ZN(new_n842_));
  OR2_X1    g641(.A1(new_n620_), .A2(G134gat), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n826_), .B2(new_n843_), .ZN(G1343gat));
  NOR2_X1   g643(.A1(new_n426_), .A2(new_n366_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n824_), .A2(new_n845_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n609_), .A2(new_n283_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n846_), .A2(new_n460_), .A3(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(G141gat), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n849_), .B(new_n850_), .ZN(G1344gat));
  NOR3_X1   g650(.A1(new_n846_), .A2(new_n606_), .A3(new_n848_), .ZN(new_n852_));
  INV_X1    g651(.A(G148gat), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n852_), .B(new_n853_), .ZN(G1345gat));
  NAND4_X1  g653(.A1(new_n824_), .A2(new_n658_), .A3(new_n845_), .A4(new_n847_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT123), .ZN(new_n856_));
  INV_X1    g655(.A(new_n845_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(new_n804_), .B2(new_n809_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT123), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n858_), .A2(new_n859_), .A3(new_n658_), .A4(new_n847_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT61), .B(G155gat), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n856_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n861_), .B1(new_n856_), .B2(new_n860_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(G1346gat));
  NOR2_X1   g663(.A1(new_n846_), .A2(new_n848_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n620_), .ZN(new_n866_));
  AOI21_X1  g665(.A(G162gat), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n543_), .A2(G162gat), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(KEYINPUT124), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n867_), .B1(new_n865_), .B2(new_n869_), .ZN(G1347gat));
  NOR2_X1   g669(.A1(new_n813_), .A2(new_n816_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n610_), .A2(new_n614_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n412_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n426_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n871_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  OAI211_X1 g676(.A(KEYINPUT62), .B(G169gat), .C1(new_n877_), .C2(new_n460_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT62), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n871_), .A2(new_n460_), .A3(new_n875_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(new_n208_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n221_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n878_), .A2(new_n881_), .A3(new_n882_), .ZN(G1348gat));
  NAND3_X1  g682(.A1(new_n874_), .A2(G176gat), .A3(new_n605_), .ZN(new_n884_));
  AOI211_X1 g683(.A(new_n686_), .B(new_n884_), .C1(new_n804_), .C2(new_n809_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n871_), .A2(new_n606_), .A3(new_n875_), .ZN(new_n886_));
  OR3_X1    g685(.A1(new_n886_), .A2(KEYINPUT125), .A3(G176gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT125), .B1(new_n886_), .B2(G176gat), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n885_), .B1(new_n887_), .B2(new_n888_), .ZN(G1349gat));
  AND4_X1   g688(.A1(new_n217_), .A2(new_n876_), .A3(new_n572_), .A4(new_n564_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n244_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n824_), .A2(new_n426_), .A3(new_n658_), .A4(new_n874_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n890_), .B1(new_n891_), .B2(new_n892_), .ZN(G1350gat));
  OAI21_X1  g692(.A(G190gat), .B1(new_n877_), .B2(new_n652_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n876_), .A2(new_n218_), .A3(new_n866_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1351gat));
  NAND3_X1  g695(.A1(new_n858_), .A2(new_n459_), .A3(new_n872_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g697(.A1(new_n858_), .A2(new_n872_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(new_n606_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(KEYINPUT126), .B(G204gat), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(G1353gat));
  NOR3_X1   g701(.A1(KEYINPUT127), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n903_));
  OAI21_X1  g702(.A(KEYINPUT127), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n905_), .A2(new_n903_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n573_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n858_), .A2(new_n872_), .A3(new_n907_), .ZN(new_n908_));
  MUX2_X1   g707(.A(new_n903_), .B(new_n906_), .S(new_n908_), .Z(G1354gat));
  OAI21_X1  g708(.A(G218gat), .B1(new_n899_), .B2(new_n652_), .ZN(new_n910_));
  OR2_X1    g709(.A1(new_n620_), .A2(G218gat), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n899_), .B2(new_n911_), .ZN(G1355gat));
endmodule


