//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n759_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n885_, new_n886_, new_n887_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n919_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT25), .B(G183gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT26), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G190gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT77), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n206_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT26), .ZN(new_n212_));
  AOI21_X1  g011(.A(KEYINPUT77), .B1(new_n208_), .B2(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n205_), .B1(new_n210_), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT78), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT78), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n216_), .B(new_n205_), .C1(new_n210_), .C2(new_n213_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n218_), .B(new_n219_), .ZN(new_n220_));
  NOR3_X1   g019(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n215_), .A2(new_n217_), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n218_), .A2(new_n219_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n224_), .B(new_n225_), .C1(G183gat), .C2(G190gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT79), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(G169gat), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT79), .B1(G183gat), .B2(G190gat), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n228_), .B(new_n230_), .C1(new_n220_), .C2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n223_), .A2(KEYINPUT30), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT30), .B1(new_n223_), .B2(new_n232_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT81), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n235_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT81), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(new_n238_), .A3(new_n233_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G227gat), .A2(G233gat), .ZN(new_n240_));
  INV_X1    g039(.A(G71gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(G99gat), .ZN(new_n243_));
  XOR2_X1   g042(.A(G15gat), .B(G43gat), .Z(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT80), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n243_), .B(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n236_), .A2(new_n239_), .A3(new_n247_), .ZN(new_n248_));
  OAI211_X1 g047(.A(KEYINPUT81), .B(new_n246_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT82), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n248_), .A2(KEYINPUT82), .A3(new_n249_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G127gat), .B(G134gat), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(G113gat), .B(G120gat), .Z(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G113gat), .B(G120gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n254_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT31), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n252_), .A2(new_n253_), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n261_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n248_), .A2(KEYINPUT82), .A3(new_n249_), .A4(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G228gat), .A2(G233gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  OR2_X1    g066(.A1(G197gat), .A2(G204gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G197gat), .A2(G204gat), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(KEYINPUT21), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT84), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G211gat), .B(G218gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G197gat), .B(G204gat), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT21), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT84), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n268_), .A2(new_n276_), .A3(KEYINPUT21), .A4(new_n269_), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n271_), .A2(new_n272_), .A3(new_n275_), .A4(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n270_), .ZN(new_n279_));
  INV_X1    g078(.A(G218gat), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n280_), .A2(G211gat), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n280_), .A2(G211gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT85), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT85), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n272_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n279_), .A2(new_n283_), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n278_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT3), .ZN(new_n289_));
  INV_X1    g088(.A(G141gat), .ZN(new_n290_));
  INV_X1    g089(.A(G148gat), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n289_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G141gat), .A2(G148gat), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT2), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n292_), .A2(new_n295_), .A3(new_n296_), .A4(new_n297_), .ZN(new_n298_));
  OR2_X1    g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G155gat), .A2(G162gat), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(KEYINPUT1), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT1), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n303_), .A2(G155gat), .A3(G162gat), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n302_), .A2(new_n304_), .A3(new_n299_), .ZN(new_n305_));
  XOR2_X1   g104(.A(G141gat), .B(G148gat), .Z(new_n306_));
  AOI22_X1  g105(.A1(new_n298_), .A2(new_n301_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT87), .B(KEYINPUT29), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n267_), .B1(new_n288_), .B2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G78gat), .B(G106gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n287_), .A2(KEYINPUT86), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT86), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n278_), .A2(new_n314_), .A3(new_n286_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n298_), .A2(new_n301_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n305_), .A2(new_n306_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n319_), .A2(KEYINPUT83), .A3(KEYINPUT29), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT83), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT29), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n321_), .B1(new_n307_), .B2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n320_), .A2(new_n323_), .A3(new_n266_), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n310_), .B(new_n312_), .C1(new_n316_), .C2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT88), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n307_), .A2(new_n322_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G22gat), .B(G50gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT28), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n328_), .B(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n327_), .A2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n310_), .B1(new_n316_), .B2(new_n324_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(new_n311_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n325_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n332_), .A2(new_n335_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n334_), .A2(KEYINPUT88), .A3(new_n325_), .A4(new_n331_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G64gat), .B(G92gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT91), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G8gat), .B(G36gat), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n343_), .B(new_n344_), .Z(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT32), .ZN(new_n346_));
  INV_X1    g145(.A(new_n315_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n314_), .B1(new_n278_), .B2(new_n286_), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n223_), .B(new_n232_), .C1(new_n347_), .C2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT20), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n230_), .A2(new_n226_), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n208_), .A2(new_n212_), .A3(KEYINPUT89), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT89), .B1(new_n208_), .B2(new_n212_), .ZN(new_n353_));
  INV_X1    g152(.A(G183gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT25), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT25), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(G183gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  NOR3_X1   g157(.A1(new_n352_), .A2(new_n353_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n221_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n205_), .A2(new_n360_), .A3(new_n224_), .A4(new_n225_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n351_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n350_), .B1(new_n362_), .B2(new_n287_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n349_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G226gat), .A2(G233gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT19), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n366_), .ZN(new_n368_));
  OAI211_X1 g167(.A(KEYINPUT20), .B(new_n368_), .C1(new_n362_), .C2(new_n287_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n347_), .A2(new_n348_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n223_), .A2(new_n232_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n369_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n346_), .A2(new_n367_), .A3(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G1gat), .B(G29gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G57gat), .B(G85gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G225gat), .A2(G233gat), .ZN(new_n381_));
  NOR3_X1   g180(.A1(new_n319_), .A2(new_n260_), .A3(KEYINPUT92), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT92), .ZN(new_n383_));
  AOI22_X1  g182(.A1(new_n307_), .A2(new_n383_), .B1(new_n259_), .B2(new_n257_), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT4), .B1(new_n382_), .B2(new_n384_), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n260_), .A2(new_n307_), .A3(KEYINPUT4), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n381_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n381_), .ZN(new_n389_));
  NOR3_X1   g188(.A1(new_n382_), .A2(new_n384_), .A3(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n380_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT4), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n257_), .A2(new_n259_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n393_), .A2(new_n307_), .A3(new_n383_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n260_), .B1(new_n319_), .B2(KEYINPUT92), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n392_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n389_), .B1(new_n396_), .B2(new_n386_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n390_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n397_), .A2(new_n398_), .A3(new_n379_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n391_), .A2(KEYINPUT101), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT101), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n397_), .A2(new_n398_), .A3(new_n401_), .A4(new_n379_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n374_), .A2(new_n400_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n370_), .A2(new_n371_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n287_), .B1(new_n362_), .B2(KEYINPUT97), .ZN(new_n405_));
  INV_X1    g204(.A(new_n353_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n208_), .A2(new_n212_), .A3(KEYINPUT89), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(new_n407_), .A3(new_n206_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n203_), .A2(new_n204_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n224_), .A2(new_n225_), .ZN(new_n410_));
  NOR3_X1   g209(.A1(new_n409_), .A2(new_n410_), .A3(new_n221_), .ZN(new_n411_));
  AOI22_X1  g210(.A1(new_n408_), .A2(new_n411_), .B1(new_n226_), .B2(new_n230_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT97), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n350_), .B1(new_n405_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT98), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n404_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  AOI211_X1 g216(.A(KEYINPUT98), .B(new_n350_), .C1(new_n405_), .C2(new_n414_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n366_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT99), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  OAI211_X1 g220(.A(KEYINPUT99), .B(new_n366_), .C1(new_n417_), .C2(new_n418_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n349_), .A2(new_n368_), .A3(new_n363_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT100), .ZN(new_n424_));
  OR2_X1    g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n424_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n421_), .A2(new_n422_), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n346_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n403_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n345_), .B1(new_n367_), .B2(new_n373_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n368_), .B1(new_n349_), .B2(new_n363_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n343_), .B(new_n344_), .ZN(new_n433_));
  NOR3_X1   g232(.A1(new_n432_), .A2(new_n433_), .A3(new_n372_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n431_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n391_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT94), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT33), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT33), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n391_), .A2(KEYINPUT94), .A3(new_n439_), .ZN(new_n440_));
  NOR3_X1   g239(.A1(new_n396_), .A2(new_n389_), .A3(new_n386_), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n441_), .A2(KEYINPUT96), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n396_), .A2(new_n386_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n443_), .A2(KEYINPUT96), .A3(new_n381_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT95), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n381_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n445_), .B1(new_n446_), .B2(new_n380_), .ZN(new_n447_));
  OR3_X1    g246(.A1(new_n446_), .A2(new_n380_), .A3(new_n445_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n442_), .A2(new_n444_), .A3(new_n447_), .A4(new_n448_), .ZN(new_n449_));
  AND4_X1   g248(.A1(new_n435_), .A2(new_n438_), .A3(new_n440_), .A4(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n339_), .B1(new_n430_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT27), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n434_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n454_), .B1(new_n428_), .B2(new_n433_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n452_), .B1(new_n431_), .B2(new_n434_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n400_), .A2(new_n402_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n338_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT102), .B1(new_n455_), .B2(new_n458_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n338_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT102), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n419_), .A2(new_n420_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n345_), .B1(new_n462_), .B2(new_n422_), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n460_), .B(new_n461_), .C1(new_n463_), .C2(new_n454_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n451_), .A2(new_n459_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n456_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n428_), .A2(new_n433_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n466_), .B1(new_n467_), .B2(new_n453_), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n262_), .A2(new_n264_), .A3(new_n457_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT103), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n468_), .A2(new_n469_), .A3(new_n470_), .A4(new_n339_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n456_), .B(new_n339_), .C1(new_n463_), .C2(new_n454_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n262_), .A2(new_n264_), .A3(new_n457_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT103), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  AOI22_X1  g273(.A1(new_n265_), .A2(new_n465_), .B1(new_n471_), .B2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G29gat), .B(G36gat), .ZN(new_n476_));
  OR2_X1    g275(.A1(new_n476_), .A2(KEYINPUT73), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(KEYINPUT73), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G43gat), .B(G50gat), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n477_), .A2(new_n478_), .A3(new_n480_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT15), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G1gat), .B(G8gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT74), .ZN(new_n487_));
  INV_X1    g286(.A(G15gat), .ZN(new_n488_));
  INV_X1    g287(.A(G22gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G15gat), .A2(G22gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G1gat), .A2(G8gat), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n490_), .A2(new_n491_), .B1(KEYINPUT14), .B2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n487_), .B(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n485_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n494_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(new_n484_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G229gat), .A2(G233gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n495_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n494_), .B(new_n484_), .Z(new_n500_));
  INV_X1    g299(.A(new_n498_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n499_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G113gat), .B(G141gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT76), .ZN(new_n505_));
  XOR2_X1   g304(.A(G169gat), .B(G197gat), .Z(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n503_), .B(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT104), .B1(new_n475_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n465_), .A2(new_n265_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n471_), .A2(new_n474_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT104), .ZN(new_n513_));
  INV_X1    g312(.A(new_n508_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n512_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(G85gat), .ZN(new_n516_));
  INV_X1    g315(.A(G92gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT9), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G85gat), .A2(G92gat), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n520_), .A2(KEYINPUT64), .A3(new_n519_), .ZN(new_n521_));
  AOI21_X1  g320(.A(KEYINPUT64), .B1(new_n520_), .B2(new_n519_), .ZN(new_n522_));
  OAI221_X1 g321(.A(new_n518_), .B1(new_n519_), .B2(new_n520_), .C1(new_n521_), .C2(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(KEYINPUT10), .B(G99gat), .Z(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT6), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT65), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT65), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT6), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G99gat), .A2(G106gat), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n533_));
  INV_X1    g332(.A(new_n531_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  OAI221_X1 g334(.A(new_n523_), .B1(G106gat), .B2(new_n525_), .C1(new_n532_), .C2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(G99gat), .A2(G106gat), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT7), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n530_), .A2(new_n531_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n533_), .A2(new_n534_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n539_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n518_), .A2(new_n520_), .ZN(new_n543_));
  NOR3_X1   g342(.A1(new_n542_), .A2(KEYINPUT8), .A3(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT8), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n537_), .B(KEYINPUT7), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n546_), .B1(new_n532_), .B2(new_n535_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n543_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n545_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n536_), .B1(new_n544_), .B2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G57gat), .B(G64gat), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT11), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT67), .ZN(new_n553_));
  XOR2_X1   g352(.A(G71gat), .B(G78gat), .Z(new_n554_));
  OAI21_X1  g353(.A(new_n554_), .B1(KEYINPUT11), .B2(new_n551_), .ZN(new_n555_));
  OR2_X1    g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n553_), .A2(new_n555_), .ZN(new_n557_));
  AND4_X1   g356(.A1(KEYINPUT12), .A2(new_n550_), .A3(new_n556_), .A4(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n557_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT66), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n550_), .A2(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(KEYINPUT8), .B1(new_n542_), .B2(new_n543_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n547_), .A2(new_n545_), .A3(new_n548_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(KEYINPUT66), .B1(new_n565_), .B2(new_n536_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n560_), .B1(new_n562_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT12), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n558_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n550_), .A2(new_n561_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n565_), .A2(KEYINPUT66), .A3(new_n536_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n570_), .A2(new_n559_), .A3(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G230gat), .A2(G233gat), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n572_), .A2(KEYINPUT69), .A3(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(KEYINPUT69), .B1(new_n572_), .B2(new_n573_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n569_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n567_), .A2(KEYINPUT68), .A3(new_n572_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT68), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n578_), .B(new_n560_), .C1(new_n562_), .C2(new_n566_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n573_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n577_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G120gat), .B(G148gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT5), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G176gat), .B(G204gat), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n583_), .B(new_n584_), .Z(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n576_), .A2(new_n581_), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(KEYINPUT70), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT70), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n576_), .A2(new_n589_), .A3(new_n581_), .A4(new_n586_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n576_), .A2(new_n581_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(new_n585_), .ZN(new_n593_));
  AND3_X1   g392(.A1(new_n591_), .A2(KEYINPUT13), .A3(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(KEYINPUT13), .B1(new_n591_), .B2(new_n593_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n509_), .A2(new_n515_), .A3(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G190gat), .B(G218gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G134gat), .B(G162gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n600_), .A2(KEYINPUT36), .ZN(new_n601_));
  XOR2_X1   g400(.A(KEYINPUT71), .B(KEYINPUT35), .Z(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G232gat), .A2(G233gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT34), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n606_), .B1(new_n485_), .B2(new_n550_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n570_), .A2(new_n571_), .A3(new_n484_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n603_), .A2(new_n605_), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n609_), .B(KEYINPUT72), .Z(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n607_), .A2(new_n608_), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n611_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n601_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n614_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n600_), .B(KEYINPUT36), .Z(new_n617_));
  NAND3_X1  g416(.A1(new_n616_), .A2(new_n612_), .A3(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n615_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT37), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT37), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n615_), .A2(new_n618_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G231gat), .A2(G233gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n559_), .B(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(new_n496_), .ZN(new_n627_));
  XOR2_X1   g426(.A(G127gat), .B(G155gat), .Z(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT16), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G183gat), .B(G211gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT17), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT75), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n631_), .A2(new_n634_), .A3(new_n632_), .ZN(new_n635_));
  OR3_X1    g434(.A1(new_n627_), .A2(new_n633_), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n627_), .A2(new_n635_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n624_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n597_), .A2(new_n639_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n640_), .A2(G1gat), .A3(new_n457_), .ZN(new_n641_));
  XOR2_X1   g440(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n642_));
  OR2_X1    g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n595_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n591_), .A2(KEYINPUT13), .A3(new_n593_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n646_), .A2(new_n638_), .A3(new_n508_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n647_), .A2(new_n619_), .A3(new_n512_), .ZN(new_n648_));
  OAI21_X1  g447(.A(G1gat), .B1(new_n648_), .B2(new_n457_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n641_), .A2(new_n642_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n643_), .A2(new_n649_), .A3(new_n650_), .ZN(G1324gat));
  OAI21_X1  g450(.A(G8gat), .B1(new_n648_), .B2(new_n468_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT39), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n468_), .A2(G8gat), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n640_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT106), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n640_), .A2(KEYINPUT106), .A3(new_n654_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n653_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT40), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  OAI211_X1 g460(.A(KEYINPUT40), .B(new_n653_), .C1(new_n657_), .C2(new_n658_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1325gat));
  OAI21_X1  g462(.A(G15gat), .B1(new_n648_), .B2(new_n265_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT41), .Z(new_n665_));
  INV_X1    g464(.A(new_n265_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(new_n488_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n665_), .B1(new_n640_), .B2(new_n667_), .ZN(G1326gat));
  OAI21_X1  g467(.A(G22gat), .B1(new_n648_), .B2(new_n339_), .ZN(new_n669_));
  XOR2_X1   g468(.A(KEYINPUT107), .B(KEYINPUT42), .Z(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n338_), .A2(new_n489_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(new_n640_), .B2(new_n672_), .ZN(G1327gat));
  NAND3_X1  g472(.A1(new_n596_), .A2(new_n638_), .A3(new_n514_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT108), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n596_), .A2(KEYINPUT108), .A3(new_n638_), .A4(new_n514_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT109), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n623_), .A2(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(KEYINPUT109), .B1(new_n620_), .B2(new_n622_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(KEYINPUT43), .B1(new_n475_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT43), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n512_), .A2(new_n624_), .A3(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n678_), .A2(new_n686_), .ZN(new_n687_));
  XOR2_X1   g486(.A(KEYINPUT110), .B(KEYINPUT44), .Z(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n678_), .A2(new_n686_), .A3(KEYINPUT44), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(G29gat), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n692_), .A2(new_n693_), .A3(new_n457_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n457_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n638_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n696_), .A2(new_n619_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n597_), .A2(new_n695_), .A3(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n694_), .B1(new_n693_), .B2(new_n698_), .ZN(G1328gat));
  INV_X1    g498(.A(new_n468_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n690_), .A2(new_n700_), .A3(new_n691_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(G36gat), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT111), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n468_), .A2(G36gat), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n597_), .A2(new_n703_), .A3(new_n697_), .A4(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT45), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n509_), .A2(new_n515_), .A3(new_n596_), .A4(new_n697_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n704_), .ZN(new_n708_));
  OAI21_X1  g507(.A(KEYINPUT111), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n705_), .A2(new_n706_), .A3(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n706_), .B1(new_n705_), .B2(new_n709_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n702_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(KEYINPUT112), .A2(KEYINPUT46), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  OAI221_X1 g513(.A(new_n702_), .B1(KEYINPUT112), .B2(KEYINPUT46), .C1(new_n710_), .C2(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1329gat));
  INV_X1    g515(.A(G43gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n717_), .B1(new_n707_), .B2(new_n265_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n265_), .A2(new_n717_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n718_), .B1(new_n692_), .B2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g521(.A(G50gat), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n692_), .A2(new_n723_), .A3(new_n339_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n597_), .A2(new_n338_), .A3(new_n697_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n723_), .B2(new_n725_), .ZN(G1331gat));
  NAND2_X1  g525(.A1(new_n646_), .A2(new_n508_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n727_), .A2(new_n475_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n728_), .A2(new_n639_), .ZN(new_n729_));
  INV_X1    g528(.A(G57gat), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n729_), .A2(new_n730_), .A3(new_n695_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n619_), .ZN(new_n732_));
  NOR4_X1   g531(.A1(new_n727_), .A2(new_n475_), .A3(new_n638_), .A4(new_n732_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n733_), .A2(new_n695_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n731_), .B1(new_n734_), .B2(new_n730_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT113), .ZN(G1332gat));
  INV_X1    g535(.A(G64gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n733_), .B2(new_n700_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT48), .Z(new_n739_));
  NAND3_X1  g538(.A1(new_n729_), .A2(new_n737_), .A3(new_n700_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1333gat));
  AOI21_X1  g540(.A(new_n241_), .B1(new_n733_), .B2(new_n666_), .ZN(new_n742_));
  XOR2_X1   g541(.A(KEYINPUT114), .B(KEYINPUT49), .Z(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n729_), .A2(new_n241_), .A3(new_n666_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1334gat));
  INV_X1    g545(.A(G78gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n733_), .B2(new_n338_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT50), .Z(new_n749_));
  NAND3_X1  g548(.A1(new_n729_), .A2(new_n747_), .A3(new_n338_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1335gat));
  NAND2_X1  g550(.A1(new_n728_), .A2(new_n697_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n753_), .A2(new_n516_), .A3(new_n695_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n646_), .A2(new_n638_), .A3(new_n508_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n683_), .B2(new_n685_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n756_), .A2(new_n695_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n754_), .B1(new_n757_), .B2(new_n516_), .ZN(G1336gat));
  AOI21_X1  g557(.A(new_n517_), .B1(new_n756_), .B2(new_n700_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n752_), .A2(G92gat), .A3(new_n468_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT115), .ZN(G1337gat));
  NOR3_X1   g561(.A1(new_n752_), .A2(new_n525_), .A3(new_n265_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n756_), .A2(new_n666_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(G99gat), .B2(new_n764_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n765_), .B(new_n766_), .ZN(G1338gat));
  INV_X1    g566(.A(G106gat), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n753_), .A2(new_n768_), .A3(new_n338_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(KEYINPUT118), .A2(KEYINPUT52), .ZN(new_n770_));
  INV_X1    g569(.A(new_n755_), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n680_), .A2(new_n681_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n684_), .B1(new_n512_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n624_), .A2(new_n684_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n475_), .A2(new_n774_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n338_), .B(new_n771_), .C1(new_n773_), .C2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT117), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n686_), .A2(KEYINPUT117), .A3(new_n338_), .A4(new_n771_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n768_), .B1(KEYINPUT118), .B2(KEYINPUT52), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n770_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n770_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n781_), .ZN(new_n784_));
  AOI211_X1 g583(.A(new_n783_), .B(new_n784_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n769_), .B1(new_n782_), .B2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT53), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n788_), .B(new_n769_), .C1(new_n782_), .C2(new_n785_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(G1339gat));
  INV_X1    g589(.A(KEYINPUT58), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n576_), .A2(new_n792_), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n569_), .B(KEYINPUT55), .C1(new_n574_), .C2(new_n575_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n567_), .A2(new_n568_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n558_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n796_), .A3(new_n572_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n580_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n793_), .A2(new_n794_), .A3(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n799_), .A2(KEYINPUT56), .A3(new_n585_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  AOI22_X1  g600(.A1(new_n576_), .A2(new_n792_), .B1(new_n580_), .B2(new_n797_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n586_), .B1(new_n802_), .B2(new_n794_), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT121), .B1(new_n803_), .B2(KEYINPUT56), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n799_), .A2(new_n585_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT121), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT56), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n805_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n801_), .B1(new_n804_), .B2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n499_), .A2(new_n502_), .A3(new_n507_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n507_), .B1(new_n500_), .B2(new_n498_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n495_), .A2(new_n497_), .A3(new_n501_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n810_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n591_), .A2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n791_), .B1(new_n809_), .B2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n806_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n818_));
  AOI211_X1 g617(.A(KEYINPUT121), .B(KEYINPUT56), .C1(new_n799_), .C2(new_n585_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n800_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n816_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(KEYINPUT58), .A3(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n817_), .A2(new_n822_), .A3(new_n624_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n805_), .A2(new_n807_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT120), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n826_), .A3(new_n800_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n508_), .B1(new_n588_), .B2(new_n590_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n799_), .A2(KEYINPUT120), .A3(KEYINPUT56), .A4(new_n585_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n591_), .A2(new_n593_), .ZN(new_n831_));
  AOI22_X1  g630(.A1(new_n827_), .A2(new_n830_), .B1(new_n831_), .B2(new_n815_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n824_), .B1(new_n832_), .B2(new_n732_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n800_), .A2(new_n826_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT56), .B1(new_n799_), .B2(new_n585_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n829_), .B(new_n828_), .C1(new_n834_), .C2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n831_), .A2(new_n815_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n838_), .A2(KEYINPUT57), .A3(new_n619_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n823_), .A2(new_n833_), .A3(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n638_), .A2(new_n514_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n644_), .A2(new_n645_), .A3(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n623_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT119), .B1(new_n596_), .B2(new_n841_), .ZN(new_n845_));
  OAI21_X1  g644(.A(KEYINPUT54), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n842_), .A2(new_n843_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n596_), .A2(KEYINPUT119), .A3(new_n841_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n847_), .A2(new_n848_), .A3(new_n849_), .A4(new_n623_), .ZN(new_n850_));
  AOI22_X1  g649(.A1(new_n840_), .A2(new_n638_), .B1(new_n846_), .B2(new_n850_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n472_), .A2(new_n265_), .A3(new_n457_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n851_), .A2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(G113gat), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n854_), .A2(new_n855_), .A3(new_n514_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(KEYINPUT59), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n851_), .B2(new_n853_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n508_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n856_), .B1(new_n860_), .B2(new_n855_), .ZN(G1340gat));
  AOI21_X1  g660(.A(new_n596_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n862_));
  INV_X1    g661(.A(G120gat), .ZN(new_n863_));
  INV_X1    g662(.A(new_n854_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n596_), .B2(KEYINPUT60), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(KEYINPUT60), .B2(new_n863_), .ZN(new_n866_));
  OAI22_X1  g665(.A1(new_n862_), .A2(new_n863_), .B1(new_n864_), .B2(new_n866_), .ZN(G1341gat));
  AOI21_X1  g666(.A(G127gat), .B1(new_n854_), .B2(new_n696_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n857_), .A2(new_n859_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n696_), .A2(G127gat), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(KEYINPUT122), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n868_), .B1(new_n869_), .B2(new_n871_), .ZN(G1342gat));
  INV_X1    g671(.A(G134gat), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n854_), .A2(new_n873_), .A3(new_n732_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n623_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(new_n873_), .ZN(G1343gat));
  NOR2_X1   g675(.A1(new_n851_), .A2(new_n666_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n700_), .A2(new_n457_), .A3(new_n339_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n879_), .A2(new_n290_), .A3(new_n514_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n877_), .A2(new_n878_), .ZN(new_n881_));
  OAI21_X1  g680(.A(G141gat), .B1(new_n881_), .B2(new_n508_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(G1344gat));
  XNOR2_X1  g682(.A(KEYINPUT123), .B(G148gat), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n879_), .A2(new_n646_), .A3(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n884_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n886_), .B1(new_n881_), .B2(new_n596_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(G1345gat));
  XNOR2_X1  g687(.A(KEYINPUT61), .B(G155gat), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n879_), .A2(new_n696_), .A3(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n889_), .B1(new_n881_), .B2(new_n638_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1346gat));
  NAND2_X1  g692(.A1(new_n879_), .A2(new_n732_), .ZN(new_n894_));
  INV_X1    g693(.A(G162gat), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n682_), .A2(new_n895_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(KEYINPUT124), .ZN(new_n897_));
  AOI22_X1  g696(.A1(new_n894_), .A2(new_n895_), .B1(new_n879_), .B2(new_n897_), .ZN(G1347gat));
  INV_X1    g697(.A(G169gat), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n468_), .A2(new_n338_), .A3(new_n473_), .ZN(new_n900_));
  AOI21_X1  g699(.A(KEYINPUT57), .B1(new_n838_), .B2(new_n619_), .ZN(new_n901_));
  AOI211_X1 g700(.A(new_n824_), .B(new_n732_), .C1(new_n836_), .C2(new_n837_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n696_), .B1(new_n903_), .B2(new_n823_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n846_), .A2(new_n850_), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n514_), .B(new_n900_), .C1(new_n904_), .C2(new_n905_), .ZN(new_n906_));
  OAI211_X1 g705(.A(KEYINPUT62), .B(new_n899_), .C1(new_n906_), .C2(KEYINPUT22), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n908_));
  INV_X1    g707(.A(new_n900_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n851_), .A2(new_n508_), .A3(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT22), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n908_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(G169gat), .B1(new_n906_), .B2(KEYINPUT62), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n907_), .B1(new_n912_), .B2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(G1348gat));
  NOR2_X1   g714(.A1(new_n851_), .A2(new_n909_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n646_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(G176gat), .ZN(G1349gat));
  AOI21_X1  g717(.A(G183gat), .B1(new_n916_), .B2(new_n696_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n916_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n638_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n919_), .B1(new_n921_), .B2(new_n358_), .ZN(G1350gat));
  OAI211_X1 g721(.A(new_n624_), .B(new_n900_), .C1(new_n904_), .C2(new_n905_), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT125), .ZN(new_n924_));
  AND3_X1   g723(.A1(new_n923_), .A2(new_n924_), .A3(G190gat), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n924_), .B1(new_n923_), .B2(G190gat), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n732_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n927_));
  OAI22_X1  g726(.A1(new_n925_), .A2(new_n926_), .B1(new_n920_), .B2(new_n927_), .ZN(G1351gat));
  INV_X1    g727(.A(G197gat), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n468_), .A2(new_n695_), .A3(new_n339_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n877_), .A2(new_n930_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n929_), .B1(new_n931_), .B2(new_n508_), .ZN(new_n932_));
  NAND4_X1  g731(.A1(new_n877_), .A2(G197gat), .A3(new_n514_), .A4(new_n930_), .ZN(new_n933_));
  AND2_X1   g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1352gat));
  INV_X1    g733(.A(KEYINPUT126), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(G204gat), .ZN(new_n936_));
  XOR2_X1   g735(.A(new_n936_), .B(KEYINPUT127), .Z(new_n937_));
  INV_X1    g736(.A(new_n937_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n938_), .B1(new_n931_), .B2(new_n596_), .ZN(new_n939_));
  NAND4_X1  g738(.A1(new_n877_), .A2(new_n646_), .A3(new_n930_), .A4(new_n937_), .ZN(new_n940_));
  AND2_X1   g739(.A1(new_n939_), .A2(new_n940_), .ZN(G1353gat));
  AND2_X1   g740(.A1(new_n877_), .A2(new_n930_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(KEYINPUT63), .B(G211gat), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n942_), .A2(new_n696_), .A3(new_n943_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n931_), .A2(new_n638_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n944_), .B1(new_n945_), .B2(new_n946_), .ZN(G1354gat));
  NAND3_X1  g746(.A1(new_n942_), .A2(new_n280_), .A3(new_n732_), .ZN(new_n948_));
  OAI21_X1  g747(.A(G218gat), .B1(new_n931_), .B2(new_n623_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n948_), .A2(new_n949_), .ZN(G1355gat));
endmodule


