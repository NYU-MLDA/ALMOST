//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 1 1 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n651_, new_n652_, new_n653_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n782_, new_n783_,
    new_n784_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_;
  XOR2_X1   g000(.A(G155gat), .B(G162gat), .Z(new_n202_));
  INV_X1    g001(.A(G141gat), .ZN(new_n203_));
  INV_X1    g002(.A(G148gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n203_), .A2(new_n204_), .A3(KEYINPUT84), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT3), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  XOR2_X1   g006(.A(new_n207_), .B(KEYINPUT2), .Z(new_n208_));
  OAI21_X1  g007(.A(new_n202_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n202_), .A2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT83), .ZN(new_n213_));
  NAND3_X1  g012(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n211_), .A2(new_n213_), .A3(new_n207_), .A4(new_n214_), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n209_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G127gat), .B(G134gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G113gat), .B(G120gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  XOR2_X1   g018(.A(new_n216_), .B(new_n219_), .Z(new_n220_));
  NAND2_X1  g019(.A1(G225gat), .A2(G233gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(new_n222_), .B(KEYINPUT91), .Z(new_n223_));
  NAND2_X1  g022(.A1(new_n220_), .A2(KEYINPUT4), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT90), .ZN(new_n225_));
  INV_X1    g024(.A(new_n221_), .ZN(new_n226_));
  OR3_X1    g025(.A1(new_n216_), .A2(KEYINPUT4), .A3(new_n219_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT90), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n220_), .A2(new_n228_), .A3(KEYINPUT4), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .A4(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n223_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G1gat), .B(G29gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(G85gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT0), .B(G57gat), .ZN(new_n234_));
  XOR2_X1   g033(.A(new_n233_), .B(new_n234_), .Z(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT97), .B1(new_n231_), .B2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n223_), .A2(new_n230_), .A3(new_n235_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n223_), .A2(KEYINPUT97), .A3(new_n235_), .A4(new_n230_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT87), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT29), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n216_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT28), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G22gat), .B(G50gat), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n244_), .A2(new_n246_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n241_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n249_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n251_), .A2(new_n247_), .A3(KEYINPUT87), .ZN(new_n252_));
  INV_X1    g051(.A(G228gat), .ZN(new_n253_));
  INV_X1    g052(.A(G233gat), .ZN(new_n254_));
  NOR3_X1   g053(.A1(new_n253_), .A2(new_n254_), .A3(KEYINPUT85), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G197gat), .B(G204gat), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n258_), .A2(KEYINPUT21), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(KEYINPUT21), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G211gat), .B(G218gat), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n260_), .A2(new_n261_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n264_), .B1(new_n216_), .B2(new_n242_), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT85), .B1(new_n253_), .B2(new_n254_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n250_), .A2(new_n252_), .A3(new_n256_), .A4(new_n268_), .ZN(new_n269_));
  OAI221_X1 g068(.A(new_n241_), .B1(new_n255_), .B2(new_n267_), .C1(new_n248_), .C2(new_n249_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G78gat), .B(G106gat), .ZN(new_n272_));
  XOR2_X1   g071(.A(new_n272_), .B(KEYINPUT86), .Z(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n269_), .A2(new_n270_), .A3(new_n273_), .ZN(new_n276_));
  AOI22_X1  g075(.A1(new_n239_), .A2(new_n240_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT27), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT25), .B(G183gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT26), .B(G190gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G183gat), .A2(G190gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT23), .ZN(new_n283_));
  OR2_X1    g082(.A1(G169gat), .A2(G176gat), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n284_), .A2(KEYINPUT24), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(KEYINPUT24), .A3(new_n286_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n281_), .A2(new_n283_), .A3(new_n285_), .A4(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT79), .B(G176gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT22), .B(G169gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(new_n286_), .ZN(new_n292_));
  AND2_X1   g091(.A1(new_n292_), .A2(KEYINPUT80), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n283_), .B1(G183gat), .B2(G190gat), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n294_), .B1(new_n292_), .B2(KEYINPUT80), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n288_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n296_), .B(KEYINPUT81), .Z(new_n297_));
  INV_X1    g096(.A(new_n264_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n292_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n300_), .A2(KEYINPUT88), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT88), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n294_), .B1(new_n292_), .B2(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n288_), .B1(new_n301_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n264_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n299_), .A2(KEYINPUT20), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G226gat), .A2(G233gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT19), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT89), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n304_), .A2(new_n264_), .ZN(new_n311_));
  OAI211_X1 g110(.A(KEYINPUT20), .B(new_n311_), .C1(new_n297_), .C2(new_n298_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n312_), .A2(new_n308_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT89), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n306_), .A2(new_n314_), .A3(new_n308_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n310_), .A2(new_n313_), .A3(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G8gat), .B(G36gat), .ZN(new_n317_));
  INV_X1    g116(.A(G92gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT18), .B(G64gat), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n319_), .B(new_n320_), .Z(new_n321_));
  NAND2_X1  g120(.A1(new_n316_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n316_), .A2(new_n321_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n278_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n324_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n312_), .A2(new_n308_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n327_), .B1(new_n308_), .B2(new_n306_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(new_n321_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n326_), .A2(KEYINPUT27), .A3(new_n329_), .ZN(new_n330_));
  XOR2_X1   g129(.A(G15gat), .B(G43gat), .Z(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT31), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n297_), .B(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(G71gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n219_), .B(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G227gat), .A2(G233gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT30), .B(G99gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n333_), .B(new_n339_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n277_), .A2(new_n325_), .A3(new_n330_), .A4(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT98), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n223_), .A2(new_n230_), .A3(KEYINPUT33), .A4(new_n235_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT92), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n235_), .B1(new_n220_), .B2(new_n226_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n225_), .A2(new_n227_), .A3(new_n229_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n346_), .B1(new_n347_), .B2(new_n226_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n345_), .A2(new_n322_), .A3(new_n326_), .A4(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT93), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n238_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT33), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n223_), .A2(new_n230_), .A3(KEYINPUT93), .A4(new_n235_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT94), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT94), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n351_), .A2(new_n356_), .A3(new_n352_), .A4(new_n353_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT32), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n321_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n328_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n239_), .A2(new_n240_), .A3(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n360_), .B(KEYINPUT95), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n310_), .A2(new_n313_), .A3(new_n315_), .A4(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT96), .ZN(new_n365_));
  OAI22_X1  g164(.A1(new_n349_), .A2(new_n358_), .B1(new_n362_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n275_), .A2(new_n276_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n325_), .A2(new_n330_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n239_), .A2(new_n240_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n370_), .A2(new_n367_), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n366_), .A2(new_n367_), .B1(new_n368_), .B2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n340_), .B(KEYINPUT82), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n343_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G71gat), .B(G78gat), .ZN(new_n376_));
  OR2_X1    g175(.A1(G57gat), .A2(G64gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G57gat), .A2(G64gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT11), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT11), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n377_), .A2(new_n381_), .A3(new_n378_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n376_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n376_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n384_), .B1(KEYINPUT11), .B2(new_n379_), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT12), .B1(new_n383_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  AND3_X1   g186(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT65), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G99gat), .A2(G106gat), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT6), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT65), .ZN(new_n394_));
  NAND3_X1  g193(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n393_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n390_), .A2(new_n396_), .ZN(new_n397_));
  AND2_X1   g196(.A1(G85gat), .A2(G92gat), .ZN(new_n398_));
  NOR2_X1   g197(.A1(G85gat), .A2(G92gat), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT9), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT9), .ZN(new_n401_));
  INV_X1    g200(.A(G85gat), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n401_), .B1(new_n402_), .B2(new_n318_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n400_), .A2(KEYINPUT64), .A3(new_n403_), .ZN(new_n404_));
  XOR2_X1   g203(.A(KEYINPUT10), .B(G99gat), .Z(new_n405_));
  INV_X1    g204(.A(G106gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT64), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n398_), .A2(new_n408_), .A3(KEYINPUT9), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n397_), .A2(new_n404_), .A3(new_n407_), .A4(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n398_), .A2(new_n399_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT8), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT7), .ZN(new_n414_));
  INV_X1    g213(.A(G99gat), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n415_), .A3(new_n406_), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n413_), .B1(new_n397_), .B2(new_n418_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n416_), .A2(new_n393_), .A3(new_n395_), .A4(new_n417_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n412_), .B1(new_n420_), .B2(new_n411_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n410_), .B(KEYINPUT66), .C1(new_n419_), .C2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n398_), .A2(new_n399_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n388_), .A2(new_n389_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n424_), .B1(new_n418_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n416_), .A2(new_n417_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n427_), .B1(new_n390_), .B2(new_n396_), .ZN(new_n428_));
  OAI22_X1  g227(.A1(new_n426_), .A2(new_n412_), .B1(new_n428_), .B2(new_n413_), .ZN(new_n429_));
  AOI21_X1  g228(.A(KEYINPUT66), .B1(new_n429_), .B2(new_n410_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n387_), .B1(new_n423_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT67), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G230gat), .A2(G233gat), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n410_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n434_));
  OR2_X1    g233(.A1(new_n383_), .A2(new_n385_), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT12), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n435_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT66), .ZN(new_n439_));
  NOR3_X1   g238(.A1(new_n388_), .A2(new_n389_), .A3(KEYINPUT65), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n394_), .B1(new_n393_), .B2(new_n395_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n418_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n413_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n420_), .A2(new_n411_), .ZN(new_n444_));
  AOI22_X1  g243(.A1(new_n442_), .A2(new_n443_), .B1(new_n444_), .B2(KEYINPUT8), .ZN(new_n445_));
  AND4_X1   g244(.A1(new_n397_), .A2(new_n404_), .A3(new_n407_), .A4(new_n409_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n439_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n422_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT67), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n448_), .A2(new_n449_), .A3(new_n387_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n432_), .A2(new_n433_), .A3(new_n438_), .A4(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n434_), .B(new_n435_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n433_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n451_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT5), .B(G176gat), .ZN(new_n456_));
  INV_X1    g255(.A(G204gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G120gat), .B(G148gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT68), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n455_), .B(new_n461_), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n462_), .A2(KEYINPUT13), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(KEYINPUT13), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G229gat), .A2(G233gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT76), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G15gat), .B(G22gat), .ZN(new_n469_));
  INV_X1    g268(.A(G1gat), .ZN(new_n470_));
  INV_X1    g269(.A(G8gat), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT14), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G1gat), .B(G8gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  XOR2_X1   g274(.A(G29gat), .B(G36gat), .Z(new_n476_));
  XNOR2_X1  g275(.A(G43gat), .B(G50gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n475_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT75), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT75), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n481_), .B1(new_n475_), .B2(new_n478_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n475_), .A2(new_n478_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n468_), .B1(new_n483_), .B2(new_n485_), .ZN(new_n486_));
  AOI211_X1 g285(.A(KEYINPUT76), .B(new_n484_), .C1(new_n480_), .C2(new_n482_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n467_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n478_), .B(KEYINPUT15), .Z(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(new_n475_), .ZN(new_n490_));
  AND3_X1   g289(.A1(new_n490_), .A2(new_n483_), .A3(new_n466_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n488_), .A2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G113gat), .B(G141gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT77), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G169gat), .B(G197gat), .ZN(new_n496_));
  XOR2_X1   g295(.A(new_n495_), .B(new_n496_), .Z(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT78), .B1(new_n493_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n482_), .ZN(new_n500_));
  NOR3_X1   g299(.A1(new_n475_), .A2(new_n478_), .A3(new_n481_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n485_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT76), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n483_), .A2(new_n468_), .A3(new_n485_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n491_), .B1(new_n505_), .B2(new_n467_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT78), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(new_n507_), .A3(new_n497_), .ZN(new_n508_));
  AOI22_X1  g307(.A1(new_n499_), .A2(new_n508_), .B1(new_n493_), .B2(new_n498_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n465_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n375_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G232gat), .A2(G233gat), .ZN(new_n512_));
  XOR2_X1   g311(.A(new_n512_), .B(KEYINPUT34), .Z(new_n513_));
  INV_X1    g312(.A(KEYINPUT35), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n448_), .A2(new_n489_), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n434_), .A2(new_n478_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n513_), .A2(new_n514_), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n518_), .B(KEYINPUT69), .Z(new_n519_));
  AOI21_X1  g318(.A(KEYINPUT70), .B1(new_n517_), .B2(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n516_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n517_), .A2(KEYINPUT70), .A3(new_n519_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n515_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n517_), .A2(new_n519_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n515_), .B(KEYINPUT71), .ZN(new_n525_));
  NOR3_X1   g324(.A1(new_n516_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n523_), .A2(new_n526_), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n527_), .A2(KEYINPUT36), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G190gat), .B(G218gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G134gat), .B(G162gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n528_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n527_), .A2(KEYINPUT36), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n528_), .A2(new_n532_), .A3(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n536_), .A2(KEYINPUT37), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT37), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n538_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G231gat), .A2(G233gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n475_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(new_n435_), .ZN(new_n543_));
  XOR2_X1   g342(.A(KEYINPUT72), .B(KEYINPUT16), .Z(new_n544_));
  XNOR2_X1  g343(.A(G127gat), .B(G155gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G183gat), .B(G211gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT17), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n543_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT73), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n548_), .A2(new_n549_), .ZN(new_n553_));
  NOR3_X1   g352(.A1(new_n543_), .A2(new_n550_), .A3(new_n553_), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT74), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n540_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n511_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n560_), .A2(new_n470_), .A3(new_n370_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT38), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n366_), .A2(new_n367_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n368_), .A2(new_n371_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n374_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n341_), .B(KEYINPUT98), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n536_), .ZN(new_n568_));
  NOR3_X1   g367(.A1(new_n567_), .A2(new_n557_), .A3(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n510_), .B(KEYINPUT99), .Z(new_n570_));
  AND2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n571_), .A2(new_n370_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n562_), .B1(new_n470_), .B2(new_n572_), .ZN(G1324gat));
  INV_X1    g372(.A(new_n368_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n471_), .B1(new_n571_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT39), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n560_), .A2(new_n471_), .A3(new_n574_), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n578_), .B(KEYINPUT100), .Z(new_n579_));
  XNOR2_X1  g378(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n577_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n580_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(G1325gat));
  INV_X1    g382(.A(G15gat), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n584_), .B1(new_n571_), .B2(new_n374_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT41), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n560_), .A2(new_n584_), .A3(new_n374_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(G1326gat));
  INV_X1    g387(.A(G22gat), .ZN(new_n589_));
  INV_X1    g388(.A(new_n367_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n589_), .B1(new_n571_), .B2(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n591_), .B(KEYINPUT42), .Z(new_n592_));
  NAND3_X1  g391(.A1(new_n560_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(G1327gat));
  NOR3_X1   g393(.A1(new_n511_), .A2(new_n556_), .A3(new_n536_), .ZN(new_n595_));
  AOI21_X1  g394(.A(G29gat), .B1(new_n595_), .B2(new_n370_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT43), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n597_), .B(new_n540_), .C1(new_n565_), .C2(new_n566_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT103), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n540_), .B(KEYINPUT102), .ZN(new_n600_));
  OAI21_X1  g399(.A(KEYINPUT43), .B1(new_n567_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT103), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n375_), .A2(new_n602_), .A3(new_n597_), .A4(new_n540_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n599_), .A2(new_n601_), .A3(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n604_), .A2(new_n570_), .A3(new_n557_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT44), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n604_), .A2(KEYINPUT44), .A3(new_n570_), .A4(new_n557_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n607_), .A2(G29gat), .A3(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n596_), .B1(new_n609_), .B2(new_n370_), .ZN(G1328gat));
  NAND3_X1  g409(.A1(new_n607_), .A2(new_n574_), .A3(new_n608_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(G36gat), .ZN(new_n612_));
  INV_X1    g411(.A(G36gat), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n536_), .A2(new_n556_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n375_), .A2(new_n613_), .A3(new_n510_), .A4(new_n614_), .ZN(new_n615_));
  OR3_X1    g414(.A1(new_n615_), .A2(KEYINPUT104), .A3(new_n368_), .ZN(new_n616_));
  OAI21_X1  g415(.A(KEYINPUT104), .B1(new_n615_), .B2(new_n368_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT45), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n612_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT46), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n612_), .A2(KEYINPUT46), .A3(new_n619_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(G1329gat));
  NAND3_X1  g423(.A1(new_n607_), .A2(new_n340_), .A3(new_n608_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(G43gat), .ZN(new_n626_));
  INV_X1    g425(.A(G43gat), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n595_), .A2(new_n627_), .A3(new_n374_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(KEYINPUT105), .B(KEYINPUT47), .Z(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n630_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n626_), .A2(new_n632_), .A3(new_n628_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(G1330gat));
  AND4_X1   g433(.A1(G50gat), .A2(new_n607_), .A3(new_n590_), .A4(new_n608_), .ZN(new_n635_));
  AOI21_X1  g434(.A(G50gat), .B1(new_n595_), .B2(new_n590_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(G1331gat));
  INV_X1    g436(.A(new_n465_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n509_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n375_), .A2(new_n558_), .A3(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(G57gat), .B1(new_n641_), .B2(new_n370_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n569_), .A2(new_n640_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n643_), .A2(G57gat), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n642_), .B1(new_n644_), .B2(new_n370_), .ZN(G1332gat));
  INV_X1    g444(.A(G64gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n646_), .B1(new_n643_), .B2(new_n574_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT48), .Z(new_n648_));
  NAND3_X1  g447(.A1(new_n641_), .A2(new_n646_), .A3(new_n574_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(G1333gat));
  AOI21_X1  g449(.A(new_n334_), .B1(new_n643_), .B2(new_n374_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT49), .Z(new_n652_));
  NAND3_X1  g451(.A1(new_n641_), .A2(new_n334_), .A3(new_n374_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1334gat));
  INV_X1    g453(.A(G78gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n655_), .B1(new_n643_), .B2(new_n590_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT50), .Z(new_n657_));
  NAND3_X1  g456(.A1(new_n641_), .A2(new_n655_), .A3(new_n590_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1335gat));
  AND3_X1   g458(.A1(new_n375_), .A2(new_n614_), .A3(new_n640_), .ZN(new_n660_));
  AOI21_X1  g459(.A(G85gat), .B1(new_n660_), .B2(new_n370_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n604_), .A2(new_n557_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n662_), .A2(new_n640_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n663_), .A2(G85gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n661_), .B1(new_n664_), .B2(new_n370_), .ZN(G1336gat));
  AOI21_X1  g464(.A(G92gat), .B1(new_n660_), .B2(new_n574_), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n666_), .B(KEYINPUT106), .Z(new_n667_));
  NOR2_X1   g466(.A1(new_n368_), .A2(new_n318_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n667_), .B1(new_n663_), .B2(new_n668_), .ZN(G1337gat));
  NAND3_X1  g468(.A1(new_n662_), .A2(new_n374_), .A3(new_n640_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(G99gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n660_), .A2(new_n405_), .A3(new_n340_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g473(.A1(new_n660_), .A2(new_n406_), .A3(new_n590_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n604_), .A2(new_n557_), .A3(new_n590_), .A4(new_n640_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT52), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n676_), .A2(new_n677_), .A3(G106gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n677_), .B1(new_n676_), .B2(G106gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n675_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g480(.A1(new_n558_), .A2(new_n509_), .A3(new_n638_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT54), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT54), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n558_), .A2(new_n684_), .A3(new_n509_), .A4(new_n638_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n505_), .A2(new_n466_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n490_), .A2(new_n483_), .A3(new_n467_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(new_n498_), .A3(new_n688_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n455_), .A2(new_n460_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n508_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n507_), .B1(new_n506_), .B2(new_n497_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n689_), .B(new_n691_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT112), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n499_), .A2(new_n508_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT112), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n696_), .A2(new_n697_), .A3(new_n689_), .A4(new_n691_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n695_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n451_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT55), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT55), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n451_), .A2(new_n700_), .A3(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT109), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n449_), .B1(new_n448_), .B2(new_n387_), .ZN(new_n706_));
  AOI211_X1 g505(.A(KEYINPUT67), .B(new_n386_), .C1(new_n447_), .C2(new_n422_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n436_), .A2(new_n437_), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n706_), .A2(new_n707_), .A3(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n705_), .B1(new_n709_), .B2(new_n433_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n432_), .A2(new_n438_), .A3(new_n450_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n711_), .A2(KEYINPUT109), .A3(new_n453_), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n702_), .A2(new_n704_), .A3(new_n710_), .A4(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(KEYINPUT56), .B1(new_n713_), .B2(new_n460_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT113), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n713_), .A2(KEYINPUT56), .A3(new_n460_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n714_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  AOI211_X1 g516(.A(KEYINPUT113), .B(KEYINPUT56), .C1(new_n713_), .C2(new_n460_), .ZN(new_n718_));
  OAI211_X1 g517(.A(KEYINPUT114), .B(new_n699_), .C1(new_n717_), .C2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT58), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n716_), .A2(new_n715_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n713_), .A2(new_n460_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT56), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n722_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n718_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT114), .B1(new_n728_), .B2(new_n699_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n540_), .B1(new_n721_), .B2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT115), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n728_), .A2(KEYINPUT58), .A3(new_n699_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT115), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n733_), .B(new_n540_), .C1(new_n721_), .C2(new_n729_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n731_), .A2(new_n732_), .A3(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT116), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n639_), .A2(new_n737_), .A3(new_n691_), .ZN(new_n738_));
  OAI21_X1  g537(.A(KEYINPUT107), .B1(new_n509_), .B2(new_n690_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n714_), .B(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n740_), .B1(new_n742_), .B2(new_n716_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n696_), .A2(new_n689_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n744_), .A2(new_n462_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n536_), .B1(new_n743_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT57), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n736_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n738_), .A2(new_n739_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n725_), .A2(new_n741_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n714_), .A2(KEYINPUT110), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(new_n716_), .A3(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n745_), .B1(new_n749_), .B2(new_n752_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n753_), .A2(new_n568_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(KEYINPUT116), .A3(KEYINPUT57), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n748_), .A2(new_n755_), .ZN(new_n756_));
  XOR2_X1   g555(.A(KEYINPUT111), .B(KEYINPUT57), .Z(new_n757_));
  NAND2_X1  g556(.A1(new_n746_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n735_), .A2(new_n756_), .A3(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n686_), .B1(new_n759_), .B2(new_n557_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  AND4_X1   g560(.A1(new_n370_), .A2(new_n368_), .A3(new_n340_), .A4(new_n367_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(G113gat), .B1(new_n763_), .B2(new_n639_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT117), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n735_), .A2(new_n765_), .A3(new_n758_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n756_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n765_), .B1(new_n735_), .B2(new_n758_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n557_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n686_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT59), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n771_), .A2(new_n772_), .A3(new_n762_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n763_), .A2(new_n772_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n773_), .A2(new_n774_), .A3(new_n509_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n764_), .B1(new_n775_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g575(.A(G120gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n777_), .B1(new_n638_), .B2(KEYINPUT60), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n763_), .B(new_n778_), .C1(KEYINPUT60), .C2(new_n777_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n773_), .A2(new_n774_), .A3(new_n638_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n779_), .B1(new_n780_), .B2(new_n777_), .ZN(G1341gat));
  AOI21_X1  g580(.A(G127gat), .B1(new_n763_), .B2(new_n556_), .ZN(new_n782_));
  INV_X1    g581(.A(G127gat), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n773_), .A2(new_n774_), .A3(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n782_), .B1(new_n784_), .B2(new_n556_), .ZN(G1342gat));
  AOI21_X1  g584(.A(G134gat), .B1(new_n763_), .B2(new_n568_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n773_), .A2(new_n774_), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n537_), .A2(new_n539_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(KEYINPUT118), .B(G134gat), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n786_), .B1(new_n787_), .B2(new_n790_), .ZN(G1343gat));
  INV_X1    g590(.A(KEYINPUT119), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n759_), .A2(new_n557_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n369_), .B1(new_n793_), .B2(new_n770_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n574_), .A2(new_n374_), .A3(new_n367_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n792_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n795_), .ZN(new_n797_));
  NOR4_X1   g596(.A1(new_n760_), .A2(KEYINPUT119), .A3(new_n369_), .A4(new_n797_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n796_), .A2(new_n798_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n799_), .A2(new_n509_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(new_n203_), .ZN(G1344gat));
  NOR2_X1   g600(.A1(new_n799_), .A2(new_n638_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(new_n204_), .ZN(G1345gat));
  OAI21_X1  g602(.A(new_n556_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT120), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT120), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n806_), .B(new_n556_), .C1(new_n796_), .C2(new_n798_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(KEYINPUT61), .B(G155gat), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n805_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n809_), .A2(new_n810_), .ZN(G1346gat));
  INV_X1    g610(.A(G162gat), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n799_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n600_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n568_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n815_));
  AOI22_X1  g614(.A1(new_n813_), .A2(new_n814_), .B1(new_n812_), .B2(new_n815_), .ZN(G1347gat));
  NOR4_X1   g615(.A1(new_n368_), .A2(new_n370_), .A3(new_n373_), .A4(new_n590_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n771_), .A2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(G169gat), .B1(new_n818_), .B2(new_n509_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT121), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT121), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n821_), .B(G169gat), .C1(new_n818_), .C2(new_n509_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n820_), .A2(KEYINPUT62), .A3(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n818_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n824_), .A2(new_n639_), .A3(new_n290_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT62), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n819_), .A2(KEYINPUT121), .A3(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n823_), .A2(new_n825_), .A3(new_n827_), .ZN(G1348gat));
  AND2_X1   g627(.A1(new_n761_), .A2(new_n817_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n829_), .A2(G176gat), .A3(new_n465_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(KEYINPUT122), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n824_), .A2(new_n465_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(new_n289_), .B2(new_n832_), .ZN(G1349gat));
  INV_X1    g632(.A(new_n279_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n824_), .A2(new_n556_), .A3(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT123), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n829_), .A2(new_n556_), .ZN(new_n837_));
  OR2_X1    g636(.A1(new_n837_), .A2(G183gat), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT123), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n824_), .A2(new_n839_), .A3(new_n556_), .A4(new_n834_), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n836_), .A2(new_n838_), .A3(new_n840_), .ZN(G1350gat));
  NAND3_X1  g640(.A1(new_n824_), .A2(new_n568_), .A3(new_n280_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT124), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n824_), .A2(new_n540_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(G190gat), .ZN(new_n845_));
  INV_X1    g644(.A(G190gat), .ZN(new_n846_));
  AOI211_X1 g645(.A(KEYINPUT124), .B(new_n846_), .C1(new_n824_), .C2(new_n540_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n842_), .B1(new_n845_), .B2(new_n847_), .ZN(G1351gat));
  NAND2_X1  g647(.A1(new_n371_), .A2(new_n373_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n849_), .A2(KEYINPUT125), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n760_), .A2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n368_), .B1(new_n849_), .B2(KEYINPUT125), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(new_n509_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(KEYINPUT126), .B(G197gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n854_), .B2(new_n857_), .ZN(G1352gat));
  NAND2_X1  g657(.A1(new_n457_), .A2(KEYINPUT127), .ZN(new_n859_));
  XOR2_X1   g658(.A(KEYINPUT127), .B(G204gat), .Z(new_n860_));
  NOR2_X1   g659(.A1(new_n853_), .A2(new_n638_), .ZN(new_n861_));
  MUX2_X1   g660(.A(new_n859_), .B(new_n860_), .S(new_n861_), .Z(G1353gat));
  INV_X1    g661(.A(new_n853_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n556_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n865_));
  AND2_X1   g664(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n864_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n867_), .B1(new_n864_), .B2(new_n865_), .ZN(G1354gat));
  AND3_X1   g667(.A1(new_n863_), .A2(G218gat), .A3(new_n540_), .ZN(new_n869_));
  AOI21_X1  g668(.A(G218gat), .B1(new_n863_), .B2(new_n568_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1355gat));
endmodule


