//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 1 0 0 0 1 1 0 1 0 0 0 0 1 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n925_, new_n927_, new_n928_, new_n929_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT23), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G183gat), .A3(G190gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(G169gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT24), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT79), .ZN(new_n215_));
  NOR3_X1   g014(.A1(new_n215_), .A2(G169gat), .A3(G176gat), .ZN(new_n216_));
  INV_X1    g015(.A(G169gat), .ZN(new_n217_));
  INV_X1    g016(.A(G176gat), .ZN(new_n218_));
  AOI21_X1  g017(.A(KEYINPUT79), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n214_), .B1(new_n216_), .B2(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT80), .B1(new_n203_), .B2(new_n205_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT80), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n222_), .B1(new_n202_), .B2(KEYINPUT23), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n220_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G190gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT26), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT26), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(G190gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT88), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT25), .B(G183gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n226_), .A2(new_n228_), .A3(KEYINPUT88), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n216_), .A2(new_n219_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n214_), .B1(G169gat), .B2(G176gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n234_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT89), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n224_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n234_), .A2(new_n237_), .A3(KEYINPUT89), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n213_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(G211gat), .B(G218gat), .Z(new_n243_));
  INV_X1    g042(.A(KEYINPUT21), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G197gat), .B(G204gat), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n243_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n245_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT21), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n247_), .A2(new_n243_), .A3(KEYINPUT21), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT90), .B1(new_n242_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT90), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n234_), .A2(new_n237_), .A3(KEYINPUT89), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT89), .B1(new_n234_), .B2(new_n237_), .ZN(new_n256_));
  NOR3_X1   g055(.A1(new_n255_), .A2(new_n256_), .A3(new_n224_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n254_), .B(new_n251_), .C1(new_n257_), .C2(new_n213_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n232_), .A2(new_n226_), .A3(new_n228_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n237_), .A2(new_n206_), .A3(new_n220_), .A4(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n208_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(new_n211_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT20), .B1(new_n263_), .B2(new_n251_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n253_), .A2(new_n258_), .A3(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G226gat), .A2(G233gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT19), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G8gat), .B(G36gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G64gat), .B(G92gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n240_), .A2(new_n241_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n276_), .A2(new_n252_), .A3(new_n212_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n268_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT20), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n279_), .B1(new_n263_), .B2(new_n251_), .ZN(new_n280_));
  AND3_X1   g079(.A1(new_n277_), .A2(new_n278_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n269_), .A2(new_n275_), .A3(new_n282_), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n283_), .A2(KEYINPUT27), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n277_), .A2(new_n280_), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n285_), .A2(new_n278_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n251_), .B1(new_n257_), .B2(new_n213_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n264_), .B1(new_n287_), .B2(KEYINPUT90), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT95), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n288_), .A2(new_n289_), .A3(new_n278_), .A4(new_n258_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n253_), .A2(new_n258_), .A3(new_n278_), .A4(new_n265_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT95), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n286_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n274_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n278_), .B1(new_n288_), .B2(new_n258_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n274_), .B1(new_n295_), .B2(new_n281_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(new_n283_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT27), .ZN(new_n298_));
  AOI22_X1  g097(.A1(new_n284_), .A2(new_n294_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT87), .ZN(new_n301_));
  INV_X1    g100(.A(G228gat), .ZN(new_n302_));
  INV_X1    g101(.A(G233gat), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n251_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT3), .ZN(new_n305_));
  INV_X1    g104(.A(G141gat), .ZN(new_n306_));
  INV_X1    g105(.A(G148gat), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G141gat), .A2(G148gat), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT2), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n308_), .A2(new_n311_), .A3(new_n312_), .A4(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(G155gat), .B(G162gat), .Z(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT82), .ZN(new_n317_));
  AND2_X1   g116(.A1(G141gat), .A2(G148gat), .ZN(new_n318_));
  NOR2_X1   g117(.A1(G141gat), .A2(G148gat), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G155gat), .B(G162gat), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n320_), .B(new_n321_), .C1(new_n322_), .C2(KEYINPUT1), .ZN(new_n323_));
  AND3_X1   g122(.A1(new_n316_), .A2(new_n317_), .A3(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n317_), .B1(new_n316_), .B2(new_n323_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT83), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n326_), .A2(new_n327_), .A3(KEYINPUT29), .ZN(new_n328_));
  INV_X1    g127(.A(new_n313_), .ZN(new_n329_));
  NOR3_X1   g128(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n312_), .ZN(new_n332_));
  AOI21_X1  g131(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n322_), .B1(new_n331_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n306_), .A2(new_n307_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n336_), .A2(new_n321_), .A3(new_n309_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT1), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n337_), .B1(new_n315_), .B2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT82), .B1(new_n335_), .B2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n316_), .A2(new_n317_), .A3(new_n323_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(KEYINPUT29), .A3(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT83), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n304_), .B1(new_n328_), .B2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT29), .B1(new_n335_), .B2(new_n339_), .ZN(new_n345_));
  AOI211_X1 g144(.A(new_n302_), .B(new_n303_), .C1(new_n251_), .C2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G78gat), .B(G106gat), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n348_), .B(KEYINPUT84), .Z(new_n349_));
  XOR2_X1   g148(.A(new_n349_), .B(KEYINPUT85), .Z(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT28), .B1(new_n326_), .B2(KEYINPUT29), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n340_), .A2(new_n341_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT28), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT29), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G22gat), .B(G50gat), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n351_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n356_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n353_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n359_));
  AOI211_X1 g158(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n340_), .C2(new_n341_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n358_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  AOI22_X1  g160(.A1(new_n347_), .A2(new_n350_), .B1(new_n357_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT86), .ZN(new_n363_));
  INV_X1    g162(.A(new_n304_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n327_), .B1(new_n326_), .B2(KEYINPUT29), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n342_), .A2(KEYINPUT83), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n364_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n346_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n350_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n363_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n363_), .B(new_n370_), .C1(new_n344_), .C2(new_n346_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n362_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n347_), .A2(new_n349_), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n344_), .A2(new_n346_), .A3(new_n370_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n357_), .B(new_n361_), .C1(new_n375_), .C2(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n301_), .B1(new_n374_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n374_), .A2(new_n377_), .A3(new_n301_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT81), .ZN(new_n382_));
  INV_X1    g181(.A(G134gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(G127gat), .ZN(new_n384_));
  INV_X1    g183(.A(G127gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(G134gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(G120gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(G113gat), .ZN(new_n389_));
  INV_X1    g188(.A(G113gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(G120gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n382_), .B1(new_n387_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n387_), .A2(new_n392_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n384_), .A2(new_n386_), .A3(new_n389_), .A4(new_n391_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n393_), .B1(new_n396_), .B2(new_n382_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n340_), .A2(new_n341_), .A3(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT92), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n396_), .A2(new_n316_), .A3(new_n323_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT92), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n340_), .A2(new_n397_), .A3(new_n401_), .A4(new_n341_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n399_), .A2(KEYINPUT4), .A3(new_n400_), .A4(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT93), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n402_), .A2(new_n400_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT93), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n405_), .A2(new_n406_), .A3(KEYINPUT4), .A4(new_n399_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n404_), .A2(new_n407_), .ZN(new_n408_));
  OR2_X1    g207(.A1(new_n398_), .A2(KEYINPUT4), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G225gat), .A2(G233gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n408_), .A2(new_n413_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n405_), .A2(new_n399_), .A3(new_n410_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G1gat), .B(G29gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(G85gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT0), .B(G57gat), .ZN(new_n419_));
  XOR2_X1   g218(.A(new_n418_), .B(new_n419_), .Z(new_n420_));
  NAND3_X1  g219(.A1(new_n414_), .A2(new_n416_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n420_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n412_), .B1(new_n404_), .B2(new_n407_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n422_), .B1(new_n423_), .B2(new_n415_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n421_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G227gat), .A2(G233gat), .ZN(new_n427_));
  INV_X1    g226(.A(G15gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT30), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n263_), .B(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(new_n397_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G71gat), .B(G99gat), .ZN(new_n433_));
  INV_X1    g232(.A(G43gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT31), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n432_), .B(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n426_), .A2(new_n437_), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n300_), .A2(new_n381_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT96), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT94), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT33), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n414_), .A2(new_n416_), .A3(new_n420_), .A4(new_n443_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n409_), .A2(new_n410_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n408_), .A2(new_n445_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n405_), .A2(new_n399_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n420_), .B1(new_n447_), .B2(new_n411_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  AND4_X1   g248(.A1(new_n444_), .A2(new_n283_), .A3(new_n296_), .A4(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n415_), .B1(new_n408_), .B2(new_n413_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n443_), .B1(new_n451_), .B2(new_n420_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n275_), .A2(KEYINPUT32), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n293_), .A2(new_n454_), .ZN(new_n455_));
  AOI211_X1 g254(.A(new_n454_), .B(new_n281_), .C1(new_n268_), .C2(new_n266_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n456_), .B1(new_n421_), .B2(new_n424_), .ZN(new_n457_));
  AOI22_X1  g256(.A1(new_n450_), .A2(new_n453_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n440_), .B1(new_n458_), .B2(new_n381_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n367_), .A2(new_n368_), .A3(new_n350_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n361_), .A2(new_n357_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT86), .B1(new_n347_), .B2(new_n350_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n462_), .B1(new_n463_), .B2(new_n372_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n349_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n369_), .A2(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n461_), .B1(new_n466_), .B2(new_n460_), .ZN(new_n467_));
  NOR3_X1   g266(.A1(new_n464_), .A2(KEYINPUT87), .A3(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n468_), .A2(new_n378_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n296_), .A2(new_n449_), .A3(new_n283_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n444_), .ZN(new_n471_));
  NOR3_X1   g270(.A1(new_n470_), .A2(new_n471_), .A3(new_n452_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n456_), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n425_), .A2(new_n455_), .A3(new_n473_), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n469_), .B(KEYINPUT96), .C1(new_n472_), .C2(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n425_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(new_n299_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n459_), .A2(new_n475_), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n437_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n439_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G29gat), .B(G36gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G43gat), .B(G50gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT15), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G15gat), .B(G22gat), .ZN(new_n486_));
  INV_X1    g285(.A(G1gat), .ZN(new_n487_));
  INV_X1    g286(.A(G8gat), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT14), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n486_), .A2(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G1gat), .B(G8gat), .Z(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n485_), .A2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT77), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G229gat), .A2(G233gat), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  XOR2_X1   g295(.A(new_n483_), .B(KEYINPUT76), .Z(new_n497_));
  AOI21_X1  g296(.A(new_n496_), .B1(new_n497_), .B2(new_n492_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n494_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n497_), .B(new_n492_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n496_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G113gat), .B(G141gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G169gat), .B(G197gat), .ZN(new_n503_));
  XOR2_X1   g302(.A(new_n502_), .B(new_n503_), .Z(new_n504_));
  AND3_X1   g303(.A1(new_n499_), .A2(new_n501_), .A3(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n504_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT78), .ZN(new_n507_));
  OR3_X1    g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n507_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT70), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G85gat), .B(G92gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT64), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT8), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G99gat), .A2(G106gat), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT6), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  OR3_X1    g317(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n514_), .B(new_n515_), .C1(new_n518_), .C2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT64), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n513_), .B(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n519_), .A2(KEYINPUT65), .A3(new_n520_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT65), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n518_), .B1(new_n526_), .B2(new_n521_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n524_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n522_), .B1(new_n528_), .B2(new_n515_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT9), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n513_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n518_), .ZN(new_n532_));
  XOR2_X1   g331(.A(KEYINPUT10), .B(G99gat), .Z(new_n533_));
  INV_X1    g332(.A(G106gat), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n530_), .A2(G85gat), .A3(G92gat), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n531_), .A2(new_n532_), .A3(new_n535_), .A4(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT66), .B(G71gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(G78gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G57gat), .B(G64gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT11), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n540_), .A2(KEYINPUT11), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n539_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(G78gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n538_), .B(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n541_), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n544_), .A2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n529_), .A2(new_n537_), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G230gat), .A2(G233gat), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(KEYINPUT69), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(KEYINPUT69), .B1(new_n549_), .B2(new_n550_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n544_), .A2(new_n547_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT68), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT12), .ZN(new_n557_));
  INV_X1    g356(.A(new_n537_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n529_), .A2(KEYINPUT67), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT67), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n560_), .B(new_n522_), .C1(new_n528_), .C2(new_n515_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n558_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n548_), .B1(new_n529_), .B2(new_n537_), .ZN(new_n563_));
  OAI22_X1  g362(.A1(new_n557_), .A2(new_n562_), .B1(new_n563_), .B2(KEYINPUT12), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n512_), .B1(new_n554_), .B2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n563_), .A2(KEYINPUT12), .ZN(new_n566_));
  INV_X1    g365(.A(new_n562_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT68), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n555_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT12), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n566_), .B1(new_n567_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n553_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(new_n551_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n572_), .A2(KEYINPUT70), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n550_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n549_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n576_), .B1(new_n577_), .B2(new_n563_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n565_), .A2(new_n575_), .A3(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(G176gat), .B(G204gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT72), .ZN(new_n581_));
  XOR2_X1   g380(.A(KEYINPUT71), .B(KEYINPUT5), .Z(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G120gat), .B(G148gat), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n583_), .B(new_n584_), .Z(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n579_), .A2(new_n586_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n565_), .A2(new_n575_), .A3(new_n578_), .A4(new_n585_), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n587_), .A2(KEYINPUT73), .A3(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(KEYINPUT73), .B1(new_n587_), .B2(new_n588_), .ZN(new_n590_));
  OAI21_X1  g389(.A(KEYINPUT13), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n587_), .A2(new_n588_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT73), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT13), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n587_), .A2(KEYINPUT73), .A3(new_n588_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n594_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n511_), .B1(new_n591_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n480_), .A2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G190gat), .B(G218gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G134gat), .B(G162gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n603_), .B(KEYINPUT36), .Z(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n529_), .A2(new_n483_), .A3(new_n537_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(G232gat), .A2(G233gat), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n607_), .B(KEYINPUT34), .Z(new_n608_));
  XOR2_X1   g407(.A(KEYINPUT74), .B(KEYINPUT35), .Z(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n606_), .B(new_n610_), .C1(new_n562_), .C2(new_n485_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n608_), .A2(new_n609_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n605_), .B1(new_n613_), .B2(KEYINPUT75), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n614_), .B1(KEYINPUT75), .B2(new_n613_), .ZN(new_n615_));
  OR3_X1    g414(.A1(new_n613_), .A2(KEYINPUT36), .A3(new_n603_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT37), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n613_), .A2(new_n604_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n616_), .A2(KEYINPUT37), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(G127gat), .B(G155gat), .Z(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT16), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G183gat), .B(G211gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT17), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(G231gat), .A2(G233gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n492_), .B(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n628_), .B1(new_n548_), .B2(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n631_), .B1(new_n548_), .B2(new_n630_), .ZN(new_n632_));
  AOI211_X1 g431(.A(new_n627_), .B(new_n626_), .C1(new_n556_), .C2(new_n630_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n633_), .B1(new_n556_), .B2(new_n630_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n622_), .A2(new_n636_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n600_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n638_), .A2(new_n487_), .A3(new_n425_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT38), .ZN(new_n640_));
  INV_X1    g439(.A(new_n617_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n480_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n642_), .A2(new_n598_), .A3(new_n635_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT97), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n487_), .B1(new_n644_), .B2(new_n425_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT98), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n645_), .A2(new_n646_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n640_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT99), .ZN(G1324gat));
  NAND3_X1  g449(.A1(new_n638_), .A2(new_n488_), .A3(new_n300_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n643_), .A2(new_n299_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n488_), .B1(new_n652_), .B2(KEYINPUT100), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n653_), .B1(KEYINPUT100), .B2(new_n652_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n654_), .A2(KEYINPUT39), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(KEYINPUT39), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n651_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n657_), .B(new_n659_), .ZN(G1325gat));
  AOI21_X1  g459(.A(new_n428_), .B1(new_n644_), .B2(new_n437_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT41), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n638_), .A2(new_n428_), .A3(new_n437_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1326gat));
  INV_X1    g463(.A(G22gat), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n665_), .B1(new_n644_), .B2(new_n381_), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n666_), .B(KEYINPUT42), .Z(new_n667_));
  NAND3_X1  g466(.A1(new_n638_), .A2(new_n665_), .A3(new_n381_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1327gat));
  NOR2_X1   g468(.A1(new_n617_), .A2(new_n635_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n600_), .A2(new_n670_), .ZN(new_n671_));
  OR3_X1    g470(.A1(new_n671_), .A2(G29gat), .A3(new_n426_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n622_), .ZN(new_n673_));
  OAI21_X1  g472(.A(KEYINPUT43), .B1(new_n480_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n469_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n676_));
  AOI22_X1  g475(.A1(new_n676_), .A2(new_n440_), .B1(new_n476_), .B2(new_n299_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n437_), .B1(new_n677_), .B2(new_n475_), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n675_), .B(new_n622_), .C1(new_n678_), .C2(new_n439_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n674_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n598_), .A2(new_n636_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT44), .B1(new_n680_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684_));
  AOI211_X1 g483(.A(new_n684_), .B(new_n681_), .C1(new_n674_), .C2(new_n679_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n686_), .A2(KEYINPUT102), .A3(new_n425_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(G29gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT102), .B1(new_n686_), .B2(new_n425_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n672_), .B1(new_n688_), .B2(new_n689_), .ZN(G1328gat));
  NAND2_X1  g489(.A1(new_n680_), .A2(new_n682_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(new_n684_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n680_), .A2(KEYINPUT44), .A3(new_n682_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n692_), .A2(new_n693_), .A3(new_n300_), .A4(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(G36gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n693_), .B1(new_n686_), .B2(new_n300_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT104), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n692_), .A2(new_n300_), .A3(new_n694_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT103), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n700_), .A2(new_n701_), .A3(G36gat), .A4(new_n695_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n698_), .A2(new_n702_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n671_), .A2(G36gat), .A3(new_n299_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT45), .Z(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n703_), .A2(KEYINPUT46), .A3(new_n705_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1329gat));
  NAND3_X1  g509(.A1(new_n686_), .A2(G43gat), .A3(new_n437_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n434_), .B1(new_n671_), .B2(new_n479_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n713_), .B(new_n714_), .ZN(G1330gat));
  OR3_X1    g514(.A1(new_n671_), .A2(G50gat), .A3(new_n469_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT106), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n686_), .A2(new_n717_), .A3(new_n381_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(G50gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n717_), .B1(new_n686_), .B2(new_n381_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n716_), .B1(new_n719_), .B2(new_n720_), .ZN(G1331gat));
  NAND2_X1  g520(.A1(new_n591_), .A2(new_n597_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n642_), .A2(new_n511_), .A3(new_n723_), .A4(new_n635_), .ZN(new_n724_));
  OAI21_X1  g523(.A(G57gat), .B1(new_n724_), .B2(new_n426_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n480_), .A2(new_n510_), .A3(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(new_n637_), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n426_), .A2(G57gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n725_), .B1(new_n727_), .B2(new_n728_), .ZN(G1332gat));
  OAI21_X1  g528(.A(G64gat), .B1(new_n724_), .B2(new_n299_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT48), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n299_), .A2(G64gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n727_), .B2(new_n732_), .ZN(G1333gat));
  OAI21_X1  g532(.A(G71gat), .B1(new_n724_), .B2(new_n479_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n734_), .A2(KEYINPUT49), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n734_), .A2(KEYINPUT49), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n479_), .A2(G71gat), .ZN(new_n737_));
  OAI22_X1  g536(.A1(new_n735_), .A2(new_n736_), .B1(new_n727_), .B2(new_n737_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT107), .Z(G1334gat));
  OAI21_X1  g538(.A(G78gat), .B1(new_n724_), .B2(new_n469_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT50), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n381_), .A2(new_n545_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n741_), .B1(new_n727_), .B2(new_n742_), .ZN(G1335gat));
  NAND2_X1  g542(.A1(new_n726_), .A2(new_n670_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(G85gat), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n745_), .A2(new_n746_), .A3(new_n425_), .ZN(new_n747_));
  AND4_X1   g546(.A1(new_n511_), .A2(new_n680_), .A3(new_n723_), .A4(new_n636_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n748_), .A2(new_n425_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n747_), .B1(new_n749_), .B2(new_n746_), .ZN(G1336gat));
  INV_X1    g549(.A(G92gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n745_), .A2(new_n751_), .A3(new_n300_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n748_), .A2(new_n300_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n752_), .B1(new_n753_), .B2(new_n751_), .ZN(G1337gat));
  INV_X1    g553(.A(G99gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n748_), .B2(new_n437_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n756_), .A2(KEYINPUT108), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n756_), .A2(KEYINPUT108), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n437_), .A2(new_n533_), .ZN(new_n759_));
  OAI22_X1  g558(.A1(new_n757_), .A2(new_n758_), .B1(new_n744_), .B2(new_n759_), .ZN(new_n760_));
  AND2_X1   g559(.A1(KEYINPUT109), .A2(KEYINPUT51), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n760_), .B(new_n761_), .ZN(G1338gat));
  AOI21_X1  g561(.A(new_n534_), .B1(new_n748_), .B2(new_n381_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n763_), .A2(new_n764_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n381_), .A2(new_n534_), .ZN(new_n767_));
  OAI22_X1  g566(.A1(new_n765_), .A2(new_n766_), .B1(new_n744_), .B2(new_n767_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g568(.A1(new_n300_), .A2(new_n381_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n770_), .A2(new_n425_), .A3(new_n437_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n508_), .A2(new_n509_), .A3(new_n635_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n508_), .A2(new_n509_), .A3(KEYINPUT110), .A4(new_n635_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n589_), .A2(new_n590_), .A3(KEYINPUT13), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n595_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n779_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n722_), .A2(KEYINPUT111), .A3(new_n779_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n622_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n773_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  AOI211_X1 g587(.A(new_n783_), .B(new_n778_), .C1(new_n591_), .C2(new_n597_), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT111), .B1(new_n722_), .B2(new_n779_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n673_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n791_), .A2(KEYINPUT113), .A3(KEYINPUT54), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n787_), .B(new_n673_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT112), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n784_), .A2(new_n785_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n795_), .A2(new_n796_), .A3(new_n787_), .A4(new_n673_), .ZN(new_n797_));
  AOI22_X1  g596(.A1(new_n788_), .A2(new_n792_), .B1(new_n794_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n554_), .A2(new_n564_), .A3(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n550_), .B1(new_n572_), .B2(new_n549_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n565_), .A2(new_n575_), .A3(new_n799_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n585_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT56), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n588_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  AOI211_X1 g605(.A(KEYINPUT56), .B(new_n585_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n806_), .A2(new_n511_), .A3(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n504_), .B1(new_n500_), .B2(new_n495_), .ZN(new_n809_));
  OR2_X1    g608(.A1(new_n809_), .A2(KEYINPUT114), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(KEYINPUT114), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n495_), .B1(new_n497_), .B2(new_n492_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n494_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n810_), .A2(new_n811_), .A3(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n505_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n617_), .B1(new_n808_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n588_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n802_), .A2(new_n803_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n586_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n821_), .B1(new_n823_), .B2(KEYINPUT56), .ZN(new_n824_));
  INV_X1    g623(.A(new_n816_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n807_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n824_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(KEYINPUT115), .A2(KEYINPUT58), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n828_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n824_), .A2(new_n830_), .A3(new_n825_), .A4(new_n826_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n829_), .A2(new_n622_), .A3(new_n831_), .ZN(new_n832_));
  OAI211_X1 g631(.A(KEYINPUT57), .B(new_n617_), .C1(new_n808_), .C2(new_n817_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n820_), .A2(new_n832_), .A3(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n636_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n772_), .B1(new_n798_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n788_), .A2(new_n792_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n794_), .A2(new_n797_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT116), .B1(new_n834_), .B2(new_n636_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n834_), .A2(KEYINPUT116), .A3(new_n636_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n840_), .A2(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n771_), .A2(KEYINPUT59), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n837_), .A2(KEYINPUT59), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n390_), .B1(new_n847_), .B2(new_n510_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n837_), .A2(G113gat), .A3(new_n511_), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT117), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n834_), .A2(KEYINPUT116), .A3(new_n636_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n851_), .A2(new_n841_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n846_), .B1(new_n798_), .B2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n771_), .B1(new_n840_), .B2(new_n835_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n853_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(G113gat), .B1(new_n856_), .B2(new_n511_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n858_));
  INV_X1    g657(.A(new_n849_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n857_), .A2(new_n858_), .A3(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n850_), .A2(new_n860_), .ZN(G1340gat));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n388_), .B1(new_n847_), .B2(new_n723_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n722_), .A2(KEYINPUT60), .ZN(new_n864_));
  MUX2_X1   g663(.A(KEYINPUT60), .B(new_n864_), .S(new_n388_), .Z(new_n865_));
  NAND2_X1  g664(.A1(new_n854_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n862_), .B1(new_n863_), .B2(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(G120gat), .B1(new_n856_), .B2(new_n722_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n869_), .A2(KEYINPUT118), .A3(new_n866_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n870_), .ZN(G1341gat));
  OAI21_X1  g670(.A(G127gat), .B1(new_n856_), .B2(new_n636_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n854_), .A2(new_n385_), .A3(new_n635_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(G1342gat));
  AOI21_X1  g673(.A(G134gat), .B1(new_n854_), .B2(new_n641_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n383_), .A2(KEYINPUT119), .ZN(new_n876_));
  OR2_X1    g675(.A1(new_n383_), .A2(KEYINPUT119), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n673_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(KEYINPUT120), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n875_), .B1(new_n847_), .B2(new_n879_), .ZN(G1343gat));
  NOR3_X1   g679(.A1(new_n300_), .A2(new_n469_), .A3(new_n426_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n479_), .B(new_n881_), .C1(new_n798_), .C2(new_n836_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n511_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(new_n306_), .ZN(G1344gat));
  NOR2_X1   g683(.A1(new_n882_), .A2(new_n722_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT121), .B(G148gat), .ZN(new_n886_));
  XOR2_X1   g685(.A(new_n885_), .B(new_n886_), .Z(G1345gat));
  OR3_X1    g686(.A1(new_n882_), .A2(KEYINPUT122), .A3(new_n636_), .ZN(new_n888_));
  OAI21_X1  g687(.A(KEYINPUT122), .B1(new_n882_), .B2(new_n636_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(KEYINPUT61), .B(G155gat), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n888_), .A2(new_n889_), .A3(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1346gat));
  OAI21_X1  g692(.A(G162gat), .B1(new_n882_), .B2(new_n673_), .ZN(new_n894_));
  OR2_X1    g693(.A1(new_n617_), .A2(G162gat), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n882_), .B2(new_n895_), .ZN(G1347gat));
  OR2_X1    g695(.A1(new_n299_), .A2(new_n438_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n381_), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n510_), .B(new_n898_), .C1(new_n798_), .C2(new_n852_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(G169gat), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(KEYINPUT62), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(KEYINPUT124), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT124), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n900_), .A2(new_n903_), .A3(KEYINPUT62), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n905_), .B1(new_n900_), .B2(KEYINPUT62), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n899_), .A2(KEYINPUT123), .A3(new_n907_), .A4(G169gat), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n902_), .A2(new_n904_), .A3(new_n906_), .A4(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n898_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n910_), .B1(new_n840_), .B2(new_n844_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(KEYINPUT22), .B(G169gat), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n911_), .A2(new_n510_), .A3(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n909_), .A2(new_n913_), .ZN(G1348gat));
  AOI21_X1  g713(.A(G176gat), .B1(new_n911_), .B2(new_n723_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n798_), .A2(new_n836_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(new_n910_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n722_), .A2(new_n218_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n915_), .B1(new_n917_), .B2(new_n918_), .ZN(G1349gat));
  AOI21_X1  g718(.A(G183gat), .B1(new_n917_), .B2(new_n635_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n636_), .A2(new_n232_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n920_), .B1(new_n911_), .B2(new_n921_), .ZN(G1350gat));
  NAND4_X1  g721(.A1(new_n911_), .A2(new_n231_), .A3(new_n233_), .A4(new_n641_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n911_), .A2(new_n622_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n923_), .B1(new_n925_), .B2(new_n225_), .ZN(G1351gat));
  NOR2_X1   g725(.A1(new_n916_), .A2(new_n437_), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n469_), .A2(new_n299_), .A3(new_n425_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n927_), .A2(new_n510_), .A3(new_n928_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g729(.A1(new_n927_), .A2(new_n723_), .A3(new_n928_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g731(.A1(new_n927_), .A2(new_n928_), .ZN(new_n933_));
  NOR3_X1   g732(.A1(KEYINPUT125), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n934_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n635_), .A2(new_n935_), .ZN(new_n936_));
  OAI21_X1  g735(.A(KEYINPUT125), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n937_));
  XOR2_X1   g736(.A(new_n937_), .B(KEYINPUT126), .Z(new_n938_));
  INV_X1    g737(.A(new_n938_), .ZN(new_n939_));
  OR3_X1    g738(.A1(new_n933_), .A2(new_n936_), .A3(new_n939_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n933_), .B2(new_n936_), .ZN(new_n941_));
  AND2_X1   g740(.A1(new_n940_), .A2(new_n941_), .ZN(G1354gat));
  INV_X1    g741(.A(G218gat), .ZN(new_n943_));
  NOR3_X1   g742(.A1(new_n933_), .A2(new_n943_), .A3(new_n673_), .ZN(new_n944_));
  AND3_X1   g743(.A1(new_n927_), .A2(new_n641_), .A3(new_n928_), .ZN(new_n945_));
  AOI21_X1  g744(.A(G218gat), .B1(new_n945_), .B2(KEYINPUT127), .ZN(new_n946_));
  INV_X1    g745(.A(KEYINPUT127), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n947_), .B1(new_n933_), .B2(new_n617_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n944_), .B1(new_n946_), .B2(new_n948_), .ZN(G1355gat));
endmodule


