//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n785_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n932_, new_n934_, new_n935_,
    new_n936_, new_n938_, new_n939_, new_n940_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n962_, new_n963_, new_n964_;
  INV_X1    g000(.A(KEYINPUT78), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT15), .ZN(new_n203_));
  XOR2_X1   g002(.A(G29gat), .B(G36gat), .Z(new_n204_));
  XNOR2_X1  g003(.A(G43gat), .B(G50gat), .ZN(new_n205_));
  OR2_X1    g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n205_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n208_));
  AND3_X1   g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n208_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n203_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n206_), .A2(new_n207_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n208_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n206_), .A2(new_n208_), .A3(new_n207_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(KEYINPUT15), .A3(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G85gat), .A2(G92gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G85gat), .A2(G92gat), .ZN(new_n219_));
  NOR3_X1   g018(.A1(new_n218_), .A2(new_n219_), .A3(KEYINPUT67), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G99gat), .A2(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT6), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT6), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(G99gat), .A3(G106gat), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT7), .ZN(new_n226_));
  INV_X1    g025(.A(G99gat), .ZN(new_n227_));
  INV_X1    g026(.A(G106gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n220_), .B1(new_n225_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT8), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n222_), .A2(new_n224_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n234_), .A2(new_n230_), .A3(new_n229_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT8), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n236_), .A3(new_n220_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n233_), .A2(new_n237_), .ZN(new_n238_));
  OR2_X1    g037(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n228_), .A3(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT64), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT64), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n239_), .A2(new_n243_), .A3(new_n228_), .A4(new_n240_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n225_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n245_));
  AND2_X1   g044(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n246_));
  NOR2_X1   g045(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n217_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT66), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n250_), .B(new_n217_), .C1(new_n246_), .C2(new_n247_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n219_), .B1(new_n218_), .B2(KEYINPUT9), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n249_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n245_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n238_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n211_), .A2(new_n216_), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n214_), .A2(new_n215_), .ZN(new_n257_));
  AOI22_X1  g056(.A1(new_n233_), .A2(new_n237_), .B1(new_n245_), .B2(new_n253_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT35), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G232gat), .A2(G233gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT34), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n257_), .A2(new_n258_), .B1(new_n259_), .B2(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n259_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n256_), .A2(new_n263_), .A3(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT76), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n256_), .A2(new_n263_), .A3(KEYINPUT76), .A4(new_n265_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT75), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n256_), .A2(new_n270_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n211_), .A2(new_n216_), .A3(new_n255_), .A4(KEYINPUT75), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(new_n272_), .A3(new_n263_), .ZN(new_n273_));
  AOI22_X1  g072(.A1(new_n268_), .A2(new_n269_), .B1(new_n273_), .B2(new_n264_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G190gat), .B(G218gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G134gat), .B(G162gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n277_), .B(KEYINPUT36), .Z(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n202_), .B1(new_n274_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n268_), .A2(new_n269_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n273_), .A2(new_n264_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n283_), .A2(KEYINPUT78), .A3(new_n278_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n277_), .A2(KEYINPUT36), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n274_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n280_), .A2(new_n284_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT37), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n288_), .B1(new_n274_), .B2(new_n285_), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n278_), .B(KEYINPUT77), .Z(new_n290_));
  NAND2_X1  g089(.A1(new_n283_), .A2(new_n290_), .ZN(new_n291_));
  AOI22_X1  g090(.A1(new_n287_), .A2(new_n288_), .B1(new_n289_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT79), .B(G8gat), .ZN(new_n294_));
  INV_X1    g093(.A(G1gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT14), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT80), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G15gat), .B(G22gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n297_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G1gat), .B(G8gat), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NOR3_X1   g102(.A1(new_n300_), .A2(new_n301_), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n296_), .A2(new_n298_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT80), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n302_), .B1(new_n306_), .B2(new_n299_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n304_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(G71gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(G78gat), .ZN(new_n310_));
  INV_X1    g109(.A(G78gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(G71gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G57gat), .B(G64gat), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n313_), .B1(new_n314_), .B2(KEYINPUT11), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT68), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n316_), .B1(new_n314_), .B2(KEYINPUT11), .ZN(new_n317_));
  INV_X1    g116(.A(G64gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(G57gat), .ZN(new_n319_));
  INV_X1    g118(.A(G57gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(G64gat), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n319_), .A2(new_n321_), .A3(new_n316_), .A4(KEYINPUT11), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n315_), .B1(new_n317_), .B2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n319_), .A2(new_n321_), .A3(KEYINPUT11), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT68), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n319_), .A2(new_n321_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT11), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n326_), .A2(new_n329_), .A3(new_n313_), .A4(new_n322_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n324_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(G231gat), .ZN(new_n332_));
  INV_X1    g131(.A(G233gat), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n331_), .A2(new_n334_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n324_), .B(new_n330_), .C1(new_n332_), .C2(new_n333_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n308_), .A2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n303_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n306_), .A2(new_n299_), .A3(new_n302_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n341_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G183gat), .B(G211gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT82), .ZN(new_n345_));
  XOR2_X1   g144(.A(G127gat), .B(G155gat), .Z(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  OR2_X1    g146(.A1(new_n344_), .A2(KEYINPUT82), .ZN(new_n348_));
  INV_X1    g147(.A(new_n346_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n344_), .A2(KEYINPUT82), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n348_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n343_), .B1(new_n347_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n347_), .A2(new_n351_), .A3(new_n343_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(KEYINPUT17), .A3(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n338_), .A2(new_n342_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT17), .ZN(new_n358_));
  INV_X1    g157(.A(new_n354_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n358_), .B1(new_n359_), .B2(new_n352_), .ZN(new_n360_));
  AOI22_X1  g159(.A1(new_n338_), .A2(new_n342_), .B1(new_n360_), .B2(new_n355_), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT83), .B1(new_n357_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n338_), .A2(new_n342_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n360_), .A2(new_n355_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT83), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(new_n366_), .A3(new_n356_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n362_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n293_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT13), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n324_), .A2(new_n330_), .ZN(new_n372_));
  AND3_X1   g171(.A1(new_n235_), .A2(new_n236_), .A3(new_n220_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n236_), .B1(new_n235_), .B2(new_n220_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n245_), .A2(new_n253_), .ZN(new_n376_));
  OAI211_X1 g175(.A(KEYINPUT12), .B(new_n372_), .C1(new_n375_), .C2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT69), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n331_), .B1(new_n238_), .B2(new_n254_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT69), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(new_n380_), .A3(KEYINPUT12), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n378_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G230gat), .A2(G233gat), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n238_), .A2(new_n254_), .A3(new_n331_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT12), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n255_), .A2(new_n372_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n382_), .A2(new_n383_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n384_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n383_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(G176gat), .B(G204gat), .Z(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(KEYINPUT71), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT72), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n393_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G120gat), .B(G148gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n388_), .A2(new_n391_), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n398_), .B1(new_n388_), .B2(new_n391_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n371_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n401_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(KEYINPUT13), .A3(new_n399_), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n370_), .A2(new_n405_), .ZN(new_n406_));
  OR2_X1    g205(.A1(new_n406_), .A2(KEYINPUT84), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G113gat), .B(G141gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G169gat), .B(G197gat), .ZN(new_n409_));
  XOR2_X1   g208(.A(new_n408_), .B(new_n409_), .Z(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT85), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G229gat), .A2(G233gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n257_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n257_), .B1(new_n340_), .B2(new_n339_), .ZN(new_n417_));
  OAI211_X1 g216(.A(new_n412_), .B(new_n414_), .C1(new_n416_), .C2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n211_), .A2(new_n216_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n413_), .B(new_n415_), .C1(new_n419_), .C2(new_n308_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n418_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n341_), .A2(new_n215_), .A3(new_n214_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n415_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n412_), .B1(new_n423_), .B2(new_n414_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n411_), .B1(new_n421_), .B2(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n416_), .A2(new_n417_), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT85), .B1(new_n426_), .B2(new_n413_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n427_), .A2(new_n420_), .A3(new_n418_), .A4(new_n410_), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n425_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G227gat), .A2(G233gat), .ZN(new_n430_));
  INV_X1    g229(.A(G15gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(G71gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(new_n227_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT89), .B(G43gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT25), .B(G183gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT26), .B(G190gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G183gat), .A2(G190gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT23), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT23), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n443_), .A2(G183gat), .A3(G190gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(G169gat), .ZN(new_n446_));
  INV_X1    g245(.A(G176gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  OR2_X1    g247(.A1(new_n448_), .A2(KEYINPUT24), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G169gat), .A2(G176gat), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(KEYINPUT24), .A3(new_n450_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n440_), .A2(new_n445_), .A3(new_n449_), .A4(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT87), .ZN(new_n453_));
  OR2_X1    g252(.A1(new_n444_), .A2(new_n453_), .ZN(new_n454_));
  OR2_X1    g253(.A1(G183gat), .A2(G190gat), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n442_), .A2(new_n444_), .A3(new_n453_), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n454_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT86), .B1(new_n446_), .B2(KEYINPUT22), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT22), .B(G169gat), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n447_), .B(new_n458_), .C1(new_n459_), .C2(KEYINPUT86), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n450_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n452_), .B1(new_n457_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT88), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT88), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n464_), .B(new_n452_), .C1(new_n457_), .C2(new_n461_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT30), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n466_), .A2(new_n467_), .ZN(new_n470_));
  AOI21_X1  g269(.A(KEYINPUT90), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n470_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT90), .ZN(new_n473_));
  NOR3_X1   g272(.A1(new_n472_), .A2(new_n473_), .A3(new_n468_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n437_), .B1(new_n471_), .B2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n469_), .A2(KEYINPUT90), .A3(new_n470_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(new_n436_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G113gat), .B(G120gat), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G127gat), .B(G134gat), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT91), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(G134gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(G127gat), .ZN(new_n484_));
  INV_X1    g283(.A(G127gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(G134gat), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n484_), .A2(new_n486_), .A3(new_n481_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n479_), .B1(new_n482_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n484_), .A2(new_n486_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT91), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n480_), .A2(new_n481_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n478_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n488_), .A2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT31), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT92), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n475_), .A2(new_n477_), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n495_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n473_), .B1(new_n472_), .B2(new_n468_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n436_), .B1(new_n498_), .B2(new_n476_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n474_), .A2(new_n437_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n497_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n496_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G226gat), .A2(G233gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT19), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT98), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G211gat), .B(G218gat), .ZN(new_n506_));
  XOR2_X1   g305(.A(new_n506_), .B(KEYINPUT97), .Z(new_n507_));
  XNOR2_X1  g306(.A(G197gat), .B(G204gat), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT21), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n507_), .A2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n506_), .B(KEYINPUT97), .ZN(new_n512_));
  INV_X1    g311(.A(new_n510_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n508_), .A2(new_n509_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n512_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n511_), .A2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT20), .B1(new_n466_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n450_), .B(KEYINPUT101), .Z(new_n519_));
  NAND2_X1  g318(.A1(new_n445_), .A2(new_n455_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n459_), .A2(new_n447_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n519_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n440_), .A2(new_n451_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n454_), .A2(new_n449_), .A3(new_n456_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT99), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT99), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n454_), .A2(new_n449_), .A3(new_n526_), .A4(new_n456_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n523_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n528_), .A2(KEYINPUT100), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT100), .ZN(new_n530_));
  AOI211_X1 g329(.A(new_n530_), .B(new_n523_), .C1(new_n525_), .C2(new_n527_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n522_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n516_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n505_), .B1(new_n518_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT20), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n504_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n537_), .B1(new_n466_), .B2(new_n516_), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n511_), .A2(new_n515_), .A3(new_n522_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n539_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(G8gat), .B(G36gat), .Z(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT18), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G64gat), .B(G92gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NOR3_X1   g346(.A1(new_n534_), .A2(new_n542_), .A3(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n518_), .A2(new_n533_), .A3(new_n505_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n466_), .A2(new_n516_), .ZN(new_n550_));
  XOR2_X1   g349(.A(KEYINPUT105), .B(KEYINPUT20), .Z(new_n551_));
  INV_X1    g350(.A(new_n528_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n551_), .B1(new_n539_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n550_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(new_n504_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n546_), .B1(new_n549_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT27), .ZN(new_n557_));
  NOR3_X1   g356(.A1(new_n548_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n547_), .B1(new_n534_), .B2(new_n542_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n517_), .B1(new_n516_), .B2(new_n532_), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n541_), .B(new_n546_), .C1(new_n560_), .C2(new_n505_), .ZN(new_n561_));
  AOI21_X1  g360(.A(KEYINPUT27), .B1(new_n559_), .B2(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(G141gat), .A2(G148gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT3), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G141gat), .A2(G148gat), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(KEYINPUT93), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT93), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n567_), .A2(G141gat), .A3(G148gat), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT2), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n566_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n565_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT2), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n564_), .A2(new_n570_), .A3(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G155gat), .A2(G162gat), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(G155gat), .A2(G162gat), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n573_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT1), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n579_), .B1(G155gat), .B2(G162gat), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n579_), .A2(G155gat), .A3(G162gat), .ZN(new_n581_));
  AOI22_X1  g380(.A1(new_n574_), .A2(new_n580_), .B1(new_n581_), .B2(KEYINPUT94), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n581_), .A2(KEYINPUT94), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n566_), .A2(new_n568_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n585_), .A2(new_n563_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n578_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT29), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n516_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT95), .B(KEYINPUT28), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(G22gat), .B(G50gat), .Z(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n589_), .A2(new_n590_), .A3(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(KEYINPUT96), .A2(G233gat), .ZN(new_n597_));
  NOR2_X1   g396(.A1(KEYINPUT96), .A2(G233gat), .ZN(new_n598_));
  OAI21_X1  g397(.A(G228gat), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(new_n311_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(new_n228_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n594_), .B1(new_n588_), .B2(KEYINPUT29), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n596_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n602_), .B1(new_n596_), .B2(new_n603_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n593_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n606_), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n591_), .A2(new_n592_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n591_), .A2(new_n592_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n608_), .A2(new_n609_), .A3(new_n610_), .A4(new_n604_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n607_), .A2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G1gat), .B(G29gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(G85gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(KEYINPUT0), .B(G57gat), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n614_), .B(new_n615_), .Z(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  AOI211_X1 g416(.A(new_n585_), .B(new_n563_), .C1(new_n582_), .C2(new_n583_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n577_), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n563_), .A2(KEYINPUT3), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n563_), .A2(KEYINPUT3), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n620_), .A2(new_n621_), .B1(new_n571_), .B2(KEYINPUT2), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n619_), .B1(new_n622_), .B2(new_n570_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n493_), .B1(new_n618_), .B2(new_n623_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n578_), .A2(new_n587_), .A3(new_n492_), .A4(new_n488_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G225gat), .A2(G233gat), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n624_), .A2(KEYINPUT4), .A3(new_n625_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n628_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT4), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n588_), .A2(new_n632_), .A3(new_n493_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n630_), .A2(KEYINPUT102), .A3(new_n631_), .A4(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n629_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n631_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(KEYINPUT102), .B1(new_n637_), .B2(new_n630_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n617_), .B1(new_n635_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT102), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n624_), .A2(KEYINPUT4), .A3(new_n625_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n640_), .B1(new_n641_), .B2(new_n636_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n642_), .A2(new_n616_), .A3(new_n629_), .A4(new_n634_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n612_), .A2(new_n639_), .A3(new_n643_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n558_), .A2(new_n562_), .A3(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n629_), .A2(new_n634_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT33), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n646_), .A2(new_n647_), .A3(new_n616_), .A4(new_n642_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n643_), .A2(KEYINPUT33), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n630_), .A2(new_n628_), .A3(new_n633_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT103), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n631_), .B1(new_n627_), .B2(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n626_), .A2(KEYINPUT103), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n617_), .B(new_n651_), .C1(new_n653_), .C2(new_n654_), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n650_), .A2(new_n561_), .A3(new_n559_), .A4(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n549_), .A2(new_n555_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n546_), .A2(KEYINPUT32), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n541_), .A2(new_n658_), .ZN(new_n661_));
  OAI21_X1  g460(.A(KEYINPUT104), .B1(new_n534_), .B2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n639_), .A2(new_n643_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT104), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n659_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n664_), .B(new_n665_), .C1(new_n560_), .C2(new_n505_), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n660_), .A2(new_n662_), .A3(new_n663_), .A4(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n612_), .B1(new_n656_), .B2(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n502_), .B1(new_n645_), .B2(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n502_), .A2(new_n663_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n612_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n558_), .A2(new_n562_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n670_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n429_), .B1(new_n669_), .B2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n406_), .A2(KEYINPUT84), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n407_), .A2(new_n674_), .A3(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n676_), .A2(new_n295_), .A3(new_n663_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT38), .ZN(new_n678_));
  INV_X1    g477(.A(new_n287_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n679_), .B1(new_n669_), .B2(new_n673_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n405_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n681_), .A2(new_n369_), .A3(new_n429_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n680_), .A2(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n295_), .B1(new_n683_), .B2(new_n663_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT106), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n678_), .A2(new_n685_), .ZN(G1324gat));
  INV_X1    g485(.A(new_n672_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n676_), .A2(new_n687_), .A3(new_n294_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n683_), .A2(new_n687_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G8gat), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n690_), .A2(KEYINPUT39), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(KEYINPUT39), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n688_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT40), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(G1325gat));
  INV_X1    g494(.A(new_n502_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n431_), .B1(new_n683_), .B2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT41), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n676_), .A2(new_n431_), .A3(new_n696_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1326gat));
  INV_X1    g499(.A(G22gat), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n612_), .B(KEYINPUT107), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n683_), .B2(new_n702_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT42), .Z(new_n704_));
  NAND3_X1  g503(.A1(new_n676_), .A2(new_n701_), .A3(new_n702_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1327gat));
  NOR2_X1   g505(.A1(new_n287_), .A2(new_n368_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n707_), .A2(new_n405_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n674_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(G29gat), .B1(new_n710_), .B2(new_n663_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n681_), .A2(new_n368_), .A3(new_n429_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT43), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n669_), .A2(new_n673_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n714_), .B2(new_n293_), .ZN(new_n715_));
  AOI211_X1 g514(.A(KEYINPUT43), .B(new_n292_), .C1(new_n669_), .C2(new_n673_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  OAI211_X1 g518(.A(KEYINPUT44), .B(new_n712_), .C1(new_n715_), .C2(new_n716_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n663_), .A2(G29gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n711_), .B1(new_n721_), .B2(new_n722_), .ZN(G1328gat));
  NOR2_X1   g522(.A1(new_n672_), .A2(G36gat), .ZN(new_n724_));
  XNOR2_X1  g523(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n710_), .A2(new_n724_), .A3(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n725_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n724_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(new_n709_), .B2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n726_), .A2(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n719_), .A2(new_n687_), .A3(new_n720_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n731_), .B2(G36gat), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT46), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n732_), .A2(KEYINPUT109), .A3(new_n733_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n733_), .A2(KEYINPUT109), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n733_), .A2(KEYINPUT109), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n732_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n734_), .A2(new_n737_), .ZN(G1329gat));
  NAND4_X1  g537(.A1(new_n719_), .A2(G43gat), .A3(new_n696_), .A4(new_n720_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n709_), .A2(new_n502_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(G43gat), .B2(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g541(.A(G50gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n710_), .A2(new_n743_), .A3(new_n702_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n721_), .A2(new_n612_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n745_), .A2(KEYINPUT110), .ZN(new_n746_));
  OAI21_X1  g545(.A(G50gat), .B1(new_n745_), .B2(KEYINPUT110), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n744_), .B1(new_n746_), .B2(new_n747_), .ZN(G1331gat));
  NAND2_X1  g547(.A1(new_n425_), .A2(new_n428_), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n405_), .A2(new_n369_), .A3(new_n749_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n680_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n663_), .ZN(new_n753_));
  OAI21_X1  g552(.A(G57gat), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  AOI211_X1 g553(.A(new_n749_), .B(new_n405_), .C1(new_n669_), .C2(new_n673_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n755_), .A2(new_n370_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n756_), .A2(new_n320_), .A3(new_n663_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n754_), .A2(new_n757_), .ZN(G1332gat));
  NAND3_X1  g557(.A1(new_n756_), .A2(new_n318_), .A3(new_n687_), .ZN(new_n759_));
  OAI21_X1  g558(.A(G64gat), .B1(new_n752_), .B2(new_n672_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n760_), .A2(KEYINPUT48), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n760_), .A2(KEYINPUT48), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n759_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT111), .ZN(G1333gat));
  AOI21_X1  g563(.A(new_n309_), .B1(new_n751_), .B2(new_n696_), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT49), .Z(new_n766_));
  NAND3_X1  g565(.A1(new_n756_), .A2(new_n309_), .A3(new_n696_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(G1334gat));
  NAND3_X1  g567(.A1(new_n756_), .A2(new_n311_), .A3(new_n702_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n751_), .A2(new_n702_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n770_), .A2(G78gat), .A3(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n770_), .B2(G78gat), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT113), .ZN(G1335gat));
  NOR3_X1   g574(.A1(new_n405_), .A2(new_n368_), .A3(new_n749_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n776_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n777_));
  OAI21_X1  g576(.A(G85gat), .B1(new_n777_), .B2(new_n753_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n755_), .A2(new_n707_), .ZN(new_n779_));
  INV_X1    g578(.A(G85gat), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n780_), .A3(new_n663_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n778_), .A2(new_n781_), .ZN(G1336gat));
  OAI21_X1  g581(.A(G92gat), .B1(new_n777_), .B2(new_n672_), .ZN(new_n783_));
  INV_X1    g582(.A(G92gat), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n779_), .A2(new_n784_), .A3(new_n687_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(G1337gat));
  NAND4_X1  g585(.A1(new_n779_), .A2(new_n696_), .A3(new_n239_), .A4(new_n240_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT114), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n787_), .A2(new_n788_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n777_), .A2(new_n502_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n792_), .A2(new_n227_), .ZN(new_n793_));
  OAI21_X1  g592(.A(KEYINPUT51), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT51), .ZN(new_n795_));
  OAI221_X1 g594(.A(new_n795_), .B1(new_n792_), .B2(new_n227_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(G1338gat));
  NAND3_X1  g596(.A1(new_n779_), .A2(new_n228_), .A3(new_n612_), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n612_), .B(new_n776_), .C1(new_n715_), .C2(new_n716_), .ZN(new_n799_));
  XOR2_X1   g598(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n800_));
  AND3_X1   g599(.A1(new_n799_), .A2(G106gat), .A3(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n799_), .B2(G106gat), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n798_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  XOR2_X1   g602(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n804_));
  XNOR2_X1  g603(.A(new_n803_), .B(new_n804_), .ZN(G1339gat));
  NOR2_X1   g604(.A1(new_n687_), .A2(new_n612_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(new_n663_), .A3(new_n696_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  XOR2_X1   g607(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n809_));
  AOI21_X1  g608(.A(new_n400_), .B1(new_n425_), .B2(new_n428_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n383_), .B1(new_n382_), .B2(new_n387_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n388_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n382_), .A2(KEYINPUT55), .A3(new_n383_), .A4(new_n387_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n398_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT56), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT56), .ZN(new_n818_));
  AOI211_X1 g617(.A(new_n818_), .B(new_n398_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n810_), .B1(new_n817_), .B2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n415_), .B1(new_n419_), .B2(new_n308_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n413_), .B1(new_n821_), .B2(KEYINPUT118), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n822_), .B1(KEYINPUT118), .B2(new_n821_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n410_), .B1(new_n423_), .B2(new_n413_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n428_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n400_), .A2(new_n401_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n820_), .A2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT57), .B1(new_n830_), .B2(new_n287_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832_));
  AOI211_X1 g631(.A(new_n832_), .B(new_n679_), .C1(new_n820_), .C2(new_n829_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n826_), .A2(new_n400_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n835_), .B1(new_n817_), .B2(new_n819_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(KEYINPUT119), .A2(KEYINPUT58), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  OAI221_X1 g637(.A(new_n835_), .B1(KEYINPUT119), .B2(KEYINPUT58), .C1(new_n817_), .C2(new_n819_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n838_), .A2(new_n839_), .A3(new_n293_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n368_), .B1(new_n834_), .B2(new_n840_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n368_), .A2(KEYINPUT117), .A3(new_n425_), .A4(new_n428_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n842_), .A2(new_n402_), .A3(new_n404_), .ZN(new_n843_));
  AOI21_X1  g642(.A(KEYINPUT117), .B1(new_n429_), .B2(new_n368_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n845_), .A2(new_n846_), .A3(new_n292_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n845_), .B2(new_n292_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n808_), .B(new_n809_), .C1(new_n841_), .C2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n749_), .A2(new_n399_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n380_), .B1(new_n379_), .B2(KEYINPUT12), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT12), .ZN(new_n853_));
  NOR4_X1   g652(.A1(new_n258_), .A2(KEYINPUT69), .A3(new_n331_), .A4(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n387_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n812_), .B1(new_n855_), .B2(new_n390_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n855_), .A2(new_n390_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n814_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n816_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n818_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n815_), .A2(KEYINPUT56), .A3(new_n816_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n851_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n287_), .B1(new_n863_), .B2(new_n828_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n832_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n830_), .A2(KEYINPUT57), .A3(new_n287_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n840_), .A3(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n849_), .B1(new_n867_), .B2(new_n369_), .ZN(new_n868_));
  OAI21_X1  g667(.A(KEYINPUT59), .B1(new_n868_), .B2(new_n807_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n850_), .A2(new_n869_), .A3(new_n749_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(G113gat), .ZN(new_n871_));
  INV_X1    g670(.A(new_n868_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n429_), .A2(G113gat), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n872_), .A2(new_n808_), .A3(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n871_), .A2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT121), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n871_), .A2(new_n877_), .A3(new_n874_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(G1340gat));
  NAND3_X1  g678(.A1(new_n850_), .A2(new_n869_), .A3(new_n681_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(G120gat), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT60), .ZN(new_n882_));
  AOI21_X1  g681(.A(G120gat), .B1(new_n681_), .B2(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n883_), .B1(new_n882_), .B2(G120gat), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n872_), .A2(new_n808_), .A3(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n881_), .A2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(KEYINPUT122), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT122), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n881_), .A2(new_n888_), .A3(new_n885_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n889_), .ZN(G1341gat));
  AND3_X1   g689(.A1(new_n850_), .A2(new_n869_), .A3(new_n368_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n872_), .A2(new_n808_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n368_), .A2(new_n485_), .ZN(new_n893_));
  OAI22_X1  g692(.A1(new_n891_), .A2(new_n485_), .B1(new_n892_), .B2(new_n893_), .ZN(G1342gat));
  AND3_X1   g693(.A1(new_n850_), .A2(new_n869_), .A3(new_n293_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n679_), .A2(new_n483_), .ZN(new_n896_));
  OAI22_X1  g695(.A1(new_n895_), .A2(new_n483_), .B1(new_n892_), .B2(new_n896_), .ZN(G1343gat));
  NOR4_X1   g696(.A1(new_n687_), .A2(new_n696_), .A3(new_n753_), .A4(new_n671_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n868_), .A2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n749_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n681_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g703(.A1(new_n900_), .A2(new_n368_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(KEYINPUT123), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n900_), .A2(new_n907_), .A3(new_n368_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n908_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(KEYINPUT61), .B(G155gat), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n909_), .B(new_n910_), .ZN(G1346gat));
  INV_X1    g710(.A(new_n900_), .ZN(new_n912_));
  OR3_X1    g711(.A1(new_n912_), .A2(G162gat), .A3(new_n287_), .ZN(new_n913_));
  OAI21_X1  g712(.A(G162gat), .B1(new_n912_), .B2(new_n292_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1347gat));
  NAND2_X1  g714(.A1(new_n687_), .A2(new_n670_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(new_n702_), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n749_), .B(new_n917_), .C1(new_n841_), .C2(new_n849_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(G169gat), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n868_), .A2(new_n702_), .A3(new_n916_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n922_), .A2(new_n459_), .A3(new_n749_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n918_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n921_), .A2(new_n923_), .A3(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(KEYINPUT124), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n927_));
  NAND4_X1  g726(.A1(new_n921_), .A2(new_n923_), .A3(new_n927_), .A4(new_n924_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n926_), .A2(new_n928_), .ZN(G1348gat));
  AOI21_X1  g728(.A(G176gat), .B1(new_n922_), .B2(new_n681_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n868_), .A2(new_n612_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n916_), .A2(new_n447_), .A3(new_n405_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n930_), .B1(new_n931_), .B2(new_n932_), .ZN(G1349gat));
  NAND4_X1  g732(.A1(new_n931_), .A2(new_n687_), .A3(new_n670_), .A4(new_n368_), .ZN(new_n934_));
  INV_X1    g733(.A(G183gat), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n369_), .A2(new_n438_), .ZN(new_n936_));
  AOI22_X1  g735(.A1(new_n934_), .A2(new_n935_), .B1(new_n922_), .B2(new_n936_), .ZN(G1350gat));
  INV_X1    g736(.A(new_n922_), .ZN(new_n938_));
  OAI21_X1  g737(.A(G190gat), .B1(new_n938_), .B2(new_n292_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n922_), .A2(new_n439_), .A3(new_n679_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(G1351gat));
  NAND3_X1  g740(.A1(new_n502_), .A2(new_n753_), .A3(new_n612_), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n943_));
  OR2_X1    g742(.A1(new_n942_), .A2(new_n943_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n942_), .A2(new_n943_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n944_), .A2(new_n687_), .A3(new_n945_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n868_), .A2(new_n946_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(new_n749_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g748(.A1(new_n947_), .A2(new_n681_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g750(.A(new_n369_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n947_), .A2(new_n952_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n953_), .A2(KEYINPUT126), .ZN(new_n954_));
  INV_X1    g753(.A(new_n954_), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n953_), .A2(KEYINPUT126), .ZN(new_n956_));
  OAI22_X1  g755(.A1(new_n955_), .A2(new_n956_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n957_));
  INV_X1    g756(.A(new_n956_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n958_), .A2(new_n959_), .A3(new_n954_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n957_), .A2(new_n960_), .ZN(G1354gat));
  INV_X1    g760(.A(new_n947_), .ZN(new_n962_));
  OR3_X1    g761(.A1(new_n962_), .A2(G218gat), .A3(new_n287_), .ZN(new_n963_));
  OAI21_X1  g762(.A(G218gat), .B1(new_n962_), .B2(new_n292_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n963_), .A2(new_n964_), .ZN(G1355gat));
endmodule


