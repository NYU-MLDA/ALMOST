//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n625_, new_n626_, new_n627_, new_n628_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n826_, new_n827_, new_n828_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n861_, new_n863_, new_n864_,
    new_n865_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT19), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT20), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT25), .B(G183gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT26), .B(G190gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT90), .ZN(new_n209_));
  AND2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n208_), .A2(new_n209_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n207_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT23), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(G183gat), .A3(G190gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n216_), .A3(KEYINPUT82), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT82), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n213_), .A2(new_n218_), .A3(KEYINPUT23), .ZN(new_n219_));
  OR3_X1    g018(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n217_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT91), .ZN(new_n222_));
  INV_X1    g021(.A(G169gat), .ZN(new_n223_));
  INV_X1    g022(.A(G176gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(KEYINPUT24), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT91), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n217_), .A2(new_n228_), .A3(new_n219_), .A4(new_n220_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n212_), .A2(new_n222_), .A3(new_n227_), .A4(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n214_), .A2(new_n216_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n231_), .B1(G183gat), .B2(G190gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT22), .B(G169gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT92), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n226_), .B(new_n232_), .C1(new_n234_), .C2(G176gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n230_), .A2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G197gat), .B(G204gat), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G211gat), .B(G218gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT88), .ZN(new_n240_));
  AOI22_X1  g039(.A1(new_n238_), .A2(KEYINPUT21), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT21), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n237_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(new_n239_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n237_), .A2(new_n242_), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n239_), .B(new_n243_), .C1(new_n246_), .C2(new_n240_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n206_), .B1(new_n236_), .B2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT78), .B(G183gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT25), .ZN(new_n252_));
  OR2_X1    g051(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT26), .ZN(new_n255_));
  OAI21_X1  g054(.A(KEYINPUT79), .B1(new_n255_), .B2(G190gat), .ZN(new_n256_));
  OR2_X1    g055(.A1(new_n208_), .A2(KEYINPUT79), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n254_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n258_), .A2(new_n231_), .A3(new_n227_), .A4(new_n220_), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n217_), .B(new_n219_), .C1(G190gat), .C2(new_n251_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT22), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT80), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT80), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT22), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n223_), .B1(new_n262_), .B2(new_n264_), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n265_), .A2(KEYINPUT81), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT81), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n267_), .B1(KEYINPUT22), .B2(new_n223_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n224_), .B1(new_n265_), .B2(new_n268_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n260_), .B(new_n226_), .C1(new_n266_), .C2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n259_), .A2(new_n248_), .A3(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n205_), .B1(new_n250_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G8gat), .B(G36gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT18), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(G64gat), .ZN(new_n276_));
  INV_X1    g075(.A(G92gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n259_), .A2(new_n270_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n249_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n230_), .A2(new_n248_), .A3(new_n235_), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n280_), .A2(KEYINPUT20), .A3(new_n205_), .A4(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n273_), .A2(new_n278_), .A3(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n278_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n282_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n284_), .B1(new_n285_), .B2(new_n272_), .ZN(new_n286_));
  AOI21_X1  g085(.A(KEYINPUT27), .B1(new_n283_), .B2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n248_), .B1(new_n259_), .B2(new_n270_), .ZN(new_n288_));
  AND2_X1   g087(.A1(KEYINPUT97), .A2(KEYINPUT20), .ZN(new_n289_));
  NOR2_X1   g088(.A1(KEYINPUT97), .A2(KEYINPUT20), .ZN(new_n290_));
  NOR3_X1   g089(.A1(new_n288_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n205_), .B1(new_n291_), .B2(new_n281_), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n250_), .A2(new_n205_), .A3(new_n271_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n284_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT101), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(new_n295_), .A3(new_n283_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n273_), .A2(KEYINPUT101), .A3(new_n278_), .A4(new_n282_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n287_), .B1(new_n298_), .B2(KEYINPUT27), .ZN(new_n299_));
  XOR2_X1   g098(.A(G78gat), .B(G106gat), .Z(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  OR2_X1    g100(.A1(G155gat), .A2(G162gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT86), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(KEYINPUT86), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n308_));
  AND2_X1   g107(.A1(G141gat), .A2(G148gat), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n307_), .B(new_n308_), .C1(new_n309_), .C2(KEYINPUT2), .ZN(new_n310_));
  NOR2_X1   g109(.A1(G141gat), .A2(G148gat), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT3), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n304_), .B1(new_n310_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n303_), .A2(KEYINPUT1), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT85), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n315_), .A2(new_n316_), .A3(new_n302_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n316_), .B1(new_n315_), .B2(new_n302_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n303_), .A2(KEYINPUT1), .ZN(new_n319_));
  NOR3_X1   g118(.A1(new_n317_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n309_), .A2(new_n311_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n314_), .B1(new_n320_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT29), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n249_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT87), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(G233gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n327_), .A2(G233gat), .ZN(new_n330_));
  OAI21_X1  g129(.A(G228gat), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n326_), .B(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT89), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT28), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n324_), .A2(new_n335_), .A3(new_n325_), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT28), .B1(new_n323_), .B2(KEYINPUT29), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G22gat), .B(G50gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n339_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n336_), .A2(new_n337_), .A3(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n334_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n331_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n326_), .B(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT89), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n334_), .A2(new_n347_), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n301_), .B(new_n344_), .C1(new_n348_), .C2(new_n343_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n343_), .B1(new_n334_), .B2(new_n347_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n334_), .A2(new_n343_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n300_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n349_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT100), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G127gat), .A2(G134gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(G127gat), .A2(G134gat), .ZN(new_n357_));
  OAI21_X1  g156(.A(G113gat), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(G127gat), .ZN(new_n359_));
  INV_X1    g158(.A(G134gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(G113gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n361_), .A2(new_n362_), .A3(new_n355_), .ZN(new_n363_));
  AND3_X1   g162(.A1(new_n358_), .A2(new_n363_), .A3(G120gat), .ZN(new_n364_));
  AOI21_X1  g163(.A(G120gat), .B1(new_n358_), .B2(new_n363_), .ZN(new_n365_));
  OR2_X1    g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n323_), .A2(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n364_), .A2(new_n365_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n315_), .A2(new_n302_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT85), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n315_), .A2(new_n302_), .A3(new_n316_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n319_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n321_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n368_), .A2(new_n374_), .A3(new_n314_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n367_), .A2(KEYINPUT4), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT4), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n323_), .A2(new_n366_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379_));
  XOR2_X1   g178(.A(new_n379_), .B(KEYINPUT93), .Z(new_n380_));
  NAND3_X1  g179(.A1(new_n376_), .A2(new_n378_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT94), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n367_), .A2(new_n375_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n379_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n376_), .A2(KEYINPUT94), .A3(new_n378_), .A4(new_n380_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n383_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT98), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(G85gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT0), .ZN(new_n391_));
  INV_X1    g190(.A(G57gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n387_), .A2(new_n388_), .A3(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n388_), .B1(new_n387_), .B2(new_n394_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n383_), .A2(new_n385_), .A3(new_n393_), .A4(new_n386_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n354_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n387_), .A2(new_n394_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT98), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n387_), .A2(new_n388_), .A3(new_n394_), .ZN(new_n402_));
  AND4_X1   g201(.A1(new_n354_), .A2(new_n401_), .A3(new_n398_), .A4(new_n402_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n299_), .B(new_n353_), .C1(new_n399_), .C2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT102), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n397_), .A2(new_n354_), .A3(new_n398_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n401_), .A2(new_n398_), .A3(new_n402_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT100), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n410_), .A2(KEYINPUT102), .A3(new_n299_), .A4(new_n353_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n376_), .A2(new_n379_), .A3(new_n378_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n384_), .A2(KEYINPUT96), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n380_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n384_), .A2(KEYINPUT96), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n394_), .B(new_n412_), .C1(new_n414_), .C2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT95), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n417_), .A2(KEYINPUT33), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n283_), .B(new_n286_), .C1(new_n398_), .C2(new_n418_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n398_), .A2(new_n418_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n278_), .A2(KEYINPUT32), .ZN(new_n422_));
  NOR3_X1   g221(.A1(new_n422_), .A2(new_n285_), .A3(new_n272_), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n292_), .A2(new_n293_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n423_), .B1(new_n424_), .B2(new_n422_), .ZN(new_n425_));
  AOI22_X1  g224(.A1(new_n416_), .A2(new_n421_), .B1(new_n408_), .B2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT99), .B1(new_n426_), .B2(new_n353_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n353_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT99), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n408_), .A2(new_n425_), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n421_), .A2(new_n416_), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n428_), .B(new_n429_), .C1(new_n430_), .C2(new_n431_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n406_), .A2(new_n411_), .A3(new_n427_), .A4(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n279_), .B(KEYINPUT30), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(G99gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G227gat), .A2(G233gat), .ZN(new_n436_));
  INV_X1    g235(.A(G15gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(G71gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT83), .B(G43gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n435_), .B(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT84), .ZN(new_n443_));
  OR2_X1    g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n366_), .B(KEYINPUT31), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n442_), .A2(new_n443_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n444_), .A2(new_n447_), .A3(new_n445_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n433_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT103), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n449_), .A2(new_n353_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n452_), .A2(new_n410_), .A3(new_n299_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT103), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n433_), .A2(new_n454_), .A3(new_n449_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n451_), .A2(new_n453_), .A3(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G29gat), .B(G36gat), .ZN(new_n457_));
  INV_X1    g256(.A(G43gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(G50gat), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT15), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(G8gat), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT74), .ZN(new_n465_));
  OR2_X1    g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G15gat), .B(G22gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n464_), .A2(new_n465_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G1gat), .B(G8gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n462_), .A2(new_n471_), .ZN(new_n472_));
  OR2_X1    g271(.A1(new_n471_), .A2(new_n460_), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G229gat), .A2(G233gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n475_), .B(KEYINPUT76), .Z(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT77), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n471_), .B(new_n460_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(G229gat), .A3(G233gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G113gat), .B(G141gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(new_n223_), .ZN(new_n483_));
  INV_X1    g282(.A(G197gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n481_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n485_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n478_), .A2(new_n480_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n456_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT13), .ZN(new_n491_));
  XOR2_X1   g290(.A(G85gat), .B(G92gat), .Z(new_n492_));
  INV_X1    g291(.A(G99gat), .ZN(new_n493_));
  INV_X1    g292(.A(G106gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT7), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G99gat), .A2(G106gat), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT6), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n492_), .B1(new_n496_), .B2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT8), .ZN(new_n501_));
  INV_X1    g300(.A(G85gat), .ZN(new_n502_));
  NOR3_X1   g301(.A1(new_n502_), .A2(new_n277_), .A3(KEYINPUT9), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n499_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n492_), .A2(KEYINPUT9), .ZN(new_n505_));
  XOR2_X1   g304(.A(KEYINPUT10), .B(G99gat), .Z(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n494_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n504_), .A2(new_n505_), .A3(new_n507_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n508_), .A2(KEYINPUT64), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(KEYINPUT64), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n501_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G57gat), .B(G64gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT11), .ZN(new_n513_));
  XOR2_X1   g312(.A(G71gat), .B(G78gat), .Z(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n515_), .B1(KEYINPUT11), .B2(new_n512_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n511_), .A2(new_n516_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n509_), .A2(new_n510_), .A3(KEYINPUT65), .ZN(new_n518_));
  AOI21_X1  g317(.A(KEYINPUT65), .B1(new_n509_), .B2(new_n510_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n501_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n520_), .A2(KEYINPUT12), .A3(new_n516_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT66), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n517_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n511_), .A2(new_n516_), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n524_), .A2(KEYINPUT12), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G230gat), .A2(G233gat), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n520_), .A2(KEYINPUT66), .A3(KEYINPUT12), .A4(new_n516_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n523_), .A2(new_n525_), .A3(new_n526_), .A4(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n526_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n529_), .B1(new_n524_), .B2(new_n517_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G120gat), .B(G148gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT5), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G176gat), .B(G204gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n535_), .B(new_n536_), .Z(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n531_), .A2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n528_), .A2(new_n530_), .A3(new_n537_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n539_), .A2(KEYINPUT69), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(KEYINPUT69), .B1(new_n539_), .B2(new_n540_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n491_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n543_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n545_), .A2(KEYINPUT13), .A3(new_n541_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n520_), .A2(new_n462_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G232gat), .A2(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT34), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n550_), .A2(KEYINPUT35), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n551_), .A2(KEYINPUT72), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(KEYINPUT72), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n552_), .B(new_n553_), .C1(new_n511_), .C2(new_n460_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n548_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT71), .ZN(new_n556_));
  OAI211_X1 g355(.A(KEYINPUT35), .B(new_n550_), .C1(new_n554_), .C2(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n555_), .B(new_n557_), .Z(new_n558_));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT73), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(G134gat), .ZN(new_n561_));
  INV_X1    g360(.A(G162gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT36), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n558_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT36), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n558_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n565_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n471_), .B(new_n516_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n571_), .B(KEYINPUT75), .Z(new_n572_));
  XNOR2_X1  g371(.A(new_n570_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G127gat), .B(G155gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT16), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(G183gat), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n576_), .B(G211gat), .Z(new_n577_));
  INV_X1    g376(.A(KEYINPUT17), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n577_), .A2(new_n578_), .ZN(new_n580_));
  NOR3_X1   g379(.A1(new_n573_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n581_), .B1(new_n579_), .B2(new_n573_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n569_), .A2(new_n583_), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n490_), .A2(new_n547_), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n410_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n202_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT104), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT70), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n547_), .B(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n569_), .B(KEYINPUT37), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n591_), .A2(new_n583_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n590_), .A2(new_n456_), .A3(new_n489_), .A4(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n593_), .A2(new_n410_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n588_), .B1(new_n594_), .B2(new_n202_), .ZN(new_n595_));
  NOR4_X1   g394(.A1(new_n593_), .A2(KEYINPUT104), .A3(G1gat), .A4(new_n410_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n587_), .B1(new_n597_), .B2(KEYINPUT38), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n490_), .A2(new_n586_), .A3(new_n590_), .A4(new_n592_), .ZN(new_n599_));
  OAI21_X1  g398(.A(KEYINPUT104), .B1(new_n599_), .B2(G1gat), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n594_), .A2(new_n588_), .A3(new_n202_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT38), .ZN(new_n603_));
  AOI21_X1  g402(.A(KEYINPUT105), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT105), .ZN(new_n605_));
  AOI211_X1 g404(.A(new_n605_), .B(KEYINPUT38), .C1(new_n600_), .C2(new_n601_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n598_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT106), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n598_), .B(KEYINPUT106), .C1(new_n604_), .C2(new_n606_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(G1324gat));
  INV_X1    g410(.A(new_n299_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n585_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(G8gat), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT107), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT39), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n614_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  OR3_X1    g416(.A1(new_n593_), .A2(G8gat), .A3(new_n299_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(KEYINPUT107), .A2(KEYINPUT39), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n615_), .A2(new_n616_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n613_), .A2(G8gat), .A3(new_n619_), .A4(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n617_), .A2(new_n618_), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT40), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(G1325gat));
  INV_X1    g423(.A(new_n449_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n437_), .B1(new_n585_), .B2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT41), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n593_), .A2(G15gat), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n627_), .B1(new_n449_), .B2(new_n628_), .ZN(G1326gat));
  INV_X1    g428(.A(G22gat), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n630_), .B1(new_n585_), .B2(new_n353_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT42), .Z(new_n632_));
  NAND2_X1  g431(.A1(new_n353_), .A2(new_n630_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n632_), .B1(new_n593_), .B2(new_n633_), .ZN(G1327gat));
  INV_X1    g433(.A(new_n489_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n456_), .A2(new_n591_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT43), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT43), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n456_), .A2(new_n638_), .A3(new_n591_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n635_), .B1(new_n637_), .B2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n641_));
  OR2_X1    g440(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n642_));
  INV_X1    g441(.A(new_n547_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n643_), .A2(new_n582_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n640_), .A2(new_n641_), .A3(new_n642_), .A4(new_n644_), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n456_), .A2(new_n638_), .A3(new_n591_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n638_), .B1(new_n456_), .B2(new_n591_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n489_), .B(new_n644_), .C1(new_n646_), .C2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n648_), .A2(KEYINPUT108), .A3(KEYINPUT44), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n645_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(G29gat), .B1(new_n651_), .B2(new_n410_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n569_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n653_), .A2(new_n582_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n490_), .A2(new_n547_), .A3(new_n654_), .ZN(new_n655_));
  OR3_X1    g454(.A1(new_n655_), .A2(G29gat), .A3(new_n410_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n652_), .A2(new_n656_), .ZN(G1328gat));
  INV_X1    g456(.A(G36gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n658_), .B1(new_n650_), .B2(new_n612_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n655_), .A2(G36gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n662_), .B1(new_n663_), .B2(new_n612_), .ZN(new_n664_));
  NOR4_X1   g463(.A1(new_n655_), .A2(G36gat), .A3(new_n299_), .A4(new_n661_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n660_), .A2(KEYINPUT46), .A3(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT46), .ZN(new_n668_));
  INV_X1    g467(.A(new_n666_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(new_n669_), .B2(new_n659_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n667_), .A2(new_n670_), .ZN(G1329gat));
  AOI21_X1  g470(.A(new_n458_), .B1(new_n650_), .B2(new_n625_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT47), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n655_), .A2(G43gat), .A3(new_n449_), .ZN(new_n674_));
  OR3_X1    g473(.A1(new_n672_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n673_), .B1(new_n672_), .B2(new_n674_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1330gat));
  OAI21_X1  g476(.A(G50gat), .B1(new_n651_), .B2(new_n428_), .ZN(new_n678_));
  OR3_X1    g477(.A1(new_n655_), .A2(G50gat), .A3(new_n428_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1331gat));
  INV_X1    g479(.A(new_n590_), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n681_), .A2(new_n635_), .A3(new_n456_), .A4(new_n584_), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n682_), .A2(new_n392_), .A3(new_n410_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n456_), .A2(new_n635_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT110), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n685_), .A2(new_n643_), .A3(new_n592_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(new_n586_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n683_), .B1(new_n687_), .B2(new_n392_), .ZN(G1332gat));
  INV_X1    g487(.A(G64gat), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n686_), .A2(new_n689_), .A3(new_n612_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G64gat), .B1(new_n682_), .B2(new_n299_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT48), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(G1333gat));
  INV_X1    g492(.A(G71gat), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n686_), .A2(new_n694_), .A3(new_n625_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G71gat), .B1(new_n682_), .B2(new_n449_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT49), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(G1334gat));
  INV_X1    g497(.A(G78gat), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n686_), .A2(new_n699_), .A3(new_n353_), .ZN(new_n700_));
  OAI21_X1  g499(.A(G78gat), .B1(new_n682_), .B2(new_n428_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT50), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(G1335gat));
  NAND2_X1  g502(.A1(new_n637_), .A2(new_n639_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n547_), .A2(new_n489_), .A3(new_n582_), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n704_), .A2(G85gat), .A3(new_n586_), .A4(new_n705_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n685_), .A2(new_n586_), .A3(new_n681_), .A4(new_n654_), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n707_), .A2(KEYINPUT111), .A3(new_n502_), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT111), .B1(new_n707_), .B2(new_n502_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n706_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT112), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  OAI211_X1 g511(.A(KEYINPUT112), .B(new_n706_), .C1(new_n708_), .C2(new_n709_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1336gat));
  NAND2_X1  g513(.A1(new_n704_), .A2(new_n705_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n715_), .A2(new_n277_), .A3(new_n299_), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n685_), .A2(new_n681_), .A3(new_n654_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(new_n612_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n716_), .B1(new_n718_), .B2(new_n277_), .ZN(G1337gat));
  NAND3_X1  g518(.A1(new_n717_), .A2(new_n506_), .A3(new_n625_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n721_));
  OAI21_X1  g520(.A(G99gat), .B1(new_n715_), .B2(new_n449_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n720_), .A2(new_n721_), .A3(new_n722_), .ZN(new_n723_));
  OR2_X1    g522(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n723_), .B(new_n724_), .ZN(G1338gat));
  NAND3_X1  g524(.A1(new_n717_), .A2(new_n494_), .A3(new_n353_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n353_), .B(new_n705_), .C1(new_n646_), .C2(new_n647_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT114), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n727_), .A2(new_n728_), .A3(G106gat), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n728_), .B1(new_n727_), .B2(G106gat), .ZN(new_n731_));
  NOR3_X1   g530(.A1(new_n730_), .A2(new_n731_), .A3(KEYINPUT52), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT52), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n727_), .A2(G106gat), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT114), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n733_), .B1(new_n735_), .B2(new_n729_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n726_), .B1(new_n732_), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT53), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT53), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n739_), .B(new_n726_), .C1(new_n732_), .C2(new_n736_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(G1339gat));
  NAND2_X1  g540(.A1(new_n489_), .A2(new_n540_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT55), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n528_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT116), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n528_), .A2(new_n743_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n528_), .A2(KEYINPUT116), .A3(new_n743_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n523_), .A2(new_n525_), .A3(new_n527_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(new_n529_), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n746_), .A2(new_n747_), .A3(new_n748_), .A4(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(KEYINPUT56), .B1(new_n751_), .B2(new_n538_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT117), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n742_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n751_), .A2(new_n538_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT56), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n751_), .A2(KEYINPUT56), .A3(new_n538_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n757_), .A2(KEYINPUT117), .A3(new_n758_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n754_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n545_), .A2(new_n541_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n487_), .B1(new_n479_), .B2(new_n476_), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT118), .Z(new_n763_));
  INV_X1    g562(.A(new_n474_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(new_n476_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n488_), .A2(new_n765_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n761_), .A2(new_n766_), .ZN(new_n767_));
  OAI211_X1 g566(.A(KEYINPUT57), .B(new_n653_), .C1(new_n760_), .C2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT57), .ZN(new_n769_));
  AOI22_X1  g568(.A1(new_n754_), .A2(new_n759_), .B1(new_n761_), .B2(new_n766_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(new_n770_), .B2(new_n569_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n757_), .A2(new_n758_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n772_), .A2(new_n540_), .A3(new_n766_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT58), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n772_), .A2(KEYINPUT58), .A3(new_n540_), .A4(new_n766_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n591_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n768_), .A2(new_n771_), .A3(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n591_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n544_), .A2(new_n546_), .A3(new_n635_), .A4(new_n582_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n780_), .A2(KEYINPUT115), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n780_), .A2(KEYINPUT115), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n779_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT54), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n785_), .B(new_n779_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n778_), .A2(new_n583_), .B1(new_n784_), .B2(new_n786_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n410_), .A2(new_n612_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n452_), .A2(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(G113gat), .B1(new_n790_), .B2(new_n489_), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n791_), .A2(KEYINPUT119), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(KEYINPUT119), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n771_), .A2(new_n777_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT120), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT120), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n771_), .A2(new_n777_), .A3(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n795_), .A2(new_n768_), .A3(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n583_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n784_), .A2(new_n786_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n789_), .A2(KEYINPUT59), .ZN(new_n802_));
  INV_X1    g601(.A(new_n787_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n789_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  AOI22_X1  g604(.A1(new_n801_), .A2(new_n802_), .B1(new_n805_), .B2(KEYINPUT59), .ZN(new_n806_));
  XNOR2_X1  g605(.A(KEYINPUT121), .B(G113gat), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n489_), .A2(new_n807_), .ZN(new_n808_));
  XOR2_X1   g607(.A(new_n808_), .B(KEYINPUT122), .Z(new_n809_));
  AOI22_X1  g608(.A1(new_n792_), .A2(new_n793_), .B1(new_n806_), .B2(new_n809_), .ZN(G1340gat));
  NAND2_X1  g609(.A1(new_n801_), .A2(new_n802_), .ZN(new_n811_));
  OAI21_X1  g610(.A(KEYINPUT59), .B1(new_n787_), .B2(new_n789_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n811_), .A2(KEYINPUT124), .A3(new_n681_), .A4(new_n812_), .ZN(new_n813_));
  AOI22_X1  g612(.A1(new_n798_), .A2(new_n583_), .B1(new_n784_), .B2(new_n786_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n802_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n681_), .B(new_n812_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT124), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n813_), .A2(new_n818_), .A3(G120gat), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT60), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n820_), .B1(new_n547_), .B2(G120gat), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n790_), .B(new_n821_), .C1(new_n820_), .C2(G120gat), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT123), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n822_), .B(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n819_), .A2(new_n824_), .ZN(G1341gat));
  NAND2_X1  g624(.A1(new_n806_), .A2(new_n582_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(G127gat), .ZN(new_n827_));
  OR4_X1    g626(.A1(G127gat), .A2(new_n800_), .A3(new_n583_), .A4(new_n789_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(G1342gat));
  NAND3_X1  g628(.A1(new_n806_), .A2(G134gat), .A3(new_n591_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n360_), .B1(new_n805_), .B2(new_n653_), .ZN(new_n831_));
  OR2_X1    g630(.A1(new_n831_), .A2(KEYINPUT125), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(KEYINPUT125), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n830_), .A2(new_n832_), .A3(new_n833_), .ZN(G1343gat));
  NOR3_X1   g633(.A1(new_n787_), .A2(new_n625_), .A3(new_n428_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n835_), .A2(new_n788_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n489_), .ZN(new_n837_));
  XOR2_X1   g636(.A(KEYINPUT126), .B(G141gat), .Z(new_n838_));
  XNOR2_X1  g637(.A(new_n837_), .B(new_n838_), .ZN(G1344gat));
  NAND2_X1  g638(.A1(new_n836_), .A2(new_n681_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g640(.A1(new_n836_), .A2(new_n582_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(KEYINPUT61), .B(G155gat), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(G1346gat));
  AOI21_X1  g643(.A(G162gat), .B1(new_n836_), .B2(new_n569_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n779_), .A2(new_n562_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n845_), .B1(new_n836_), .B2(new_n846_), .ZN(G1347gat));
  NOR2_X1   g646(.A1(new_n586_), .A2(new_n299_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n452_), .A2(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n814_), .A2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n223_), .B1(new_n850_), .B2(new_n489_), .ZN(new_n851_));
  NOR4_X1   g650(.A1(new_n814_), .A2(new_n635_), .A3(new_n234_), .A4(new_n849_), .ZN(new_n852_));
  OAI21_X1  g651(.A(KEYINPUT62), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT62), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n814_), .A2(new_n635_), .A3(new_n849_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n223_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n853_), .A2(new_n856_), .ZN(G1348gat));
  NAND3_X1  g656(.A1(new_n850_), .A2(new_n224_), .A3(new_n643_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n787_), .A2(new_n590_), .A3(new_n849_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n224_), .B2(new_n859_), .ZN(G1349gat));
  NOR3_X1   g659(.A1(new_n800_), .A2(new_n583_), .A3(new_n849_), .ZN(new_n861_));
  MUX2_X1   g660(.A(new_n251_), .B(new_n207_), .S(new_n861_), .Z(G1350gat));
  OAI211_X1 g661(.A(new_n850_), .B(new_n569_), .C1(new_n211_), .C2(new_n210_), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n814_), .A2(new_n779_), .A3(new_n849_), .ZN(new_n864_));
  INV_X1    g663(.A(G190gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n863_), .B1(new_n864_), .B2(new_n865_), .ZN(G1351gat));
  NAND3_X1  g665(.A1(new_n835_), .A2(new_n489_), .A3(new_n848_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT127), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n867_), .A2(new_n868_), .A3(new_n484_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n867_), .B2(new_n484_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n867_), .A2(new_n484_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n869_), .A2(new_n870_), .A3(new_n871_), .ZN(G1352gat));
  NAND4_X1  g671(.A1(new_n803_), .A2(new_n449_), .A3(new_n353_), .A4(new_n848_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n681_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g675(.A(KEYINPUT63), .B(G211gat), .C1(new_n874_), .C2(new_n582_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(KEYINPUT63), .B(G211gat), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n873_), .A2(new_n583_), .A3(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n877_), .A2(new_n879_), .ZN(G1354gat));
  INV_X1    g679(.A(G218gat), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n873_), .A2(new_n881_), .A3(new_n779_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n874_), .A2(new_n569_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(new_n881_), .ZN(G1355gat));
endmodule


