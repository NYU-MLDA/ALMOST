//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n633_, new_n634_, new_n635_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n869_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_;
  INV_X1    g000(.A(G141gat), .ZN(new_n202_));
  INV_X1    g001(.A(G148gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT2), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  AOI22_X1  g005(.A1(new_n204_), .A2(KEYINPUT3), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  NAND3_X1  g006(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT86), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND4_X1  g009(.A1(KEYINPUT86), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT85), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n213_), .B1(new_n204_), .B2(KEYINPUT3), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(KEYINPUT85), .A3(new_n216_), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n207_), .A2(new_n212_), .A3(new_n214_), .A4(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n218_), .A2(new_n222_), .ZN(new_n223_));
  NOR3_X1   g022(.A1(new_n220_), .A2(new_n221_), .A3(KEYINPUT1), .ZN(new_n224_));
  NAND3_X1  g023(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n204_), .A2(new_n225_), .A3(new_n206_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT84), .B1(new_n224_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n221_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(new_n229_), .A3(new_n219_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n206_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n231_), .A2(new_n215_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT84), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n230_), .A2(new_n232_), .A3(new_n233_), .A4(new_n225_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n227_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n223_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT87), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  AOI22_X1  g037(.A1(new_n222_), .A2(new_n218_), .B1(new_n227_), .B2(new_n234_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT87), .ZN(new_n240_));
  XOR2_X1   g039(.A(G127gat), .B(G134gat), .Z(new_n241_));
  XOR2_X1   g040(.A(G113gat), .B(G120gat), .Z(new_n242_));
  XOR2_X1   g041(.A(new_n241_), .B(new_n242_), .Z(new_n243_));
  NAND3_X1  g042(.A1(new_n238_), .A2(new_n240_), .A3(new_n243_), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n236_), .A2(new_n243_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G225gat), .A2(G233gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n244_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G1gat), .B(G29gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(G85gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT0), .B(G57gat), .ZN(new_n250_));
  XOR2_X1   g049(.A(new_n249_), .B(new_n250_), .Z(new_n251_));
  AND3_X1   g050(.A1(new_n244_), .A2(KEYINPUT4), .A3(new_n245_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT4), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n238_), .A2(new_n240_), .A3(new_n253_), .A4(new_n243_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n246_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n247_), .B(new_n251_), .C1(new_n252_), .C2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n244_), .A2(new_n245_), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n255_), .B(new_n254_), .C1(new_n259_), .C2(new_n253_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n251_), .B1(new_n260_), .B2(new_n247_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n258_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT23), .ZN(new_n264_));
  INV_X1    g063(.A(G183gat), .ZN(new_n265_));
  INV_X1    g064(.A(G190gat), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n264_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT24), .ZN(new_n269_));
  INV_X1    g068(.A(G169gat), .ZN(new_n270_));
  INV_X1    g069(.A(G176gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  AND3_X1   g071(.A1(new_n267_), .A2(new_n268_), .A3(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT81), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT81), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n278_), .A2(G169gat), .A3(G176gat), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n275_), .A2(new_n277_), .A3(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT26), .B(G190gat), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT80), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT25), .B(G183gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT26), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n282_), .B1(new_n285_), .B2(G190gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n273_), .B(new_n280_), .C1(new_n283_), .C2(new_n287_), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n267_), .B(new_n268_), .C1(G183gat), .C2(G190gat), .ZN(new_n289_));
  AND2_X1   g088(.A1(new_n277_), .A2(new_n279_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT22), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n291_), .A2(KEYINPUT83), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(KEYINPUT83), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n270_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT82), .B1(new_n291_), .B2(G169gat), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT82), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n296_), .A2(new_n270_), .A3(KEYINPUT22), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n295_), .A2(new_n297_), .A3(new_n271_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n289_), .B(new_n290_), .C1(new_n294_), .C2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n288_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G71gat), .B(G99gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(G43gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n300_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(new_n243_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G227gat), .A2(G233gat), .ZN(new_n305_));
  INV_X1    g104(.A(G15gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT30), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT31), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n304_), .B(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n263_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G226gat), .A2(G233gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT19), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT90), .ZN(new_n314_));
  INV_X1    g113(.A(G211gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n315_), .A2(G218gat), .ZN(new_n316_));
  INV_X1    g115(.A(G218gat), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n317_), .A2(G211gat), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n314_), .B1(new_n316_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(G211gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n315_), .A2(G218gat), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n320_), .A2(new_n321_), .A3(KEYINPUT90), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n319_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT21), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT89), .ZN(new_n325_));
  INV_X1    g124(.A(G204gat), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n325_), .B1(new_n326_), .B2(G197gat), .ZN(new_n327_));
  INV_X1    g126(.A(G197gat), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n328_), .A2(KEYINPUT89), .A3(G204gat), .ZN(new_n329_));
  AOI22_X1  g128(.A1(new_n327_), .A2(new_n329_), .B1(G197gat), .B2(new_n326_), .ZN(new_n330_));
  NOR3_X1   g129(.A1(new_n323_), .A2(new_n324_), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n327_), .A2(new_n329_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n326_), .A2(G197gat), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(new_n324_), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT88), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n335_), .B1(new_n328_), .B2(G204gat), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n326_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n328_), .A2(G204gat), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT21), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n323_), .A2(new_n334_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT91), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n323_), .A2(new_n334_), .A3(new_n340_), .A4(KEYINPUT91), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n331_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n277_), .A2(new_n279_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT22), .B(G169gat), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n346_), .B1(new_n271_), .B2(new_n347_), .ZN(new_n348_));
  AOI22_X1  g147(.A1(new_n281_), .A2(new_n284_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n349_));
  AOI22_X1  g148(.A1(new_n348_), .A2(new_n289_), .B1(new_n349_), .B2(new_n273_), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT20), .B1(new_n345_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n331_), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n324_), .A2(new_n330_), .B1(new_n319_), .B2(new_n322_), .ZN(new_n353_));
  AOI21_X1  g152(.A(KEYINPUT91), .B1(new_n353_), .B2(new_n340_), .ZN(new_n354_));
  AND4_X1   g153(.A1(KEYINPUT91), .A2(new_n323_), .A3(new_n340_), .A4(new_n334_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n352_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n356_), .A2(new_n300_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n313_), .B1(new_n351_), .B2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT96), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G8gat), .B(G36gat), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n360_), .A2(new_n361_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G64gat), .B(G92gat), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  OR3_X1    g164(.A1(new_n362_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n365_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT20), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n369_), .B1(new_n345_), .B2(new_n350_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n313_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n356_), .A2(new_n300_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n358_), .A2(new_n368_), .A3(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT27), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT99), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n368_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n366_), .A2(new_n367_), .A3(KEYINPUT99), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n352_), .B(new_n350_), .C1(new_n354_), .C2(new_n355_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT20), .ZN(new_n381_));
  INV_X1    g180(.A(new_n300_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n343_), .A2(new_n344_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n382_), .B1(new_n383_), .B2(new_n352_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n313_), .B1(new_n381_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n350_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n369_), .B1(new_n356_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n345_), .A2(new_n382_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n387_), .A2(new_n371_), .A3(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n379_), .B1(new_n385_), .B2(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n375_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n368_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n371_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n381_), .A2(new_n313_), .A3(new_n384_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n392_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT97), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n368_), .B1(new_n358_), .B2(new_n373_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT97), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n399_), .A3(new_n374_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT100), .B(KEYINPUT27), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n391_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT94), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT93), .ZN(new_n404_));
  XOR2_X1   g203(.A(KEYINPUT92), .B(KEYINPUT29), .Z(new_n405_));
  OAI21_X1  g204(.A(new_n404_), .B1(new_n239_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n405_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n236_), .A2(KEYINPUT93), .A3(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n356_), .A2(new_n406_), .A3(new_n408_), .ZN(new_n409_));
  AND2_X1   g208(.A1(G228gat), .A2(G233gat), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n345_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n238_), .A2(new_n240_), .A3(KEYINPUT29), .ZN(new_n412_));
  AOI22_X1  g211(.A1(new_n409_), .A2(new_n410_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G78gat), .B(G106gat), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n403_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n238_), .A2(new_n240_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT29), .ZN(new_n418_));
  XOR2_X1   g217(.A(G22gat), .B(G50gat), .Z(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT28), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n417_), .A2(new_n418_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n420_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n409_), .A2(new_n410_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n411_), .A2(new_n412_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n425_), .A2(new_n415_), .A3(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n415_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n428_));
  OAI22_X1  g227(.A1(new_n416_), .A2(new_n424_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n428_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n413_), .A2(new_n415_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n422_), .A2(new_n423_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .A4(new_n403_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n429_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n311_), .A2(new_n402_), .A3(new_n434_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n262_), .A2(new_n433_), .A3(new_n429_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n389_), .A2(new_n385_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n437_), .A2(KEYINPUT32), .A3(new_n368_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n368_), .A2(KEYINPUT32), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n358_), .A2(new_n373_), .A3(new_n439_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n438_), .B(new_n440_), .C1(new_n258_), .C2(new_n261_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(KEYINPUT98), .B(KEYINPUT33), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n257_), .A2(new_n442_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n260_), .A2(KEYINPUT33), .A3(new_n247_), .A4(new_n251_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n251_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n254_), .A2(new_n246_), .ZN(new_n446_));
  OAI221_X1 g245(.A(new_n445_), .B1(new_n259_), .B2(new_n246_), .C1(new_n252_), .C2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n443_), .A2(new_n444_), .A3(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n441_), .B1(new_n400_), .B2(new_n448_), .ZN(new_n449_));
  AOI22_X1  g248(.A1(new_n436_), .A2(new_n402_), .B1(new_n449_), .B2(new_n434_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n310_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n435_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(G29gat), .B(G36gat), .Z(new_n454_));
  XNOR2_X1  g253(.A(G43gat), .B(G50gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(new_n456_), .B(KEYINPUT15), .Z(new_n457_));
  XNOR2_X1  g256(.A(G15gat), .B(G22gat), .ZN(new_n458_));
  INV_X1    g257(.A(G1gat), .ZN(new_n459_));
  INV_X1    g258(.A(G8gat), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT14), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n458_), .A2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G1gat), .B(G8gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n457_), .A2(new_n464_), .ZN(new_n465_));
  OR2_X1    g264(.A1(new_n464_), .A2(new_n456_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G229gat), .A2(G233gat), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n464_), .B(new_n456_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n467_), .ZN(new_n470_));
  AOI22_X1  g269(.A1(new_n465_), .A2(new_n468_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(G113gat), .B(G141gat), .Z(new_n472_));
  XNOR2_X1  g271(.A(G169gat), .B(G197gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n471_), .A2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n471_), .A2(new_n474_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n453_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT69), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G230gat), .A2(G233gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G99gat), .A2(G106gat), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT6), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(KEYINPUT10), .B(G99gat), .Z(new_n485_));
  INV_X1    g284(.A(G106gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G85gat), .B(G92gat), .Z(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT9), .ZN(new_n489_));
  INV_X1    g288(.A(G85gat), .ZN(new_n490_));
  INV_X1    g289(.A(G92gat), .ZN(new_n491_));
  OR3_X1    g290(.A1(new_n490_), .A2(new_n491_), .A3(KEYINPUT9), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n484_), .A2(new_n487_), .A3(new_n489_), .A4(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(G99gat), .A2(G106gat), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT7), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n488_), .B1(new_n497_), .B2(new_n483_), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n498_), .A2(KEYINPUT8), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(KEYINPUT8), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n494_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G57gat), .B(G64gat), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n502_), .A2(KEYINPUT11), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(KEYINPUT11), .ZN(new_n504_));
  XOR2_X1   g303(.A(G71gat), .B(G78gat), .Z(new_n505_));
  NAND3_X1  g304(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n504_), .A2(new_n505_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n501_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT12), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n498_), .A2(KEYINPUT8), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n498_), .A2(KEYINPUT8), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n493_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n508_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n510_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT65), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n517_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n499_), .A2(KEYINPUT65), .A3(new_n500_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(new_n493_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n514_), .A2(KEYINPUT12), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(KEYINPUT66), .B1(new_n521_), .B2(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n494_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT66), .ZN(new_n526_));
  NOR3_X1   g325(.A1(new_n525_), .A2(new_n526_), .A3(new_n522_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n480_), .B(new_n516_), .C1(new_n524_), .C2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT64), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n509_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n501_), .A2(KEYINPUT64), .A3(new_n508_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n515_), .A3(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n532_), .A2(G230gat), .A3(G233gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n528_), .A2(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(KEYINPUT67), .B(KEYINPUT5), .Z(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT68), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G120gat), .B(G148gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G176gat), .B(G204gat), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n538_), .B(new_n539_), .Z(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n479_), .B1(new_n534_), .B2(new_n541_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n528_), .A2(KEYINPUT69), .A3(new_n533_), .A4(new_n540_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n534_), .A2(new_n541_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n547_), .A2(KEYINPUT13), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(KEYINPUT13), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n521_), .A2(new_n457_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G232gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT71), .ZN(new_n554_));
  XOR2_X1   g353(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT35), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT74), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n513_), .A2(new_n456_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n552_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(KEYINPUT73), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n556_), .A2(new_n557_), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n564_), .B(KEYINPUT72), .Z(new_n565_));
  AND3_X1   g364(.A1(new_n562_), .A2(new_n563_), .A3(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n562_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G190gat), .B(G218gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT75), .ZN(new_n570_));
  XOR2_X1   g369(.A(G134gat), .B(G162gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT76), .B(KEYINPUT36), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n568_), .A2(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n572_), .B(KEYINPUT36), .Z(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n577_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n579_), .A2(KEYINPUT37), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT37), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n576_), .B(KEYINPUT77), .Z(new_n582_));
  OAI21_X1  g381(.A(new_n582_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n581_), .B1(new_n575_), .B2(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n580_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n508_), .B(new_n464_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G231gat), .A2(G233gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT17), .ZN(new_n589_));
  XOR2_X1   g388(.A(G127gat), .B(G155gat), .Z(new_n590_));
  XNOR2_X1  g389(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G183gat), .B(G211gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  OR3_X1    g393(.A1(new_n588_), .A2(new_n589_), .A3(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(KEYINPUT17), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n588_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT79), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n585_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n478_), .A2(new_n551_), .A3(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT101), .Z(new_n602_));
  NAND3_X1  g401(.A1(new_n602_), .A2(new_n459_), .A3(new_n263_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT38), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n602_), .A2(KEYINPUT38), .A3(new_n459_), .A4(new_n263_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n452_), .A2(new_n579_), .ZN(new_n607_));
  NOR4_X1   g406(.A1(new_n550_), .A2(new_n607_), .A3(new_n477_), .A4(new_n598_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(G1gat), .B1(new_n609_), .B2(new_n262_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n605_), .A2(new_n606_), .A3(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT102), .ZN(G1324gat));
  INV_X1    g411(.A(KEYINPUT40), .ZN(new_n613_));
  INV_X1    g412(.A(new_n402_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n460_), .B1(new_n608_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT103), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n615_), .A2(new_n616_), .ZN(new_n618_));
  OAI21_X1  g417(.A(KEYINPUT104), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n615_), .A2(new_n616_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT104), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n615_), .A2(new_n616_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n620_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n619_), .A2(new_n623_), .A3(KEYINPUT39), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT39), .ZN(new_n625_));
  OAI211_X1 g424(.A(KEYINPUT104), .B(new_n625_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n602_), .A2(new_n460_), .A3(new_n614_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n613_), .B1(new_n624_), .B2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n619_), .A2(new_n623_), .A3(KEYINPUT39), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n630_), .A2(KEYINPUT40), .A3(new_n626_), .A4(new_n627_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n629_), .A2(new_n631_), .ZN(G1325gat));
  NAND3_X1  g431(.A1(new_n602_), .A2(new_n306_), .A3(new_n451_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n306_), .B1(new_n608_), .B2(new_n451_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT41), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(G1326gat));
  INV_X1    g435(.A(G22gat), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n429_), .A2(new_n433_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n608_), .B2(new_n638_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT42), .Z(new_n640_));
  NAND3_X1  g439(.A1(new_n602_), .A2(new_n637_), .A3(new_n638_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT105), .Z(G1327gat));
  OR2_X1    g442(.A1(new_n580_), .A2(new_n584_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n453_), .A2(new_n644_), .A3(KEYINPUT43), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n449_), .A2(new_n434_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n374_), .B1(new_n398_), .B2(KEYINPUT97), .ZN(new_n648_));
  AOI211_X1 g447(.A(new_n396_), .B(new_n368_), .C1(new_n358_), .C2(new_n373_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n401_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n391_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n638_), .A2(new_n650_), .A3(new_n651_), .A4(new_n262_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n451_), .B1(new_n647_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n435_), .ZN(new_n654_));
  OAI21_X1  g453(.A(KEYINPUT106), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT106), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n656_), .B(new_n435_), .C1(new_n450_), .C2(new_n451_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n655_), .A2(new_n657_), .A3(new_n585_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT107), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n658_), .A2(new_n659_), .A3(KEYINPUT43), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n658_), .B2(KEYINPUT43), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n646_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n599_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n550_), .A2(new_n477_), .A3(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n662_), .A2(KEYINPUT44), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(G29gat), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n262_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n662_), .A2(new_n664_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n669_));
  AOI21_X1  g468(.A(KEYINPUT108), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT108), .ZN(new_n671_));
  AOI211_X1 g470(.A(new_n671_), .B(KEYINPUT44), .C1(new_n662_), .C2(new_n664_), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n665_), .B(new_n667_), .C1(new_n670_), .C2(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n663_), .A2(new_n579_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n478_), .A2(new_n551_), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n666_), .B1(new_n676_), .B2(new_n262_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n673_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT109), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT109), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n673_), .A2(new_n680_), .A3(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(G1328gat));
  INV_X1    g481(.A(G36gat), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n675_), .A2(new_n683_), .A3(new_n614_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT45), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n665_), .A2(new_n614_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n658_), .A2(KEYINPUT43), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT107), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n658_), .A2(new_n659_), .A3(KEYINPUT43), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n645_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n664_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n669_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(new_n671_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n668_), .A2(KEYINPUT108), .A3(new_n669_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n686_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n685_), .B1(new_n695_), .B2(new_n683_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  OAI221_X1 g497(.A(new_n685_), .B1(KEYINPUT110), .B2(KEYINPUT46), .C1(new_n695_), .C2(new_n683_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1329gat));
  AND2_X1   g499(.A1(new_n451_), .A2(G43gat), .ZN(new_n701_));
  OAI211_X1 g500(.A(new_n665_), .B(new_n701_), .C1(new_n670_), .C2(new_n672_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(KEYINPUT111), .B(G43gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n703_), .B1(new_n676_), .B2(new_n310_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT47), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT47), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n702_), .A2(new_n707_), .A3(new_n704_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(G1330gat));
  AOI21_X1  g508(.A(G50gat), .B1(new_n675_), .B2(new_n638_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n665_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n711_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n638_), .A2(G50gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n710_), .B1(new_n712_), .B2(new_n713_), .ZN(G1331gat));
  INV_X1    g513(.A(new_n477_), .ZN(new_n715_));
  OR4_X1    g514(.A1(new_n715_), .A2(new_n551_), .A3(new_n599_), .A4(new_n607_), .ZN(new_n716_));
  INV_X1    g515(.A(G57gat), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n716_), .A2(new_n717_), .A3(new_n262_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n551_), .A2(new_n453_), .A3(new_n715_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n600_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n721_), .A2(KEYINPUT112), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(KEYINPUT112), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n722_), .A2(new_n263_), .A3(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n718_), .B1(new_n724_), .B2(new_n717_), .ZN(G1332gat));
  OAI21_X1  g524(.A(G64gat), .B1(new_n716_), .B2(new_n402_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT48), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n402_), .A2(G64gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(new_n720_), .B2(new_n728_), .ZN(G1333gat));
  OAI21_X1  g528(.A(G71gat), .B1(new_n716_), .B2(new_n310_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT49), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n310_), .A2(G71gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n720_), .B2(new_n732_), .ZN(G1334gat));
  OAI21_X1  g532(.A(G78gat), .B1(new_n716_), .B2(new_n434_), .ZN(new_n734_));
  XOR2_X1   g533(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n735_));
  XNOR2_X1  g534(.A(new_n734_), .B(new_n735_), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n434_), .A2(G78gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n720_), .B2(new_n737_), .ZN(G1335gat));
  NAND2_X1  g537(.A1(new_n719_), .A2(new_n674_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n490_), .B1(new_n739_), .B2(new_n262_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT114), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n551_), .A2(new_n715_), .A3(new_n663_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n662_), .A2(new_n742_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n262_), .A2(new_n490_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n741_), .B1(new_n743_), .B2(new_n744_), .ZN(G1336gat));
  INV_X1    g544(.A(new_n739_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n746_), .A2(new_n491_), .A3(new_n614_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n743_), .A2(new_n614_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(new_n491_), .ZN(G1337gat));
  AND3_X1   g548(.A1(new_n746_), .A2(new_n451_), .A3(new_n485_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n743_), .A2(new_n451_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n751_), .B2(G99gat), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n752_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n662_), .A2(new_n638_), .A3(new_n742_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n755_), .A2(KEYINPUT116), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT116), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n662_), .A2(new_n757_), .A3(new_n638_), .A4(new_n742_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(G106gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n754_), .B1(new_n756_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n755_), .A2(KEYINPUT116), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n761_), .A2(KEYINPUT52), .A3(G106gat), .A4(new_n758_), .ZN(new_n762_));
  AND4_X1   g561(.A1(new_n486_), .A2(new_n719_), .A3(new_n638_), .A4(new_n674_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT115), .Z(new_n764_));
  NAND3_X1  g563(.A1(new_n760_), .A2(new_n762_), .A3(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT53), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n760_), .A2(new_n764_), .A3(new_n767_), .A4(new_n762_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1339gat));
  NAND3_X1  g568(.A1(new_n465_), .A2(new_n466_), .A3(new_n470_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n474_), .B1(new_n469_), .B2(new_n467_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n475_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n544_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n521_), .A2(KEYINPUT66), .A3(new_n523_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n526_), .B1(new_n525_), .B2(new_n522_), .ZN(new_n777_));
  AOI22_X1  g576(.A1(new_n776_), .A2(new_n777_), .B1(new_n515_), .B2(new_n510_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT117), .B1(new_n778_), .B2(new_n480_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780_));
  OAI22_X1  g579(.A1(new_n779_), .A2(new_n780_), .B1(new_n480_), .B2(new_n778_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n528_), .A2(new_n782_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n783_), .A2(KEYINPUT55), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n541_), .B1(new_n781_), .B2(new_n784_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n775_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n778_), .A2(new_n480_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n788_), .B1(new_n783_), .B2(KEYINPUT55), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n779_), .A2(new_n780_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n540_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n786_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n773_), .B1(new_n787_), .B2(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n585_), .B1(new_n794_), .B2(KEYINPUT58), .ZN(new_n795_));
  INV_X1    g594(.A(new_n773_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n774_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n785_), .A2(new_n786_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n796_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT58), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n579_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT56), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT118), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n803_), .B1(new_n791_), .B2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n785_), .A2(KEYINPUT118), .A3(KEYINPUT56), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n477_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n805_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n546_), .A2(new_n772_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n802_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  OAI22_X1  g609(.A1(new_n795_), .A2(new_n801_), .B1(new_n810_), .B2(KEYINPUT57), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n808_), .A2(new_n809_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n579_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT57), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n598_), .B1(new_n811_), .B2(new_n815_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n600_), .A2(new_n549_), .A3(new_n477_), .A4(new_n548_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(KEYINPUT54), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n614_), .A2(new_n638_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n821_), .A2(new_n263_), .A3(new_n451_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n820_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(G113gat), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n715_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT59), .ZN(new_n826_));
  INV_X1    g625(.A(new_n822_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n826_), .B1(new_n819_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT122), .ZN(new_n829_));
  XOR2_X1   g628(.A(new_n817_), .B(KEYINPUT54), .Z(new_n830_));
  INV_X1    g629(.A(KEYINPUT121), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n811_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n813_), .A2(new_n814_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n794_), .A2(KEYINPUT58), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n799_), .A2(new_n800_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n834_), .A2(new_n835_), .A3(new_n585_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n833_), .A2(new_n836_), .A3(KEYINPUT121), .ZN(new_n837_));
  INV_X1    g636(.A(new_n815_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n832_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n830_), .B1(new_n839_), .B2(new_n599_), .ZN(new_n840_));
  OR2_X1    g639(.A1(new_n822_), .A2(KEYINPUT120), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n822_), .A2(KEYINPUT120), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n841_), .A2(new_n826_), .A3(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n829_), .B1(new_n840_), .B2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n815_), .B1(new_n811_), .B2(new_n831_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n663_), .B1(new_n846_), .B2(new_n837_), .ZN(new_n847_));
  OAI211_X1 g646(.A(KEYINPUT122), .B(new_n843_), .C1(new_n847_), .C2(new_n830_), .ZN(new_n848_));
  AOI211_X1 g647(.A(new_n477_), .B(new_n828_), .C1(new_n845_), .C2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n825_), .B1(new_n849_), .B2(new_n824_), .ZN(G1340gat));
  INV_X1    g649(.A(G120gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n551_), .B2(KEYINPUT60), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n823_), .B(new_n852_), .C1(KEYINPUT60), .C2(new_n851_), .ZN(new_n853_));
  AOI211_X1 g652(.A(new_n551_), .B(new_n828_), .C1(new_n845_), .C2(new_n848_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n854_), .B2(new_n851_), .ZN(G1341gat));
  INV_X1    g654(.A(G127gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n823_), .A2(new_n856_), .A3(new_n663_), .ZN(new_n857_));
  AOI211_X1 g656(.A(new_n598_), .B(new_n828_), .C1(new_n845_), .C2(new_n848_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n856_), .ZN(G1342gat));
  AOI21_X1  g658(.A(G134gat), .B1(new_n823_), .B2(new_n802_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n828_), .B1(new_n845_), .B2(new_n848_), .ZN(new_n861_));
  XOR2_X1   g660(.A(KEYINPUT123), .B(G134gat), .Z(new_n862_));
  NOR2_X1   g661(.A1(new_n644_), .A2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n860_), .B1(new_n861_), .B2(new_n863_), .ZN(G1343gat));
  NOR3_X1   g663(.A1(new_n434_), .A2(new_n451_), .A3(new_n262_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n819_), .A2(new_n402_), .A3(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n477_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(new_n202_), .ZN(G1344gat));
  NOR2_X1   g667(.A1(new_n866_), .A2(new_n551_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(new_n203_), .ZN(G1345gat));
  NOR2_X1   g669(.A1(new_n866_), .A2(new_n599_), .ZN(new_n871_));
  XOR2_X1   g670(.A(KEYINPUT61), .B(G155gat), .Z(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(G1346gat));
  OAI21_X1  g672(.A(G162gat), .B1(new_n866_), .B2(new_n644_), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n579_), .A2(G162gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n866_), .B2(new_n875_), .ZN(G1347gat));
  NAND2_X1  g675(.A1(new_n614_), .A2(new_n311_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(new_n638_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(KEYINPUT124), .B1(new_n840_), .B2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n881_), .B(new_n878_), .C1(new_n847_), .C2(new_n830_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n715_), .A2(new_n347_), .ZN(new_n885_));
  XOR2_X1   g684(.A(new_n885_), .B(KEYINPUT125), .Z(new_n886_));
  OAI211_X1 g685(.A(new_n715_), .B(new_n878_), .C1(new_n847_), .C2(new_n830_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n888_));
  AND3_X1   g687(.A1(new_n887_), .A2(new_n888_), .A3(G169gat), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n888_), .B1(new_n887_), .B2(G169gat), .ZN(new_n890_));
  OAI22_X1  g689(.A1(new_n884_), .A2(new_n886_), .B1(new_n889_), .B2(new_n890_), .ZN(G1348gat));
  NAND2_X1  g690(.A1(new_n883_), .A2(new_n550_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n820_), .A2(new_n638_), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n550_), .A2(G176gat), .A3(new_n614_), .A4(new_n311_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n892_), .A2(new_n271_), .B1(new_n893_), .B2(new_n895_), .ZN(G1349gat));
  NOR2_X1   g695(.A1(new_n877_), .A2(new_n599_), .ZN(new_n897_));
  AOI21_X1  g696(.A(G183gat), .B1(new_n893_), .B2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n598_), .A2(new_n284_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n883_), .B2(new_n899_), .ZN(G1350gat));
  NAND3_X1  g699(.A1(new_n883_), .A2(new_n281_), .A3(new_n802_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n644_), .B1(new_n880_), .B2(new_n882_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n266_), .B2(new_n902_), .ZN(G1351gat));
  AND4_X1   g702(.A1(new_n436_), .A2(new_n819_), .A3(new_n614_), .A4(new_n310_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n715_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n550_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g707(.A1(new_n904_), .A2(new_n595_), .A3(new_n597_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(KEYINPUT63), .B(G211gat), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n911_), .B1(new_n909_), .B2(new_n912_), .ZN(G1354gat));
  NAND2_X1  g712(.A1(new_n904_), .A2(new_n802_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(KEYINPUT126), .B(G218gat), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n644_), .A2(new_n915_), .ZN(new_n916_));
  AOI22_X1  g715(.A1(new_n914_), .A2(new_n915_), .B1(new_n904_), .B2(new_n916_), .ZN(G1355gat));
endmodule


