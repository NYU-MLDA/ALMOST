//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 0 0 1 0 1 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 0 1 0 1 0 1 0 1 1 1 0 0 0 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n855_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n928_;
  XNOR2_X1  g000(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(KEYINPUT23), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT80), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n206_), .B(KEYINPUT77), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT23), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT22), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(KEYINPUT79), .A3(G169gat), .ZN(new_n216_));
  INV_X1    g015(.A(G176gat), .ZN(new_n217_));
  AND2_X1   g016(.A1(KEYINPUT79), .A2(G169gat), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n216_), .B(new_n217_), .C1(new_n215_), .C2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n213_), .A2(new_n214_), .A3(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(G197gat), .B(G204gat), .Z(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT21), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G211gat), .B(G218gat), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G197gat), .B(G204gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT21), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n222_), .A2(new_n227_), .A3(new_n223_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n224_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n209_), .A2(KEYINPUT23), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT78), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n206_), .A2(KEYINPUT23), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT78), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n234_), .B1(new_n209_), .B2(KEYINPUT23), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n232_), .A2(new_n235_), .ZN(new_n236_));
  OR2_X1    g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n237_), .A2(KEYINPUT24), .A3(new_n214_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n238_), .B1(KEYINPUT24), .B2(new_n237_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT26), .B(G190gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT25), .B(G183gat), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n239_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n236_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n220_), .A2(new_n230_), .A3(new_n243_), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n244_), .A2(KEYINPUT20), .ZN(new_n245_));
  XOR2_X1   g044(.A(new_n241_), .B(KEYINPUT91), .Z(new_n246_));
  AOI21_X1  g045(.A(new_n239_), .B1(new_n246_), .B2(new_n240_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(new_n211_), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n236_), .A2(new_n212_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT22), .B(G169gat), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n214_), .B1(new_n251_), .B2(G176gat), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n248_), .B1(new_n249_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(new_n229_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n205_), .B1(new_n245_), .B2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n248_), .B(new_n230_), .C1(new_n249_), .C2(new_n252_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n220_), .A2(new_n243_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(new_n229_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n257_), .A2(new_n259_), .A3(KEYINPUT20), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n260_), .A2(new_n204_), .ZN(new_n261_));
  XOR2_X1   g060(.A(G8gat), .B(G36gat), .Z(new_n262_));
  XNOR2_X1  g061(.A(G64gat), .B(G92gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n256_), .A2(new_n261_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT27), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n260_), .A2(new_n204_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n245_), .A2(new_n254_), .A3(new_n205_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n267_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NOR3_X1   g072(.A1(new_n269_), .A2(new_n270_), .A3(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n260_), .A2(new_n204_), .ZN(new_n275_));
  OR4_X1    g074(.A1(KEYINPUT93), .A2(new_n275_), .A3(new_n255_), .A4(new_n266_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n266_), .B1(new_n275_), .B2(new_n255_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n268_), .A2(KEYINPUT93), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT98), .B1(new_n279_), .B2(KEYINPUT27), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT98), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n276_), .A2(new_n278_), .A3(new_n281_), .A4(new_n270_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n274_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(G141gat), .B(G148gat), .Z(new_n284_));
  NAND2_X1  g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT83), .B1(new_n285_), .B2(KEYINPUT1), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(KEYINPUT1), .ZN(new_n287_));
  OR2_X1    g086(.A1(G155gat), .A2(G162gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n286_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  NOR3_X1   g088(.A1(new_n285_), .A2(KEYINPUT83), .A3(KEYINPUT1), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n284_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(G141gat), .A2(G148gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT3), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G141gat), .A2(G148gat), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT2), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n294_), .A2(new_n297_), .A3(new_n298_), .A4(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n300_), .A2(new_n285_), .A3(new_n288_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n291_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT29), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n229_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n304_), .B1(G228gat), .B2(G233gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT85), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n304_), .A2(G228gat), .A3(G233gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT86), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G78gat), .B(G106gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n310_), .B(KEYINPUT87), .Z(new_n311_));
  XOR2_X1   g110(.A(new_n311_), .B(KEYINPUT88), .Z(new_n312_));
  XNOR2_X1  g111(.A(new_n309_), .B(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n302_), .A2(KEYINPUT29), .ZN(new_n314_));
  XOR2_X1   g113(.A(G22gat), .B(G50gat), .Z(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(KEYINPUT84), .B(KEYINPUT28), .Z(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n313_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n311_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n309_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n306_), .A2(new_n308_), .A3(new_n312_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n321_), .A2(new_n322_), .A3(new_n318_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT89), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n321_), .A2(KEYINPUT89), .A3(new_n322_), .A4(new_n318_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n319_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G127gat), .B(G134gat), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n330_), .A2(KEYINPUT82), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(KEYINPUT82), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G113gat), .B(G120gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n302_), .A2(KEYINPUT94), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G225gat), .A2(G233gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n339_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT4), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n335_), .A2(new_n342_), .A3(new_n302_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n341_), .B(new_n343_), .C1(new_n337_), .C2(new_n342_), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n340_), .A2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G1gat), .B(G29gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(G85gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT0), .B(G57gat), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n347_), .B(new_n348_), .Z(new_n349_));
  OR2_X1    g148(.A1(new_n345_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n340_), .A2(new_n344_), .A3(new_n349_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n335_), .B(KEYINPUT31), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(G99gat), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n258_), .B(KEYINPUT30), .ZN(new_n356_));
  XOR2_X1   g155(.A(KEYINPUT81), .B(G43gat), .Z(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G227gat), .A2(G233gat), .ZN(new_n359_));
  INV_X1    g158(.A(G15gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(G71gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n358_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n358_), .A2(new_n363_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n355_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n366_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n368_), .A2(new_n354_), .A3(new_n364_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n352_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n283_), .A2(new_n329_), .A3(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n352_), .B1(new_n319_), .B2(new_n327_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n256_), .A2(new_n261_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n267_), .A2(KEYINPUT32), .ZN(new_n374_));
  OR3_X1    g173(.A1(new_n373_), .A2(KEYINPUT97), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n271_), .A2(new_n272_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n374_), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT97), .B1(new_n373_), .B2(new_n374_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n352_), .A2(new_n375_), .A3(new_n377_), .A4(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n349_), .B1(new_n338_), .B2(new_n341_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n380_), .A2(KEYINPUT96), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(KEYINPUT96), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n343_), .B1(new_n337_), .B2(new_n342_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n382_), .B1(new_n341_), .B2(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n279_), .B1(new_n381_), .B2(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(KEYINPUT95), .A2(KEYINPUT33), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n351_), .B(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n379_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n388_));
  AOI22_X1  g187(.A1(new_n283_), .A2(new_n372_), .B1(new_n388_), .B2(new_n329_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n367_), .A2(new_n369_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n371_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G15gat), .B(G22gat), .ZN(new_n392_));
  INV_X1    g191(.A(G1gat), .ZN(new_n393_));
  INV_X1    g192(.A(G8gat), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT14), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n392_), .A2(new_n395_), .ZN(new_n396_));
  XOR2_X1   g195(.A(G1gat), .B(G8gat), .Z(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n398_), .B(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G231gat), .A2(G233gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G71gat), .B(G78gat), .ZN(new_n404_));
  INV_X1    g203(.A(G64gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(G57gat), .ZN(new_n406_));
  INV_X1    g205(.A(G57gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(G64gat), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n404_), .A2(KEYINPUT11), .A3(new_n406_), .A4(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n406_), .A2(new_n408_), .A3(KEYINPUT11), .ZN(new_n410_));
  INV_X1    g209(.A(G78gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(G71gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n362_), .A2(G78gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(KEYINPUT11), .B1(new_n406_), .B2(new_n408_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n409_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n403_), .B(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G127gat), .B(G155gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT16), .ZN(new_n420_));
  XOR2_X1   g219(.A(G183gat), .B(G211gat), .Z(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT17), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n423_), .A2(KEYINPUT64), .ZN(new_n424_));
  OR2_X1    g223(.A1(new_n418_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT64), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n423_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n422_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT17), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n429_), .A2(KEYINPUT76), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(KEYINPUT76), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n418_), .A2(new_n427_), .A3(new_n430_), .A4(new_n431_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n425_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G190gat), .B(G218gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G134gat), .B(G162gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n437_), .A2(KEYINPUT36), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G232gat), .A2(G233gat), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT34), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT35), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT71), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT15), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G43gat), .B(G50gat), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G29gat), .B(G36gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(G29gat), .B(G36gat), .Z(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n447_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n450_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n453_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n446_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n450_), .A2(new_n452_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n453_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n450_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(KEYINPUT15), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n456_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G99gat), .A2(G106gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT6), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT6), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n465_), .A2(G99gat), .A3(G106gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  OR2_X1    g266(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n468_));
  INV_X1    g267(.A(G106gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n468_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(G85gat), .ZN(new_n472_));
  INV_X1    g271(.A(G92gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G85gat), .A2(G92gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(KEYINPUT9), .A3(new_n475_), .ZN(new_n476_));
  OR2_X1    g275(.A1(new_n475_), .A2(KEYINPUT9), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n467_), .A2(new_n471_), .A3(new_n476_), .A4(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n474_), .A2(new_n475_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT7), .ZN(new_n480_));
  INV_X1    g279(.A(G99gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n480_), .A2(new_n481_), .A3(new_n469_), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  AOI211_X1 g283(.A(KEYINPUT8), .B(new_n479_), .C1(new_n484_), .C2(new_n467_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT8), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n467_), .A2(new_n483_), .A3(new_n482_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n479_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n486_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n478_), .B1(new_n485_), .B2(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n445_), .B1(new_n462_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n478_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n464_), .A2(new_n466_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n482_), .A2(new_n483_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n488_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT8), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n487_), .A2(new_n486_), .A3(new_n488_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n492_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n454_), .A2(new_n455_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n491_), .A2(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n442_), .A2(new_n443_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT72), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n502_), .A2(KEYINPUT72), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n501_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n491_), .A2(KEYINPUT72), .A3(new_n502_), .A4(new_n500_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n439_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT73), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n437_), .B(KEYINPUT36), .Z(new_n510_));
  NAND3_X1  g309(.A1(new_n505_), .A2(new_n506_), .A3(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n508_), .A2(new_n509_), .A3(new_n511_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n505_), .A2(KEYINPUT73), .A3(new_n506_), .A4(new_n510_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n391_), .A2(new_n434_), .A3(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT13), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n516_), .A2(KEYINPUT68), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n516_), .A2(KEYINPUT68), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G120gat), .B(G148gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT5), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G176gat), .B(G204gat), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n520_), .B(new_n521_), .Z(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT65), .B(KEYINPUT12), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n417_), .A2(KEYINPUT64), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n409_), .B(new_n426_), .C1(new_n415_), .C2(new_n416_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n523_), .B1(new_n498_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G230gat), .A2(G233gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n498_), .A2(new_n526_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT11), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n407_), .A2(G64gat), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n405_), .A2(G57gat), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n530_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n533_), .A2(new_n410_), .A3(new_n414_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n534_), .A2(KEYINPUT12), .A3(new_n409_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n490_), .A2(new_n536_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n527_), .A2(new_n528_), .A3(new_n529_), .A4(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT66), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n529_), .A2(new_n537_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n541_), .A2(KEYINPUT66), .A3(new_n528_), .A4(new_n527_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n525_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n426_), .B1(new_n534_), .B2(new_n409_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n490_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n528_), .B1(new_n547_), .B2(new_n529_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n522_), .B1(new_n543_), .B2(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n548_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n522_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n549_), .A2(KEYINPUT67), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT67), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n550_), .A2(new_n551_), .ZN(new_n555_));
  AOI211_X1 g354(.A(new_n548_), .B(new_n522_), .C1(new_n540_), .C2(new_n542_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n554_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  AOI211_X1 g356(.A(new_n517_), .B(new_n518_), .C1(new_n553_), .C2(new_n557_), .ZN(new_n558_));
  AND4_X1   g357(.A1(KEYINPUT68), .A2(new_n553_), .A3(new_n557_), .A4(new_n516_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n401_), .A2(new_n499_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n398_), .B(new_n399_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n499_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G229gat), .A2(G233gat), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n562_), .A2(new_n462_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n567_), .B1(new_n401_), .B2(new_n499_), .ZN(new_n569_));
  AOI22_X1  g368(.A1(new_n565_), .A2(new_n567_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(G113gat), .B(G141gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(G169gat), .B(G197gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n570_), .B(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n560_), .A2(new_n574_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n575_), .A2(KEYINPUT99), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(KEYINPUT99), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n515_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n352_), .ZN(new_n580_));
  OAI21_X1  g379(.A(G1gat), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT38), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n391_), .A2(new_n574_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT37), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n511_), .A2(new_n509_), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n584_), .B(new_n513_), .C1(new_n585_), .C2(new_n507_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n508_), .A2(KEYINPUT37), .A3(new_n511_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n588_), .A2(new_n433_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n583_), .A2(new_n589_), .A3(new_n560_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(new_n393_), .A3(new_n352_), .ZN(new_n591_));
  AND3_X1   g390(.A1(new_n591_), .A2(KEYINPUT100), .A3(new_n582_), .ZN(new_n592_));
  AOI21_X1  g391(.A(KEYINPUT100), .B1(new_n591_), .B2(new_n582_), .ZN(new_n593_));
  OAI221_X1 g392(.A(new_n581_), .B1(new_n582_), .B2(new_n591_), .C1(new_n592_), .C2(new_n593_), .ZN(G1324gat));
  INV_X1    g393(.A(new_n283_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n590_), .A2(new_n394_), .A3(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n515_), .A2(new_n595_), .A3(new_n578_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT39), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n597_), .A2(new_n598_), .A3(G8gat), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n598_), .B1(new_n597_), .B2(G8gat), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n596_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g401(.A1(new_n515_), .A2(new_n390_), .A3(new_n578_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(G15gat), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n604_), .A2(KEYINPUT101), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(KEYINPUT101), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(KEYINPUT41), .A3(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n590_), .A2(new_n360_), .A3(new_n390_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(KEYINPUT41), .B1(new_n605_), .B2(new_n606_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n609_), .A2(new_n610_), .ZN(G1326gat));
  OAI21_X1  g410(.A(G22gat), .B1(new_n579_), .B2(new_n329_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT42), .ZN(new_n613_));
  INV_X1    g412(.A(G22gat), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n590_), .A2(new_n614_), .A3(new_n328_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(G1327gat));
  INV_X1    g415(.A(new_n560_), .ZN(new_n617_));
  NOR3_X1   g416(.A1(new_n617_), .A2(new_n434_), .A3(new_n514_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n583_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(G29gat), .B1(new_n620_), .B2(new_n352_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(KEYINPUT102), .A2(KEYINPUT43), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n283_), .A2(new_n372_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n388_), .A2(new_n329_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n390_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n371_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n588_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(KEYINPUT102), .A2(KEYINPUT43), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n623_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT103), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(KEYINPUT43), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n632_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n631_), .B(new_n371_), .C1(new_n389_), .C2(new_n390_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n633_), .A2(new_n634_), .A3(new_n588_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n630_), .A2(new_n635_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n576_), .A2(new_n433_), .A3(new_n577_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n636_), .A2(KEYINPUT104), .A3(KEYINPUT44), .A4(new_n637_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n630_), .A2(new_n635_), .A3(KEYINPUT44), .A4(new_n637_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT104), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n638_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n630_), .A2(new_n635_), .A3(new_n637_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT44), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n642_), .A2(new_n645_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n352_), .A2(G29gat), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n621_), .B1(new_n646_), .B2(new_n647_), .ZN(G1328gat));
  INV_X1    g447(.A(KEYINPUT46), .ZN(new_n649_));
  INV_X1    g448(.A(G36gat), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n283_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n642_), .B2(new_n651_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n583_), .A2(new_n650_), .A3(new_n595_), .A4(new_n618_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT45), .Z(new_n654_));
  OAI21_X1  g453(.A(new_n649_), .B1(new_n652_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n654_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n645_), .A2(new_n595_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n657_), .B1(new_n641_), .B2(new_n638_), .ZN(new_n658_));
  OAI211_X1 g457(.A(KEYINPUT46), .B(new_n656_), .C1(new_n658_), .C2(new_n650_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n655_), .A2(new_n659_), .ZN(G1329gat));
  AND2_X1   g459(.A1(new_n390_), .A2(G43gat), .ZN(new_n661_));
  INV_X1    g460(.A(new_n641_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n639_), .A2(new_n640_), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n645_), .B(new_n661_), .C1(new_n662_), .C2(new_n663_), .ZN(new_n664_));
  XOR2_X1   g463(.A(KEYINPUT105), .B(G43gat), .Z(new_n665_));
  INV_X1    g464(.A(new_n390_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n619_), .B2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT106), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n664_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT47), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT47), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n664_), .A2(new_n668_), .A3(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(G1330gat));
  OR3_X1    g472(.A1(new_n619_), .A2(G50gat), .A3(new_n329_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n329_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n675_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n676_), .A2(KEYINPUT107), .A3(G50gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT107), .B1(new_n676_), .B2(G50gat), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n674_), .B1(new_n677_), .B2(new_n678_), .ZN(G1331gat));
  INV_X1    g478(.A(new_n574_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n391_), .A2(new_n680_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n681_), .A2(new_n589_), .A3(new_n617_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n682_), .A2(new_n407_), .A3(new_n352_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n560_), .A2(new_n574_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n515_), .A2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G57gat), .B1(new_n685_), .B2(new_n580_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n683_), .A2(new_n686_), .ZN(G1332gat));
  NAND3_X1  g486(.A1(new_n682_), .A2(new_n405_), .A3(new_n595_), .ZN(new_n688_));
  OAI21_X1  g487(.A(G64gat), .B1(new_n685_), .B2(new_n283_), .ZN(new_n689_));
  XOR2_X1   g488(.A(KEYINPUT108), .B(KEYINPUT48), .Z(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n689_), .A2(new_n691_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n688_), .B1(new_n692_), .B2(new_n693_), .ZN(G1333gat));
  OAI21_X1  g493(.A(G71gat), .B1(new_n685_), .B2(new_n666_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT49), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n682_), .A2(new_n362_), .A3(new_n390_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1334gat));
  OAI21_X1  g497(.A(G78gat), .B1(new_n685_), .B2(new_n329_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT50), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n682_), .A2(new_n411_), .A3(new_n328_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1335gat));
  NOR3_X1   g501(.A1(new_n560_), .A2(new_n434_), .A3(new_n514_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n681_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n704_), .A2(new_n472_), .A3(new_n352_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n636_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n684_), .A2(new_n433_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n706_), .A2(new_n580_), .A3(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n705_), .B1(new_n708_), .B2(new_n472_), .ZN(G1336gat));
  NAND3_X1  g508(.A1(new_n704_), .A2(new_n473_), .A3(new_n595_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n706_), .A2(new_n283_), .A3(new_n707_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n710_), .B1(new_n711_), .B2(new_n473_), .ZN(G1337gat));
  NAND4_X1  g511(.A1(new_n704_), .A2(new_n390_), .A3(new_n468_), .A4(new_n470_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n706_), .A2(new_n666_), .A3(new_n707_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n713_), .B1(new_n714_), .B2(new_n481_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g515(.A1(new_n636_), .A2(new_n328_), .A3(new_n433_), .A4(new_n684_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n717_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n681_), .A2(new_n469_), .A3(new_n328_), .A4(new_n703_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT109), .Z(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT52), .B1(new_n717_), .B2(G106gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT53), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n722_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT53), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n724_), .A2(new_n725_), .A3(new_n718_), .A4(new_n720_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n723_), .A2(new_n726_), .ZN(G1339gat));
  NAND2_X1  g526(.A1(new_n574_), .A2(new_n552_), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT55), .B1(new_n540_), .B2(new_n542_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n529_), .A2(new_n537_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n523_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n546_), .B2(new_n490_), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n528_), .A2(KEYINPUT111), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n730_), .A2(new_n732_), .A3(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(KEYINPUT55), .B1(G230gat), .B2(G233gat), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n527_), .A2(new_n529_), .A3(new_n537_), .A4(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n734_), .B1(new_n733_), .B2(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n522_), .B1(new_n729_), .B2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT56), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n739_), .A2(KEYINPUT112), .A3(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT112), .B1(new_n739_), .B2(new_n740_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  OAI211_X1 g542(.A(KEYINPUT56), .B(new_n522_), .C1(new_n729_), .C2(new_n738_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT113), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n744_), .B(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n728_), .B1(new_n743_), .B2(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n573_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n568_), .A2(new_n561_), .A3(new_n567_), .ZN(new_n749_));
  AOI22_X1  g548(.A1(new_n570_), .A2(new_n573_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n553_), .A2(new_n557_), .A3(new_n750_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n514_), .B1(new_n747_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT57), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n750_), .A2(new_n552_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n739_), .A2(new_n740_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n755_), .B2(new_n744_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n588_), .B1(new_n756_), .B2(KEYINPUT58), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT58), .ZN(new_n758_));
  AOI211_X1 g557(.A(new_n758_), .B(new_n754_), .C1(new_n755_), .C2(new_n744_), .ZN(new_n759_));
  OAI21_X1  g558(.A(KEYINPUT114), .B1(new_n757_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n754_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n540_), .A2(new_n542_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT55), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n737_), .A2(new_n733_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n541_), .A2(new_n527_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(new_n733_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n764_), .A2(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(KEYINPUT56), .B1(new_n768_), .B2(new_n522_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n744_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n761_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n758_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n756_), .A2(KEYINPUT58), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n772_), .A2(new_n773_), .A3(new_n588_), .A4(new_n774_), .ZN(new_n775_));
  AOI22_X1  g574(.A1(new_n752_), .A2(new_n753_), .B1(new_n760_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n755_), .A2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n739_), .A2(KEYINPUT112), .A3(new_n740_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n744_), .A2(KEYINPUT113), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n768_), .A2(new_n745_), .A3(KEYINPUT56), .A4(new_n522_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n778_), .A2(new_n779_), .A3(new_n780_), .A4(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n728_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n751_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n514_), .A2(KEYINPUT57), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT115), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n787_));
  INV_X1    g586(.A(new_n785_), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n787_), .B(new_n788_), .C1(new_n747_), .C2(new_n751_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n786_), .A2(new_n789_), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n776_), .A2(KEYINPUT116), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT116), .B1(new_n776_), .B2(new_n790_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n791_), .A2(new_n792_), .A3(new_n434_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n560_), .A2(new_n680_), .A3(new_n589_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(KEYINPUT110), .B(KEYINPUT54), .ZN(new_n795_));
  XOR2_X1   g594(.A(new_n794_), .B(new_n795_), .Z(new_n796_));
  OAI21_X1  g595(.A(KEYINPUT117), .B1(new_n793_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n786_), .A2(new_n789_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n760_), .A2(new_n775_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n514_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n753_), .B1(new_n784_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n798_), .B1(new_n799_), .B2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n776_), .A2(new_n790_), .A3(KEYINPUT116), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(new_n433_), .A3(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT117), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n794_), .B(new_n795_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n806_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n797_), .A2(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n283_), .A2(new_n329_), .A3(new_n352_), .A4(new_n390_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(KEYINPUT118), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n810_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(G113gat), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n814_), .A2(new_n815_), .A3(new_n574_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n757_), .A2(new_n759_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n817_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n434_), .B1(new_n818_), .B2(new_n790_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT119), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n808_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n823_), .A2(KEYINPUT59), .A3(new_n813_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n776_), .A2(new_n790_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n434_), .B1(new_n825_), .B2(new_n798_), .ZN(new_n826_));
  AOI211_X1 g625(.A(KEYINPUT117), .B(new_n796_), .C1(new_n826_), .C2(new_n805_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n807_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n812_), .ZN(new_n830_));
  AOI211_X1 g629(.A(new_n680_), .B(new_n824_), .C1(new_n830_), .C2(KEYINPUT59), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n816_), .B1(new_n831_), .B2(new_n815_), .ZN(G1340gat));
  INV_X1    g631(.A(G120gat), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n833_), .B1(new_n560_), .B2(KEYINPUT60), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n814_), .B(new_n834_), .C1(KEYINPUT60), .C2(new_n833_), .ZN(new_n835_));
  AOI211_X1 g634(.A(new_n560_), .B(new_n824_), .C1(new_n830_), .C2(KEYINPUT59), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(new_n833_), .ZN(G1341gat));
  NAND3_X1  g636(.A1(new_n829_), .A2(new_n434_), .A3(new_n812_), .ZN(new_n838_));
  INV_X1    g637(.A(G127gat), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT120), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n838_), .A2(KEYINPUT120), .A3(new_n839_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n824_), .B1(new_n830_), .B2(KEYINPUT59), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n433_), .A2(new_n839_), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n842_), .A2(new_n843_), .B1(new_n844_), .B2(new_n845_), .ZN(G1342gat));
  AOI21_X1  g645(.A(G134gat), .B1(new_n814_), .B2(new_n801_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n588_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT121), .B(G134gat), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n847_), .B1(new_n844_), .B2(new_n850_), .ZN(G1343gat));
  NOR4_X1   g650(.A1(new_n595_), .A2(new_n390_), .A3(new_n580_), .A4(new_n329_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n829_), .A2(new_n574_), .A3(new_n852_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g653(.A1(new_n829_), .A2(new_n617_), .A3(new_n852_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g655(.A1(new_n829_), .A2(new_n434_), .A3(new_n852_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(KEYINPUT61), .B(G155gat), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(G1346gat));
  NAND4_X1  g658(.A1(new_n797_), .A2(new_n588_), .A3(new_n809_), .A4(new_n852_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(G162gat), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n514_), .A2(G162gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n829_), .A2(new_n852_), .A3(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n861_), .A2(new_n863_), .A3(KEYINPUT122), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1347gat));
  INV_X1    g667(.A(new_n823_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n283_), .A2(new_n666_), .A3(new_n352_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n870_), .A2(new_n329_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n873_), .A2(new_n574_), .A3(new_n250_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n870_), .A2(new_n574_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(KEYINPUT123), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n329_), .ZN(new_n877_));
  OAI21_X1  g676(.A(G169gat), .B1(new_n823_), .B2(new_n877_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n878_), .A2(KEYINPUT62), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(KEYINPUT62), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n874_), .B1(new_n879_), .B2(new_n880_), .ZN(G1348gat));
  OAI211_X1 g680(.A(new_n617_), .B(new_n871_), .C1(new_n821_), .C2(new_n822_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n217_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(KEYINPUT124), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n810_), .A2(KEYINPUT125), .A3(new_n328_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT125), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n886_), .B1(new_n829_), .B2(new_n329_), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n885_), .A2(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n870_), .A2(G176gat), .A3(new_n617_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n884_), .B1(new_n888_), .B2(new_n890_), .ZN(G1349gat));
  OR3_X1    g690(.A1(new_n872_), .A2(new_n246_), .A3(new_n433_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n434_), .B(new_n870_), .C1(new_n885_), .C2(new_n887_), .ZN(new_n894_));
  INV_X1    g693(.A(G183gat), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n894_), .B2(new_n895_), .ZN(G1350gat));
  NAND3_X1  g695(.A1(new_n873_), .A2(new_n240_), .A3(new_n801_), .ZN(new_n897_));
  OAI21_X1  g696(.A(G190gat), .B1(new_n872_), .B2(new_n848_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n898_), .A2(KEYINPUT126), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n898_), .A2(KEYINPUT126), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n897_), .B1(new_n899_), .B2(new_n900_), .ZN(G1351gat));
  NOR4_X1   g700(.A1(new_n283_), .A2(new_n329_), .A3(new_n352_), .A4(new_n390_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n797_), .A2(new_n809_), .A3(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(KEYINPUT127), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT127), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n797_), .A2(new_n905_), .A3(new_n809_), .A4(new_n902_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(G197gat), .B1(new_n907_), .B2(new_n574_), .ZN(new_n908_));
  INV_X1    g707(.A(G197gat), .ZN(new_n909_));
  AOI211_X1 g708(.A(new_n909_), .B(new_n680_), .C1(new_n904_), .C2(new_n906_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n908_), .A2(new_n910_), .ZN(G1352gat));
  AOI21_X1  g710(.A(new_n905_), .B1(new_n829_), .B2(new_n902_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n906_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n617_), .B1(new_n912_), .B2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(G204gat), .ZN(new_n915_));
  INV_X1    g714(.A(G204gat), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n907_), .A2(new_n916_), .A3(new_n617_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n915_), .A2(new_n917_), .ZN(G1353gat));
  NOR2_X1   g717(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n433_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n920_), .B1(new_n907_), .B2(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n921_), .ZN(new_n923_));
  AOI211_X1 g722(.A(new_n919_), .B(new_n923_), .C1(new_n904_), .C2(new_n906_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n922_), .A2(new_n924_), .ZN(G1354gat));
  INV_X1    g724(.A(G218gat), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n907_), .A2(new_n926_), .A3(new_n801_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n848_), .B1(new_n904_), .B2(new_n906_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n927_), .B1(new_n926_), .B2(new_n928_), .ZN(G1355gat));
endmodule


