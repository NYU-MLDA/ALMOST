//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n572_, new_n573_, new_n574_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n805_, new_n806_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n814_, new_n816_,
    new_n818_, new_n819_, new_n820_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n866_, new_n868_, new_n869_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_;
  XNOR2_X1  g000(.A(KEYINPUT18), .B(G64gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G92gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G8gat), .B(G36gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  AND2_X1   g004(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n206_));
  AND2_X1   g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT22), .B(G169gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT89), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT79), .B(G176gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n207_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT90), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT23), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n215_), .B1(G183gat), .B2(G190gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT24), .ZN(new_n219_));
  NOR3_X1   g018(.A1(new_n207_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT25), .B(G183gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT26), .B(G190gat), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n220_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT88), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n218_), .A2(new_n219_), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n215_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n217_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(G197gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT85), .B(G197gat), .ZN(new_n230_));
  MUX2_X1   g029(.A(new_n229_), .B(new_n230_), .S(G204gat), .Z(new_n231_));
  INV_X1    g030(.A(KEYINPUT21), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G211gat), .B(G218gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G197gat), .A2(G204gat), .ZN(new_n235_));
  OAI211_X1 g034(.A(KEYINPUT21), .B(new_n235_), .C1(new_n230_), .C2(G204gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n233_), .A2(new_n234_), .A3(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT86), .ZN(new_n238_));
  OR3_X1    g037(.A1(new_n231_), .A2(new_n232_), .A3(new_n234_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n228_), .A2(new_n240_), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n241_), .A2(KEYINPUT91), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT20), .ZN(new_n243_));
  INV_X1    g042(.A(new_n240_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n226_), .A2(new_n223_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n207_), .B1(new_n211_), .B2(new_n208_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n216_), .A2(new_n246_), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n243_), .B1(new_n244_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n241_), .A2(KEYINPUT91), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n242_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G226gat), .A2(G233gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n252_), .B(KEYINPUT19), .Z(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT87), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n251_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT94), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n228_), .B(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(new_n244_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n248_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n243_), .B1(new_n240_), .B2(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n253_), .B1(new_n259_), .B2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n206_), .B1(new_n256_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n251_), .A2(new_n255_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n244_), .A2(new_n227_), .A3(new_n217_), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n265_), .A2(new_n253_), .A3(new_n261_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n264_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G141gat), .A2(G148gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT82), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT2), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(G141gat), .A2(G148gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT3), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n272_), .B(new_n274_), .C1(new_n271_), .C2(new_n269_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G155gat), .A2(G162gat), .ZN(new_n276_));
  INV_X1    g075(.A(G155gat), .ZN(new_n277_));
  INV_X1    g076(.A(G162gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n275_), .A2(new_n276_), .A3(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n276_), .A2(KEYINPUT1), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT83), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n279_), .B1(KEYINPUT1), .B2(new_n276_), .ZN(new_n283_));
  OAI221_X1 g082(.A(new_n270_), .B1(G141gat), .B2(G148gat), .C1(new_n282_), .C2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n280_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G127gat), .B(G134gat), .ZN(new_n286_));
  INV_X1    g085(.A(G113gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(G120gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n285_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(G120gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n288_), .B(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n292_), .B1(new_n280_), .B2(new_n284_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n290_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G225gat), .A2(G233gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT92), .B1(new_n294_), .B2(KEYINPUT4), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT4), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n298_), .B1(new_n299_), .B2(new_n293_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n294_), .A2(KEYINPUT92), .A3(KEYINPUT4), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n297_), .B1(new_n302_), .B2(new_n296_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT0), .B(G57gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(G85gat), .ZN(new_n305_));
  XOR2_X1   g104(.A(G1gat), .B(G29gat), .Z(new_n306_));
  XOR2_X1   g105(.A(new_n305_), .B(new_n306_), .Z(new_n307_));
  AND2_X1   g106(.A1(new_n303_), .A2(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n303_), .A2(new_n307_), .ZN(new_n309_));
  OAI221_X1 g108(.A(new_n263_), .B1(new_n268_), .B2(new_n206_), .C1(new_n308_), .C2(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n205_), .B1(new_n264_), .B2(new_n267_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n205_), .ZN(new_n312_));
  AOI211_X1 g111(.A(new_n312_), .B(new_n266_), .C1(new_n251_), .C2(new_n255_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n294_), .A2(new_n296_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n307_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n300_), .A2(new_n295_), .A3(new_n301_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT93), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n314_), .B1(new_n316_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n309_), .A2(KEYINPUT33), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT33), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n321_), .B1(new_n303_), .B2(new_n307_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n310_), .B1(new_n319_), .B2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n248_), .B(KEYINPUT30), .ZN(new_n325_));
  XOR2_X1   g124(.A(G15gat), .B(G43gat), .Z(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G227gat), .A2(G233gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT80), .ZN(new_n329_));
  XOR2_X1   g128(.A(G71gat), .B(G99gat), .Z(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n327_), .B(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT81), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n289_), .B(KEYINPUT31), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n332_), .A2(new_n333_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n334_), .A2(new_n337_), .A3(new_n335_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n285_), .A2(KEYINPUT29), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n240_), .A2(new_n340_), .ZN(new_n341_));
  XOR2_X1   g140(.A(G78gat), .B(G106gat), .Z(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G228gat), .A2(G233gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT84), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n285_), .A2(KEYINPUT29), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT28), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G22gat), .B(G50gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n346_), .B(new_n350_), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n324_), .A2(new_n339_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n339_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT95), .B(KEYINPUT27), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n355_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n312_), .B1(new_n256_), .B2(new_n262_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n264_), .A2(new_n205_), .A3(new_n267_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n357_), .A2(KEYINPUT27), .A3(new_n358_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n356_), .A2(new_n359_), .A3(KEYINPUT96), .ZN(new_n360_));
  AOI21_X1  g159(.A(KEYINPUT96), .B1(new_n356_), .B2(new_n359_), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n353_), .B(new_n351_), .C1(new_n360_), .C2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n351_), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n363_), .A2(new_n339_), .A3(new_n356_), .A4(new_n359_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n308_), .A2(new_n309_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n352_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT11), .ZN(new_n369_));
  AND2_X1   g168(.A1(G57gat), .A2(G64gat), .ZN(new_n370_));
  NOR2_X1   g169(.A1(G57gat), .A2(G64gat), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT66), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(G57gat), .ZN(new_n373_));
  INV_X1    g172(.A(G64gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT66), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G57gat), .A2(G64gat), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n369_), .B1(new_n372_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n372_), .A2(new_n378_), .A3(new_n369_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT67), .ZN(new_n382_));
  XOR2_X1   g181(.A(G71gat), .B(G78gat), .Z(new_n383_));
  AND3_X1   g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n382_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n380_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n381_), .A2(new_n383_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT67), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(new_n389_), .A3(new_n379_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n386_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G231gat), .A2(G233gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT14), .ZN(new_n394_));
  AND2_X1   g193(.A1(KEYINPUT74), .A2(G1gat), .ZN(new_n395_));
  NOR2_X1   g194(.A1(KEYINPUT74), .A2(G1gat), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n394_), .B1(new_n397_), .B2(G8gat), .ZN(new_n398_));
  XOR2_X1   g197(.A(G15gat), .B(G22gat), .Z(new_n399_));
  NOR3_X1   g198(.A1(new_n398_), .A2(KEYINPUT75), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT75), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT74), .B(G1gat), .ZN(new_n402_));
  INV_X1    g201(.A(G8gat), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT14), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n399_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n401_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(G1gat), .B1(new_n400_), .B2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT75), .B1(new_n398_), .B2(new_n399_), .ZN(new_n408_));
  INV_X1    g207(.A(G1gat), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n404_), .A2(new_n401_), .A3(new_n405_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n408_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n407_), .A2(G8gat), .A3(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(G8gat), .B1(new_n407_), .B2(new_n411_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n393_), .B(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT76), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT16), .B(G183gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(G211gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G127gat), .B(G155gat), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n419_), .B(new_n420_), .Z(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT17), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n417_), .B(new_n423_), .ZN(new_n424_));
  OR3_X1    g223(.A1(new_n416_), .A2(KEYINPUT17), .A3(new_n422_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G85gat), .B(G92gat), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G99gat), .A2(G106gat), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT6), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(KEYINPUT8), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT7), .ZN(new_n435_));
  INV_X1    g234(.A(G99gat), .ZN(new_n436_));
  INV_X1    g235(.A(G106gat), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n435_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n429_), .B1(new_n434_), .B2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n441_), .A2(KEYINPUT65), .A3(KEYINPUT8), .ZN(new_n442_));
  NAND2_X1  g241(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n429_), .B(new_n443_), .C1(new_n434_), .C2(new_n440_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT9), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(G85gat), .A3(G92gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT10), .B(G99gat), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n446_), .B1(new_n447_), .B2(G106gat), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n428_), .A2(new_n445_), .ZN(new_n449_));
  OAI22_X1  g248(.A1(new_n448_), .A2(new_n449_), .B1(KEYINPUT8), .B2(new_n440_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n432_), .A2(new_n433_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT64), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n442_), .A2(new_n444_), .B1(new_n450_), .B2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n454_), .A2(new_n386_), .A3(new_n390_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G230gat), .A2(G233gat), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n442_), .A2(new_n444_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n450_), .A2(new_n453_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NOR3_X1   g259(.A1(new_n384_), .A2(new_n385_), .A3(new_n380_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n379_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n460_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT12), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n391_), .A2(KEYINPUT12), .A3(new_n460_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n457_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n463_), .A2(new_n455_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n456_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(G120gat), .B(G148gat), .Z(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G176gat), .B(G204gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n474_), .B(new_n475_), .Z(new_n476_));
  XNOR2_X1  g275(.A(new_n471_), .B(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT13), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G229gat), .A2(G233gat), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NOR3_X1   g280(.A1(new_n400_), .A2(new_n406_), .A3(G1gat), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n409_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n403_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT69), .B(G29gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(G36gat), .ZN(new_n486_));
  XOR2_X1   g285(.A(G43gat), .B(G50gat), .Z(new_n487_));
  AND2_X1   g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n486_), .A2(new_n487_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  AND3_X1   g289(.A1(new_n484_), .A2(new_n490_), .A3(new_n412_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n490_), .B1(new_n484_), .B2(new_n412_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n481_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n486_), .B(new_n487_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n494_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n490_), .A2(KEYINPUT15), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT15), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n494_), .A2(new_n497_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n484_), .A2(new_n496_), .A3(new_n412_), .A4(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n495_), .A2(new_n499_), .A3(new_n480_), .ZN(new_n500_));
  XOR2_X1   g299(.A(G113gat), .B(G141gat), .Z(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(G169gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(new_n229_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n493_), .A2(new_n500_), .A3(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT78), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n505_), .A2(new_n506_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT77), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n493_), .A2(new_n500_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n509_), .B1(new_n510_), .B2(new_n503_), .ZN(new_n511_));
  AOI211_X1 g310(.A(KEYINPUT77), .B(new_n504_), .C1(new_n493_), .C2(new_n500_), .ZN(new_n512_));
  OAI22_X1  g311(.A1(new_n507_), .A2(new_n508_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NOR3_X1   g313(.A1(new_n427_), .A2(new_n479_), .A3(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT37), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n496_), .A2(new_n460_), .A3(new_n498_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n494_), .A2(new_n454_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G232gat), .A2(G233gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT34), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n517_), .B(new_n518_), .C1(KEYINPUT35), .C2(new_n520_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n520_), .A2(KEYINPUT35), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n522_), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n523_), .A2(KEYINPUT73), .A3(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT73), .B1(new_n523_), .B2(new_n524_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT70), .B(G134gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(G162gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G190gat), .B(G218gat), .ZN(new_n529_));
  XOR2_X1   g328(.A(new_n528_), .B(new_n529_), .Z(new_n530_));
  XOR2_X1   g329(.A(new_n530_), .B(KEYINPUT36), .Z(new_n531_));
  NOR3_X1   g330(.A1(new_n525_), .A2(new_n526_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n523_), .A2(new_n524_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT71), .B(KEYINPUT36), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n530_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT72), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n534_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n516_), .B1(new_n532_), .B2(new_n539_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n538_), .B(KEYINPUT37), .C1(new_n534_), .C2(new_n531_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n368_), .A2(new_n515_), .A3(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n366_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n545_), .A2(new_n546_), .A3(new_n402_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT38), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT97), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n367_), .B1(new_n549_), .B2(new_n515_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n532_), .A2(new_n539_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n550_), .B(new_n552_), .C1(new_n549_), .C2(new_n515_), .ZN(new_n553_));
  OAI21_X1  g352(.A(G1gat), .B1(new_n553_), .B2(new_n366_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n548_), .A2(new_n554_), .ZN(G1324gat));
  NOR2_X1   g354(.A1(new_n360_), .A2(new_n361_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n545_), .A2(new_n403_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n556_), .ZN(new_n558_));
  OAI21_X1  g357(.A(G8gat), .B1(new_n553_), .B2(new_n558_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n559_), .A2(KEYINPUT39), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(KEYINPUT39), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n557_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT40), .Z(G1325gat));
  NOR3_X1   g362(.A1(new_n544_), .A2(G15gat), .A3(new_n339_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT98), .ZN(new_n565_));
  OAI21_X1  g364(.A(G15gat), .B1(new_n553_), .B2(new_n339_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT41), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n566_), .A2(new_n567_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n565_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n570_), .B(KEYINPUT99), .Z(G1326gat));
  OAI21_X1  g370(.A(G22gat), .B1(new_n553_), .B2(new_n351_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT42), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n351_), .A2(G22gat), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n573_), .B1(new_n544_), .B2(new_n574_), .ZN(G1327gat));
  NOR2_X1   g374(.A1(new_n479_), .A2(new_n514_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(new_n427_), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n367_), .A2(new_n552_), .A3(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(G29gat), .B1(new_n578_), .B2(new_n546_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT44), .ZN(new_n580_));
  INV_X1    g379(.A(new_n577_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n581_), .A2(KEYINPUT101), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT43), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT100), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n583_), .B1(new_n542_), .B2(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n585_), .B1(new_n367_), .B2(new_n543_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n546_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n587_));
  OAI221_X1 g386(.A(new_n542_), .B1(new_n584_), .B2(new_n583_), .C1(new_n587_), .C2(new_n352_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n580_), .B(new_n582_), .C1(new_n589_), .C2(KEYINPUT101), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  AOI211_X1 g390(.A(KEYINPUT101), .B(new_n580_), .C1(new_n589_), .C2(new_n581_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n593_), .A2(new_n366_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n579_), .B1(new_n594_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g394(.A(G36gat), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT101), .B1(new_n589_), .B2(new_n581_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(KEYINPUT44), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(new_n590_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n596_), .B1(new_n599_), .B2(new_n556_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n578_), .A2(new_n596_), .A3(new_n556_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n602_), .A2(KEYINPUT102), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(KEYINPUT102), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n603_), .A2(KEYINPUT45), .A3(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(KEYINPUT45), .B1(new_n603_), .B2(new_n604_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT103), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT46), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n601_), .A2(new_n608_), .A3(new_n609_), .A4(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n609_), .A2(new_n610_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n607_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(new_n605_), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n612_), .B(new_n613_), .C1(new_n615_), .C2(new_n600_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n611_), .A2(new_n616_), .ZN(G1329gat));
  INV_X1    g416(.A(KEYINPUT47), .ZN(new_n618_));
  OAI211_X1 g417(.A(G43gat), .B(new_n353_), .C1(new_n591_), .C2(new_n592_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT104), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n578_), .A2(new_n353_), .ZN(new_n621_));
  INV_X1    g420(.A(G43gat), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n619_), .A2(new_n620_), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n620_), .B1(new_n619_), .B2(new_n623_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n618_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n626_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(KEYINPUT47), .A3(new_n624_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(G1330gat));
  OAI21_X1  g429(.A(G50gat), .B1(new_n593_), .B2(new_n351_), .ZN(new_n631_));
  INV_X1    g430(.A(G50gat), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n578_), .A2(new_n632_), .A3(new_n363_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT105), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(G1331gat));
  NOR2_X1   g435(.A1(new_n367_), .A2(new_n513_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(new_n552_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n479_), .A2(new_n426_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n641_), .A2(new_n373_), .A3(new_n366_), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n637_), .A2(KEYINPUT106), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n637_), .A2(KEYINPUT106), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n540_), .A2(new_n426_), .A3(new_n541_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n645_), .A2(new_n479_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(new_n546_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n642_), .B1(new_n650_), .B2(new_n373_), .ZN(G1332gat));
  AOI21_X1  g450(.A(new_n374_), .B1(new_n640_), .B2(new_n556_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT48), .Z(new_n653_));
  NAND2_X1  g452(.A1(new_n556_), .A2(new_n374_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n653_), .B1(new_n648_), .B2(new_n654_), .ZN(G1333gat));
  INV_X1    g454(.A(G71gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n649_), .A2(new_n656_), .A3(new_n353_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n656_), .B1(new_n640_), .B2(new_n353_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT107), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n659_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n660_), .A2(KEYINPUT49), .A3(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT49), .B1(new_n660_), .B2(new_n661_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n657_), .B1(new_n662_), .B2(new_n663_), .ZN(G1334gat));
  INV_X1    g463(.A(G78gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n649_), .A2(new_n665_), .A3(new_n363_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n640_), .B2(new_n363_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT108), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n668_), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n669_), .A2(KEYINPUT50), .A3(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(KEYINPUT50), .B1(new_n669_), .B2(new_n670_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n666_), .B1(new_n671_), .B2(new_n672_), .ZN(G1335gat));
  NOR2_X1   g472(.A1(new_n426_), .A2(new_n478_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n643_), .A2(new_n551_), .A3(new_n644_), .A4(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT109), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n675_), .B(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(G85gat), .B1(new_n677_), .B2(new_n546_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n674_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n679_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(new_n514_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n681_), .A2(new_n366_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n678_), .B1(G85gat), .B2(new_n682_), .ZN(G1336gat));
  INV_X1    g482(.A(G92gat), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n681_), .A2(new_n684_), .A3(new_n558_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n677_), .A2(new_n556_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n686_), .B2(new_n684_), .ZN(G1337gat));
  INV_X1    g486(.A(new_n447_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n675_), .A2(new_n676_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n675_), .A2(new_n676_), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n688_), .B(new_n353_), .C1(new_n689_), .C2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n680_), .A2(new_n514_), .A3(new_n353_), .ZN(new_n692_));
  AOI21_X1  g491(.A(KEYINPUT110), .B1(new_n692_), .B2(G99gat), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n692_), .A2(KEYINPUT110), .A3(G99gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n691_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT111), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n695_), .A2(new_n696_), .A3(KEYINPUT51), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(KEYINPUT51), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n691_), .B(new_n698_), .C1(new_n693_), .C2(new_n694_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(G1338gat));
  NAND3_X1  g499(.A1(new_n680_), .A2(new_n514_), .A3(new_n363_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT112), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT112), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n680_), .A2(new_n703_), .A3(new_n514_), .A4(new_n363_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n702_), .A2(G106gat), .A3(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT52), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT52), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n702_), .A2(new_n707_), .A3(G106gat), .A4(new_n704_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n677_), .A2(new_n437_), .A3(new_n363_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT53), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT53), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n709_), .A2(new_n710_), .A3(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(G1339gat));
  NAND2_X1  g514(.A1(new_n478_), .A2(new_n514_), .ZN(new_n716_));
  OR3_X1    g515(.A1(new_n646_), .A2(KEYINPUT113), .A3(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(KEYINPUT113), .B1(new_n646_), .B2(new_n716_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n717_), .A2(KEYINPUT54), .A3(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT54), .B1(new_n717_), .B2(new_n718_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n471_), .A2(new_n476_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n513_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT114), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n465_), .A2(new_n455_), .A3(new_n466_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n467_), .A2(KEYINPUT55), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT55), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n457_), .A2(new_n465_), .A3(new_n729_), .A4(new_n466_), .ZN(new_n730_));
  AOI221_X4 g529(.A(new_n726_), .B1(new_n469_), .B2(new_n727_), .C1(new_n728_), .C2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n728_), .A2(new_n730_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n727_), .A2(new_n469_), .ZN(new_n733_));
  AOI21_X1  g532(.A(KEYINPUT114), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n476_), .B1(new_n731_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT56), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  AOI221_X4 g536(.A(new_n464_), .B1(new_n458_), .B2(new_n459_), .C1(new_n386_), .C2(new_n390_), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT12), .B1(new_n391_), .B2(new_n460_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n729_), .B1(new_n740_), .B2(new_n457_), .ZN(new_n741_));
  AND4_X1   g540(.A1(new_n729_), .A2(new_n457_), .A3(new_n465_), .A4(new_n466_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n733_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(new_n726_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n732_), .A2(KEYINPUT114), .A3(new_n733_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n746_), .A2(KEYINPUT56), .A3(new_n476_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n725_), .B1(new_n737_), .B2(new_n747_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n491_), .A2(new_n492_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n749_), .A2(new_n481_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n495_), .A2(new_n499_), .A3(new_n481_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n750_), .A2(new_n751_), .A3(new_n504_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n508_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n505_), .A2(new_n506_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n752_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n477_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n552_), .B1(new_n748_), .B2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT57), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n513_), .A2(new_n724_), .ZN(new_n761_));
  AOI21_X1  g560(.A(KEYINPUT56), .B1(new_n746_), .B2(new_n476_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n476_), .ZN(new_n763_));
  AOI211_X1 g562(.A(new_n736_), .B(new_n763_), .C1(new_n744_), .C2(new_n745_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n761_), .B1(new_n762_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n756_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n766_), .A2(KEYINPUT57), .A3(new_n552_), .ZN(new_n767_));
  AOI211_X1 g566(.A(new_n723_), .B(new_n752_), .C1(new_n753_), .C2(new_n754_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n768_), .B1(new_n762_), .B2(new_n764_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT58), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  OAI211_X1 g570(.A(KEYINPUT58), .B(new_n768_), .C1(new_n762_), .C2(new_n764_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n542_), .A3(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n760_), .A2(new_n767_), .A3(new_n773_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT115), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n722_), .B1(new_n775_), .B2(new_n426_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n362_), .A2(new_n366_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(G113gat), .B1(new_n779_), .B2(new_n513_), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n771_), .A2(new_n542_), .A3(new_n772_), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT57), .B1(new_n766_), .B2(new_n552_), .ZN(new_n782_));
  OAI21_X1  g581(.A(KEYINPUT117), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT117), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n760_), .A2(new_n773_), .A3(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n783_), .A2(new_n767_), .A3(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT118), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n786_), .A2(new_n787_), .A3(new_n427_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n786_), .B2(new_n427_), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n721_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n777_), .B(KEYINPUT116), .ZN(new_n791_));
  OR3_X1    g590(.A1(new_n790_), .A2(KEYINPUT59), .A3(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n778_), .A2(KEYINPUT59), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n794_), .A2(new_n514_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n780_), .B1(new_n795_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g595(.A(new_n291_), .B1(new_n478_), .B2(KEYINPUT60), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n779_), .B(new_n797_), .C1(KEYINPUT60), .C2(new_n291_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n794_), .A2(new_n478_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(new_n291_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT119), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(KEYINPUT119), .B(new_n798_), .C1(new_n799_), .C2(new_n291_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(G1341gat));
  AOI21_X1  g603(.A(G127gat), .B1(new_n779_), .B2(new_n426_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n794_), .A2(new_n427_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g606(.A(G134gat), .B1(new_n779_), .B2(new_n551_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n794_), .A2(new_n543_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n809_), .B2(G134gat), .ZN(G1343gat));
  AND3_X1   g609(.A1(new_n776_), .A2(new_n339_), .A3(new_n363_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n811_), .A2(new_n546_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n558_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(new_n514_), .ZN(new_n814_));
  XOR2_X1   g613(.A(new_n814_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g614(.A1(new_n813_), .A2(new_n478_), .ZN(new_n816_));
  XOR2_X1   g615(.A(new_n816_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g616(.A1(new_n813_), .A2(new_n427_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(new_n277_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n818_), .B(new_n820_), .ZN(G1346gat));
  NOR3_X1   g620(.A1(new_n813_), .A2(new_n278_), .A3(new_n543_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n812_), .A2(new_n558_), .A3(new_n551_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n278_), .B2(new_n823_), .ZN(G1347gat));
  AND3_X1   g623(.A1(new_n760_), .A2(new_n784_), .A3(new_n773_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n784_), .B1(new_n760_), .B2(new_n773_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n767_), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n825_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT118), .B1(new_n828_), .B2(new_n426_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n786_), .A2(new_n787_), .A3(new_n427_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n722_), .A3(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n558_), .A2(new_n546_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n353_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n833_), .A2(new_n363_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n831_), .A2(new_n834_), .ZN(new_n835_));
  OR3_X1    g634(.A1(new_n835_), .A2(KEYINPUT121), .A3(new_n514_), .ZN(new_n836_));
  OAI21_X1  g635(.A(KEYINPUT121), .B1(new_n835_), .B2(new_n514_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(G169gat), .A3(new_n837_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(KEYINPUT62), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT122), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n831_), .A2(new_n840_), .A3(new_n834_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n840_), .B1(new_n831_), .B2(new_n834_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n513_), .A2(new_n210_), .ZN(new_n844_));
  XOR2_X1   g643(.A(new_n844_), .B(KEYINPUT123), .Z(new_n845_));
  OAI21_X1  g644(.A(new_n839_), .B1(new_n843_), .B2(new_n845_), .ZN(G1348gat));
  AND2_X1   g645(.A1(new_n776_), .A2(new_n351_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n833_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n847_), .A2(G176gat), .A3(new_n479_), .A4(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n834_), .ZN(new_n850_));
  OAI21_X1  g649(.A(KEYINPUT122), .B1(new_n790_), .B2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n831_), .A2(new_n840_), .A3(new_n834_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n478_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n211_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n853_), .A2(KEYINPUT124), .A3(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT124), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n479_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(new_n211_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n849_), .B1(new_n855_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT125), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  OAI211_X1 g660(.A(KEYINPUT125), .B(new_n849_), .C1(new_n855_), .C2(new_n858_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1349gat));
  NOR3_X1   g662(.A1(new_n843_), .A2(new_n427_), .A3(new_n221_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n833_), .A2(new_n427_), .ZN(new_n865_));
  AOI21_X1  g664(.A(G183gat), .B1(new_n847_), .B2(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n864_), .A2(new_n866_), .ZN(G1350gat));
  OAI21_X1  g666(.A(G190gat), .B1(new_n843_), .B2(new_n543_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n551_), .A2(new_n222_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n843_), .B2(new_n869_), .ZN(G1351gat));
  NAND2_X1  g669(.A1(new_n811_), .A2(new_n832_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n513_), .ZN(new_n873_));
  OR2_X1    g672(.A1(new_n229_), .A2(KEYINPUT126), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n229_), .A2(KEYINPUT126), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n873_), .A2(new_n874_), .A3(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n873_), .B2(new_n875_), .ZN(G1352gat));
  NAND2_X1  g676(.A1(new_n872_), .A2(new_n479_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g678(.A1(new_n872_), .A2(new_n426_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n881_));
  AND2_X1   g680(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n880_), .A2(new_n881_), .A3(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n883_), .B1(new_n880_), .B2(new_n881_), .ZN(G1354gat));
  AOI21_X1  g683(.A(G218gat), .B1(new_n872_), .B2(new_n551_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n542_), .A2(G218gat), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(KEYINPUT127), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n885_), .B1(new_n872_), .B2(new_n887_), .ZN(G1355gat));
endmodule


