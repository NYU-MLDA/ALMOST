//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n785_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n893_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n944_, new_n945_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n954_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n965_, new_n966_;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G113gat), .B(G120gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT91), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT31), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n206_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n207_), .A2(KEYINPUT90), .A3(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G227gat), .A2(G233gat), .ZN(new_n210_));
  INV_X1    g009(.A(G15gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT30), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n209_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n213_), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n207_), .A2(KEYINPUT90), .A3(new_n208_), .A4(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(G169gat), .ZN(new_n219_));
  OR2_X1    g018(.A1(KEYINPUT87), .A2(G190gat), .ZN(new_n220_));
  INV_X1    g019(.A(G183gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(KEYINPUT87), .A2(G190gat), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n219_), .B1(new_n223_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT24), .ZN(new_n228_));
  OR3_X1    g027(.A1(KEYINPUT89), .A2(G169gat), .A3(G176gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT89), .B1(G169gat), .B2(G176gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n226_), .B1(new_n228_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n231_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n228_), .B1(G169gat), .B2(G176gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n232_), .A2(new_n235_), .ZN(new_n236_));
  OR3_X1    g035(.A1(new_n221_), .A2(KEYINPUT86), .A3(KEYINPUT25), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT25), .B1(new_n221_), .B2(KEYINPUT86), .ZN(new_n238_));
  INV_X1    g037(.A(G190gat), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n237_), .B(new_n238_), .C1(KEYINPUT26), .C2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n220_), .A2(KEYINPUT26), .A3(new_n222_), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n241_), .A2(KEYINPUT88), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(KEYINPUT88), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n240_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n227_), .B1(new_n236_), .B2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G71gat), .B(G99gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(G43gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n245_), .B(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n217_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n214_), .A2(new_n248_), .A3(new_n216_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT2), .ZN(new_n254_));
  INV_X1    g053(.A(G141gat), .ZN(new_n255_));
  INV_X1    g054(.A(G148gat), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n254_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT3), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n257_), .A2(new_n259_), .A3(new_n260_), .A4(new_n261_), .ZN(new_n262_));
  OR2_X1    g061(.A1(G155gat), .A2(G162gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G155gat), .A2(G162gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT92), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n263_), .A2(KEYINPUT92), .A3(new_n264_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n262_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  XOR2_X1   g068(.A(G141gat), .B(G148gat), .Z(new_n270_));
  NAND2_X1  g069(.A1(new_n264_), .A2(KEYINPUT1), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n263_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n264_), .A2(KEYINPUT1), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n270_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n269_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT93), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT93), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n269_), .A2(new_n274_), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT29), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT28), .ZN(new_n282_));
  XOR2_X1   g081(.A(G22gat), .B(G50gat), .Z(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(G78gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G228gat), .A2(G233gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT95), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n280_), .B1(new_n269_), .B2(new_n274_), .ZN(new_n289_));
  INV_X1    g088(.A(G197gat), .ZN(new_n290_));
  INV_X1    g089(.A(G204gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G197gat), .A2(G204gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT21), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n292_), .A2(KEYINPUT21), .A3(new_n293_), .ZN(new_n297_));
  INV_X1    g096(.A(G211gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT96), .B1(new_n298_), .B2(G218gat), .ZN(new_n299_));
  INV_X1    g098(.A(G218gat), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n300_), .A2(G211gat), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n296_), .A2(new_n297_), .A3(new_n302_), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n292_), .A2(new_n293_), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n304_), .B(KEYINPUT21), .C1(new_n301_), .C2(new_n299_), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n288_), .B1(new_n289_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT97), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT97), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n309_), .B(new_n288_), .C1(new_n289_), .C2(new_n306_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT98), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n306_), .A2(new_n288_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n313_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n311_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n312_), .B1(new_n311_), .B2(new_n314_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n286_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n303_), .A2(new_n305_), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n269_), .A2(new_n274_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n318_), .B1(new_n319_), .B2(new_n280_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n309_), .B1(new_n320_), .B2(new_n288_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n310_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n314_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT98), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n311_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(G78gat), .A3(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n317_), .A2(new_n326_), .A3(G106gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT94), .ZN(new_n328_));
  AOI21_X1  g127(.A(G106gat), .B1(new_n317_), .B2(new_n326_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n285_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n329_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n331_), .A2(KEYINPUT94), .A3(new_n327_), .A4(new_n284_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G226gat), .A2(G233gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT19), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT20), .B1(new_n245_), .B2(new_n318_), .ZN(new_n336_));
  OR2_X1    g135(.A1(new_n234_), .A2(KEYINPUT100), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n234_), .A2(KEYINPUT100), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n233_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(KEYINPUT25), .B(G183gat), .Z(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT99), .ZN(new_n341_));
  XOR2_X1   g140(.A(KEYINPUT26), .B(G190gat), .Z(new_n342_));
  OAI211_X1 g141(.A(new_n339_), .B(new_n232_), .C1(new_n341_), .C2(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(G183gat), .A2(G190gat), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n219_), .B1(new_n226_), .B2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n306_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n335_), .B1(new_n336_), .B2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G8gat), .B(G36gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT18), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G64gat), .B(G92gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n352_), .A2(KEYINPUT32), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n245_), .A2(new_n318_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n343_), .A2(new_n306_), .A3(new_n345_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n335_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n355_), .A2(new_n356_), .A3(KEYINPUT20), .A4(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n347_), .A2(new_n354_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT103), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NOR3_X1   g160(.A1(new_n336_), .A2(new_n335_), .A3(new_n346_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n355_), .A2(KEYINPUT20), .A3(new_n356_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n362_), .B1(new_n335_), .B2(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT103), .B1(new_n364_), .B2(new_n354_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n361_), .B1(new_n365_), .B2(new_n359_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n204_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n276_), .A2(new_n278_), .A3(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n368_), .B1(new_n370_), .B2(KEYINPUT4), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n319_), .A2(new_n204_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(KEYINPUT4), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT101), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n370_), .A2(KEYINPUT101), .A3(KEYINPUT4), .A4(new_n372_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n371_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT102), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n370_), .A2(new_n372_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n380_), .A2(new_n368_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n381_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G1gat), .B(G29gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(G85gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT0), .B(G57gat), .ZN(new_n385_));
  XOR2_X1   g184(.A(new_n384_), .B(new_n385_), .Z(new_n386_));
  NAND3_X1  g185(.A1(new_n379_), .A2(new_n382_), .A3(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n386_), .B1(new_n379_), .B2(new_n382_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n366_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT33), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n387_), .A2(new_n391_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n379_), .A2(new_n382_), .A3(KEYINPUT33), .A4(new_n386_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n347_), .A2(new_n358_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n351_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n347_), .A2(new_n352_), .A3(new_n358_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n386_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n398_), .B1(new_n380_), .B2(new_n367_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n375_), .A2(new_n376_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n370_), .A2(KEYINPUT4), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n401_), .A2(new_n368_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n399_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n397_), .A2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n392_), .A2(new_n393_), .A3(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n333_), .B1(new_n390_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n379_), .A2(new_n382_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n398_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n387_), .ZN(new_n409_));
  OAI211_X1 g208(.A(KEYINPUT27), .B(new_n396_), .C1(new_n364_), .C2(new_n352_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT27), .ZN(new_n411_));
  AOI21_X1  g210(.A(KEYINPUT104), .B1(new_n397_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT104), .ZN(new_n413_));
  AOI211_X1 g212(.A(new_n413_), .B(KEYINPUT27), .C1(new_n395_), .C2(new_n396_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n410_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n415_));
  AOI211_X1 g214(.A(new_n409_), .B(new_n415_), .C1(new_n332_), .C2(new_n330_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n253_), .B1(new_n406_), .B2(new_n416_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n330_), .A2(new_n332_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT105), .ZN(new_n419_));
  INV_X1    g218(.A(new_n410_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n412_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n414_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n420_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n408_), .A2(new_n387_), .A3(new_n252_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n418_), .A2(new_n419_), .A3(new_n423_), .A4(new_n424_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n423_), .A2(new_n424_), .A3(new_n332_), .A4(new_n330_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT105), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n417_), .A2(new_n428_), .ZN(new_n429_));
  XOR2_X1   g228(.A(G1gat), .B(G8gat), .Z(new_n430_));
  INV_X1    g229(.A(KEYINPUT14), .ZN(new_n431_));
  XNOR2_X1  g230(.A(KEYINPUT77), .B(G1gat), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  XOR2_X1   g232(.A(KEYINPUT78), .B(G8gat), .Z(new_n434_));
  AOI21_X1  g233(.A(new_n431_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(G15gat), .B(G22gat), .Z(new_n436_));
  OAI21_X1  g235(.A(new_n430_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT79), .B(KEYINPUT80), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT78), .B(G8gat), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT14), .B1(new_n432_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n430_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n436_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n437_), .A2(new_n438_), .A3(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n438_), .B1(new_n437_), .B2(new_n443_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  XOR2_X1   g245(.A(G29gat), .B(G36gat), .Z(new_n447_));
  XOR2_X1   g246(.A(G43gat), .B(G50gat), .Z(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT15), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n446_), .A2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n449_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G229gat), .A2(G233gat), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n451_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT84), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n437_), .A2(new_n443_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n438_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n449_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n437_), .A2(new_n438_), .A3(new_n443_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n452_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n453_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n455_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  AOI211_X1 g263(.A(KEYINPUT84), .B(new_n453_), .C1(new_n452_), .C2(new_n461_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n454_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G113gat), .B(G141gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G169gat), .B(G197gat), .ZN(new_n468_));
  XOR2_X1   g267(.A(new_n467_), .B(new_n468_), .Z(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n466_), .A2(new_n470_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n454_), .B(new_n469_), .C1(new_n464_), .C2(new_n465_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(KEYINPUT85), .A3(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT85), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n466_), .A2(new_n474_), .A3(new_n470_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G57gat), .B(G64gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT11), .ZN(new_n479_));
  XOR2_X1   g278(.A(G71gat), .B(G78gat), .Z(new_n480_));
  OR2_X1    g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n478_), .A2(KEYINPUT11), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n479_), .A2(new_n480_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n481_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G231gat), .A2(G233gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n458_), .A2(new_n460_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT82), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n446_), .A2(new_n486_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(G127gat), .B(G155gat), .Z(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G183gat), .B(G211gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT17), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n492_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n498_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .A4(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n489_), .A2(new_n491_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n497_), .A2(KEYINPUT17), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT83), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT83), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n502_), .A2(new_n508_), .A3(new_n505_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT64), .B(G92gat), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT9), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n512_), .A3(G85gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G85gat), .B(G92gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT10), .B(G99gat), .ZN(new_n515_));
  OAI221_X1 g314(.A(new_n513_), .B1(new_n512_), .B2(new_n514_), .C1(G106gat), .C2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT6), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT65), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT65), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT6), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G99gat), .A2(G106gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  AND2_X1   g322(.A1(G99gat), .A2(G106gat), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n518_), .A2(new_n520_), .A3(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n516_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT69), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n528_), .A2(KEYINPUT6), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n517_), .A2(KEYINPUT69), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n522_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(G99gat), .ZN(new_n532_));
  INV_X1    g331(.A(G106gat), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(new_n533_), .A3(KEYINPUT66), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT7), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT7), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n536_), .A2(new_n532_), .A3(new_n533_), .A4(KEYINPUT66), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n517_), .A2(KEYINPUT69), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n528_), .A2(KEYINPUT6), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n538_), .A2(new_n539_), .A3(new_n524_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n531_), .A2(new_n535_), .A3(new_n537_), .A4(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n514_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT70), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT70), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n541_), .A2(new_n545_), .A3(new_n542_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n544_), .A2(KEYINPUT8), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT8), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n548_), .A2(KEYINPUT68), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(KEYINPUT68), .ZN(new_n550_));
  NOR3_X1   g349(.A1(new_n514_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n535_), .A2(new_n537_), .ZN(new_n552_));
  NOR3_X1   g351(.A1(new_n526_), .A2(KEYINPUT67), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT67), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n518_), .A2(new_n520_), .A3(new_n524_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n524_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n535_), .A2(new_n537_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n554_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n551_), .B1(new_n553_), .B2(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n527_), .B1(new_n547_), .B2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n449_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G232gat), .A2(G233gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n565_), .A2(KEYINPUT35), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n562_), .A2(new_n566_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n538_), .A2(new_n539_), .A3(new_n524_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n524_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n514_), .B1(new_n570_), .B2(new_n558_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n548_), .B1(new_n571_), .B2(new_n545_), .ZN(new_n572_));
  OAI21_X1  g371(.A(KEYINPUT67), .B1(new_n526_), .B2(new_n552_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n557_), .A2(new_n558_), .A3(new_n554_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  AOI22_X1  g374(.A1(new_n572_), .A2(new_n544_), .B1(new_n575_), .B2(new_n551_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n450_), .B1(new_n576_), .B2(new_n527_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT76), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n565_), .A2(KEYINPUT35), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n579_), .B(KEYINPUT75), .Z(new_n580_));
  OAI211_X1 g379(.A(new_n567_), .B(new_n577_), .C1(new_n578_), .C2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n577_), .A2(new_n562_), .A3(new_n566_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n580_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n562_), .A2(new_n566_), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n582_), .B(new_n583_), .C1(KEYINPUT76), .C2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G190gat), .B(G218gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G134gat), .B(G162gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n588_), .A2(KEYINPUT36), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n581_), .A2(new_n585_), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n588_), .B(KEYINPUT36), .Z(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n593_), .B1(new_n581_), .B2(new_n585_), .ZN(new_n594_));
  OAI21_X1  g393(.A(KEYINPUT37), .B1(new_n591_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT37), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n581_), .A2(new_n585_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n596_), .B(new_n590_), .C1(new_n597_), .C2(new_n593_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n510_), .B1(new_n595_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(G230gat), .A2(G233gat), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n547_), .A2(new_n560_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n527_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n602_), .A2(new_n484_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT71), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n561_), .A2(KEYINPUT71), .A3(new_n484_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n561_), .A2(new_n484_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n601_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(KEYINPUT72), .B(KEYINPUT12), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n611_), .B1(new_n561_), .B2(new_n484_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n601_), .B1(new_n561_), .B2(new_n484_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n484_), .ZN(new_n614_));
  OAI211_X1 g413(.A(KEYINPUT12), .B(new_n614_), .C1(new_n576_), .C2(new_n527_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n612_), .A2(new_n613_), .A3(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT73), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT73), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n612_), .A2(new_n613_), .A3(new_n615_), .A4(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n610_), .A2(new_n617_), .A3(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G120gat), .B(G148gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT5), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G176gat), .B(G204gat), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n622_), .B(new_n623_), .Z(new_n624_));
  NAND2_X1  g423(.A1(new_n620_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n624_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n610_), .A2(new_n617_), .A3(new_n619_), .A4(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT13), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n625_), .A2(KEYINPUT13), .A3(new_n627_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n600_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n429_), .A2(new_n477_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT106), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT106), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n429_), .A2(new_n636_), .A3(new_n477_), .A4(new_n633_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n409_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n638_), .A2(new_n433_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n635_), .A2(new_n637_), .A3(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(KEYINPUT107), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT107), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n635_), .A2(new_n642_), .A3(new_n637_), .A4(new_n639_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT38), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT109), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n644_), .A2(KEYINPUT109), .A3(new_n645_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n641_), .A2(KEYINPUT38), .A3(new_n643_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n405_), .A2(new_n390_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n418_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n333_), .A2(new_n638_), .A3(new_n423_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  AOI22_X1  g453(.A1(new_n654_), .A2(new_n253_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n591_), .A2(new_n594_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT108), .Z(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n655_), .A2(new_n510_), .A3(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n632_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(new_n477_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n659_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(new_n409_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(G1gat), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n648_), .A2(new_n649_), .A3(new_n650_), .A4(new_n665_), .ZN(G1324gat));
  NAND3_X1  g465(.A1(new_n659_), .A2(new_n415_), .A3(new_n662_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT39), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n667_), .A2(new_n668_), .A3(G8gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n667_), .B2(G8gat), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n635_), .A2(new_n637_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n415_), .A2(new_n439_), .ZN(new_n672_));
  OAI22_X1  g471(.A1(new_n669_), .A2(new_n670_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT40), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(G1325gat));
  NAND3_X1  g474(.A1(new_n659_), .A2(new_n252_), .A3(new_n662_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n676_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT41), .B1(new_n676_), .B2(G15gat), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n252_), .A2(new_n211_), .ZN(new_n679_));
  OAI22_X1  g478(.A1(new_n677_), .A2(new_n678_), .B1(new_n634_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT110), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(G1326gat));
  OR3_X1    g481(.A1(new_n634_), .A2(G22gat), .A3(new_n418_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n663_), .A2(new_n333_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(G22gat), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n685_), .A2(KEYINPUT42), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(KEYINPUT42), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n683_), .B1(new_n686_), .B2(new_n687_), .ZN(G1327gat));
  INV_X1    g487(.A(KEYINPUT111), .ZN(new_n689_));
  INV_X1    g488(.A(new_n510_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n661_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n595_), .A2(new_n598_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n692_), .B1(new_n429_), .B2(new_n694_), .ZN(new_n695_));
  AOI211_X1 g494(.A(KEYINPUT43), .B(new_n693_), .C1(new_n417_), .C2(new_n428_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n691_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(KEYINPUT43), .B1(new_n655_), .B2(new_n693_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n425_), .A2(new_n427_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n252_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n692_), .B(new_n694_), .C1(new_n701_), .C2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n700_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n704_), .A2(KEYINPUT44), .A3(new_n691_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n699_), .A2(new_n409_), .A3(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(G29gat), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n655_), .A2(new_n476_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n656_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n632_), .A2(new_n690_), .A3(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n711_), .A2(G29gat), .A3(new_n638_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n689_), .B1(new_n707_), .B2(new_n713_), .ZN(new_n714_));
  AOI211_X1 g513(.A(KEYINPUT111), .B(new_n712_), .C1(new_n706_), .C2(G29gat), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1328gat));
  XNOR2_X1  g515(.A(KEYINPUT112), .B(KEYINPUT46), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(G36gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT44), .B1(new_n704_), .B2(new_n691_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n691_), .ZN(new_n721_));
  AOI211_X1 g520(.A(new_n698_), .B(new_n721_), .C1(new_n700_), .C2(new_n703_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n719_), .B1(new_n723_), .B2(new_n415_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n423_), .A2(G36gat), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  OR3_X1    g525(.A1(new_n711_), .A2(KEYINPUT45), .A3(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(KEYINPUT45), .B1(new_n711_), .B2(new_n726_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n718_), .B1(new_n724_), .B2(new_n730_), .ZN(new_n731_));
  NOR3_X1   g530(.A1(new_n720_), .A2(new_n722_), .A3(new_n423_), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n729_), .B(new_n717_), .C1(new_n732_), .C2(new_n719_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1329gat));
  AND2_X1   g533(.A1(new_n252_), .A2(G43gat), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n699_), .A2(new_n705_), .A3(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n711_), .ZN(new_n737_));
  AOI21_X1  g536(.A(G43gat), .B1(new_n737_), .B2(new_n252_), .ZN(new_n738_));
  OR3_X1    g537(.A1(new_n736_), .A2(KEYINPUT47), .A3(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(KEYINPUT47), .B1(new_n736_), .B2(new_n738_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1330gat));
  AOI21_X1  g540(.A(G50gat), .B1(new_n737_), .B2(new_n333_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n333_), .A2(G50gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n723_), .B2(new_n743_), .ZN(G1331gat));
  NAND2_X1  g543(.A1(new_n632_), .A2(new_n476_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n659_), .A2(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G57gat), .B1(new_n747_), .B2(new_n638_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n655_), .A2(new_n477_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n660_), .A2(new_n600_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n638_), .A2(G57gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(G1332gat));
  OR3_X1    g552(.A1(new_n751_), .A2(G64gat), .A3(new_n423_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n747_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n415_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT48), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n756_), .A2(new_n757_), .A3(G64gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n756_), .B2(G64gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n754_), .B1(new_n758_), .B2(new_n759_), .ZN(G1333gat));
  INV_X1    g559(.A(new_n751_), .ZN(new_n761_));
  INV_X1    g560(.A(G71gat), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(new_n762_), .A3(new_n252_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT49), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n755_), .A2(new_n252_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(G71gat), .ZN(new_n766_));
  AOI211_X1 g565(.A(KEYINPUT49), .B(new_n762_), .C1(new_n755_), .C2(new_n252_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n763_), .B1(new_n766_), .B2(new_n767_), .ZN(G1334gat));
  NAND3_X1  g567(.A1(new_n761_), .A2(new_n286_), .A3(new_n333_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n755_), .A2(new_n333_), .ZN(new_n770_));
  XOR2_X1   g569(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n771_));
  AND3_X1   g570(.A1(new_n770_), .A2(G78gat), .A3(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n770_), .B2(G78gat), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(G1335gat));
  NAND2_X1  g573(.A1(new_n746_), .A2(new_n510_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n775_), .B1(new_n700_), .B2(new_n703_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(G85gat), .B1(new_n777_), .B2(new_n638_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n660_), .A2(new_n690_), .A3(new_n709_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n749_), .A2(new_n779_), .ZN(new_n780_));
  OR3_X1    g579(.A1(new_n780_), .A2(G85gat), .A3(new_n638_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n778_), .A2(new_n781_), .ZN(G1336gat));
  NAND3_X1  g581(.A1(new_n776_), .A2(new_n415_), .A3(new_n511_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n780_), .A2(new_n423_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n783_), .B1(G92gat), .B2(new_n784_), .ZN(new_n785_));
  XOR2_X1   g584(.A(new_n785_), .B(KEYINPUT114), .Z(G1337gat));
  NOR2_X1   g585(.A1(new_n777_), .A2(new_n253_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n787_), .A2(new_n532_), .ZN(new_n788_));
  OR2_X1    g587(.A1(new_n253_), .A2(new_n515_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n780_), .A2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(KEYINPUT51), .B1(new_n788_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792_));
  OAI221_X1 g591(.A(new_n792_), .B1(new_n780_), .B2(new_n789_), .C1(new_n787_), .C2(new_n532_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(G1338gat));
  NAND4_X1  g593(.A1(new_n749_), .A2(new_n533_), .A3(new_n333_), .A4(new_n779_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n776_), .A2(new_n333_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(G106gat), .ZN(new_n798_));
  AOI211_X1 g597(.A(KEYINPUT52), .B(new_n533_), .C1(new_n776_), .C2(new_n333_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n795_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT53), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n802_), .B(new_n795_), .C1(new_n798_), .C2(new_n799_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n803_), .ZN(G1339gat));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n473_), .A2(new_n475_), .A3(new_n627_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n612_), .A2(new_n613_), .A3(new_n615_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n606_), .A2(new_n612_), .A3(new_n607_), .A4(new_n615_), .ZN(new_n808_));
  AOI22_X1  g607(.A1(KEYINPUT55), .A2(new_n807_), .B1(new_n808_), .B2(new_n601_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n617_), .A2(new_n810_), .A3(new_n619_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n626_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n812_), .A2(KEYINPUT56), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT56), .ZN(new_n814_));
  AOI211_X1 g613(.A(new_n814_), .B(new_n626_), .C1(new_n809_), .C2(new_n811_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n806_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n462_), .A2(new_n453_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n451_), .A2(new_n452_), .A3(new_n463_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n470_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n472_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n472_), .A2(KEYINPUT117), .A3(new_n819_), .ZN(new_n823_));
  AOI22_X1  g622(.A1(new_n625_), .A2(new_n627_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n656_), .B1(new_n816_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n805_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  AND3_X1   g627(.A1(new_n617_), .A2(new_n810_), .A3(new_n619_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n808_), .A2(new_n601_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n612_), .A2(new_n613_), .A3(new_n615_), .A4(KEYINPUT55), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n624_), .B1(new_n829_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n814_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n812_), .A2(KEYINPUT56), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n824_), .B1(new_n836_), .B2(new_n806_), .ZN(new_n837_));
  OAI211_X1 g636(.A(KEYINPUT118), .B(KEYINPUT57), .C1(new_n837_), .C2(new_n656_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n828_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n627_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n840_), .B1(new_n823_), .B2(new_n822_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT58), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT58), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n841_), .B(new_n844_), .C1(new_n813_), .C2(new_n815_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n694_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n690_), .B1(new_n839_), .B2(new_n847_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n599_), .A2(new_n476_), .A3(new_n631_), .A4(new_n630_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT54), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT116), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n849_), .A2(new_n852_), .A3(KEYINPUT54), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n633_), .A2(KEYINPUT115), .A3(new_n854_), .A4(new_n476_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n856_), .B1(new_n849_), .B2(KEYINPUT54), .ZN(new_n857_));
  AOI22_X1  g656(.A1(new_n851_), .A2(new_n853_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n848_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n333_), .A2(new_n415_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n861_), .A2(new_n409_), .A3(new_n252_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n859_), .A2(new_n860_), .A3(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n847_), .A2(KEYINPUT119), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n846_), .A2(new_n866_), .A3(new_n694_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n865_), .A2(new_n839_), .A3(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n858_), .B1(new_n868_), .B2(new_n510_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n862_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n864_), .B1(new_n870_), .B2(new_n860_), .ZN(new_n871_));
  OAI21_X1  g670(.A(G113gat), .B1(new_n871_), .B2(new_n476_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n870_), .ZN(new_n873_));
  OR3_X1    g672(.A1(new_n873_), .A2(G113gat), .A3(new_n476_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n874_), .ZN(G1340gat));
  OAI21_X1  g674(.A(G120gat), .B1(new_n871_), .B2(new_n660_), .ZN(new_n876_));
  INV_X1    g675(.A(G120gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(new_n660_), .B2(KEYINPUT60), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n870_), .B(new_n878_), .C1(KEYINPUT60), .C2(new_n877_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n876_), .A2(new_n879_), .ZN(G1341gat));
  OAI21_X1  g679(.A(G127gat), .B1(new_n871_), .B2(new_n510_), .ZN(new_n881_));
  OR3_X1    g680(.A1(new_n873_), .A2(G127gat), .A3(new_n510_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(G1342gat));
  OAI21_X1  g682(.A(G134gat), .B1(new_n871_), .B2(new_n693_), .ZN(new_n884_));
  OR3_X1    g683(.A1(new_n873_), .A2(G134gat), .A3(new_n657_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1343gat));
  INV_X1    g685(.A(new_n869_), .ZN(new_n887_));
  NAND4_X1  g686(.A1(new_n333_), .A2(new_n409_), .A3(new_n423_), .A4(new_n253_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(KEYINPUT120), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n476_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(new_n255_), .ZN(G1344gat));
  NOR2_X1   g691(.A1(new_n890_), .A2(new_n660_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(new_n256_), .ZN(G1345gat));
  XOR2_X1   g693(.A(KEYINPUT61), .B(G155gat), .Z(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n887_), .A2(new_n690_), .A3(new_n889_), .A4(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n866_), .B1(new_n846_), .B2(new_n694_), .ZN(new_n898_));
  AOI211_X1 g697(.A(KEYINPUT119), .B(new_n693_), .C1(new_n843_), .C2(new_n845_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n690_), .B1(new_n900_), .B2(new_n839_), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n690_), .B(new_n889_), .C1(new_n901_), .C2(new_n858_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n895_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT121), .B(KEYINPUT122), .ZN(new_n904_));
  AND3_X1   g703(.A1(new_n897_), .A2(new_n903_), .A3(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n904_), .B1(new_n897_), .B2(new_n903_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1346gat));
  OAI21_X1  g706(.A(G162gat), .B1(new_n890_), .B2(new_n693_), .ZN(new_n908_));
  OR2_X1    g707(.A1(new_n657_), .A2(G162gat), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n890_), .B2(new_n909_), .ZN(G1347gat));
  NAND2_X1  g709(.A1(new_n424_), .A2(new_n415_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(new_n333_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n859_), .A2(new_n477_), .A3(new_n912_), .ZN(new_n913_));
  OAI21_X1  g712(.A(KEYINPUT62), .B1(new_n913_), .B2(KEYINPUT22), .ZN(new_n914_));
  OAI21_X1  g713(.A(G169gat), .B1(new_n913_), .B2(KEYINPUT62), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(G169gat), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(new_n914_), .ZN(G1348gat));
  NOR2_X1   g717(.A1(new_n869_), .A2(new_n333_), .ZN(new_n919_));
  INV_X1    g718(.A(G176gat), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n660_), .A2(new_n920_), .A3(new_n911_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n919_), .A2(new_n921_), .ZN(new_n922_));
  OAI211_X1 g721(.A(new_n632_), .B(new_n912_), .C1(new_n848_), .C2(new_n858_), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT123), .ZN(new_n924_));
  AND3_X1   g723(.A1(new_n923_), .A2(new_n924_), .A3(new_n920_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n924_), .B1(new_n923_), .B2(new_n920_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n922_), .B1(new_n925_), .B2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(KEYINPUT124), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n929_));
  OAI211_X1 g728(.A(new_n922_), .B(new_n929_), .C1(new_n925_), .C2(new_n926_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n928_), .A2(new_n930_), .ZN(G1349gat));
  NOR2_X1   g730(.A1(new_n911_), .A2(new_n510_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n919_), .A2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(new_n221_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n859_), .A2(new_n912_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n690_), .A2(new_n341_), .ZN(new_n936_));
  OR2_X1    g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n934_), .A2(new_n937_), .A3(KEYINPUT125), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT125), .ZN(new_n939_));
  AOI21_X1  g738(.A(G183gat), .B1(new_n919_), .B2(new_n932_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n935_), .A2(new_n936_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n939_), .B1(new_n940_), .B2(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n938_), .A2(new_n942_), .ZN(G1350gat));
  OAI21_X1  g742(.A(G190gat), .B1(new_n935_), .B2(new_n693_), .ZN(new_n944_));
  OR2_X1    g743(.A1(new_n657_), .A2(new_n342_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n944_), .B1(new_n935_), .B2(new_n945_), .ZN(G1351gat));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n947_));
  NOR4_X1   g746(.A1(new_n418_), .A2(new_n409_), .A3(new_n423_), .A4(new_n252_), .ZN(new_n948_));
  INV_X1    g747(.A(new_n948_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n947_), .B1(new_n869_), .B2(new_n949_), .ZN(new_n950_));
  OAI211_X1 g749(.A(KEYINPUT126), .B(new_n948_), .C1(new_n901_), .C2(new_n858_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n476_), .B1(new_n950_), .B2(new_n951_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n952_), .B(new_n290_), .ZN(G1352gat));
  AOI21_X1  g752(.A(new_n660_), .B1(new_n950_), .B2(new_n951_), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n954_), .B(new_n291_), .ZN(G1353gat));
  NAND2_X1  g754(.A1(new_n950_), .A2(new_n951_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n510_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n956_), .A2(new_n957_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n959_), .B(KEYINPUT127), .ZN(new_n960_));
  INV_X1    g759(.A(new_n960_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n958_), .A2(new_n961_), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n956_), .A2(new_n960_), .A3(new_n957_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n962_), .A2(new_n963_), .ZN(G1354gat));
  NAND3_X1  g763(.A1(new_n956_), .A2(new_n300_), .A3(new_n658_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n693_), .B1(new_n950_), .B2(new_n951_), .ZN(new_n966_));
  OAI21_X1  g765(.A(new_n965_), .B1(new_n300_), .B2(new_n966_), .ZN(G1355gat));
endmodule


