//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0 0 1 0 0 1 0 1 1 1 0 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n904_, new_n905_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n954_, new_n955_, new_n956_, new_n958_, new_n959_, new_n961_,
    new_n962_, new_n964_, new_n965_, new_n966_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n978_, new_n979_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT0), .B(G57gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G127gat), .B(G134gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G113gat), .B(G120gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT81), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n207_), .B(new_n208_), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n211_), .B1(new_n212_), .B2(new_n210_), .ZN(new_n213_));
  INV_X1    g012(.A(G141gat), .ZN(new_n214_));
  INV_X1    g013(.A(G148gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n218_));
  AND3_X1   g017(.A1(new_n216_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G155gat), .B(G162gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n219_), .B1(KEYINPUT1), .B2(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT84), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n223_), .B(new_n224_), .C1(G141gat), .C2(G148gat), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n214_), .B(new_n215_), .C1(KEYINPUT84), .C2(KEYINPUT3), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n222_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT85), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT85), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n230_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n220_), .B1(new_n227_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT86), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n221_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  AOI211_X1 g034(.A(KEYINPUT86), .B(new_n220_), .C1(new_n227_), .C2(new_n232_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n213_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n225_), .A2(new_n226_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n222_), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n238_), .A2(new_n239_), .A3(new_n229_), .A4(new_n231_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n220_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT86), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n233_), .A2(new_n234_), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n243_), .A2(new_n212_), .A3(new_n244_), .A4(new_n221_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n237_), .A2(new_n245_), .A3(KEYINPUT4), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G225gat), .A2(G233gat), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT4), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n249_), .B(new_n213_), .C1(new_n235_), .C2(new_n236_), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n246_), .A2(KEYINPUT93), .A3(new_n248_), .A4(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n237_), .A2(new_n245_), .A3(new_n247_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n250_), .A2(new_n248_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT93), .B1(new_n255_), .B2(new_n246_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n206_), .B1(new_n253_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT93), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n237_), .A2(new_n245_), .A3(KEYINPUT4), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n258_), .B1(new_n259_), .B2(new_n254_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n260_), .A2(new_n205_), .A3(new_n252_), .A4(new_n251_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n257_), .A2(KEYINPUT96), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT96), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n263_), .B(new_n206_), .C1(new_n253_), .C2(new_n256_), .ZN(new_n264_));
  OR2_X1    g063(.A1(G183gat), .A2(G190gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G183gat), .A2(G190gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT79), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT79), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n268_), .A2(G183gat), .A3(G190gat), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT23), .B1(new_n267_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n266_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT23), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n265_), .B1(new_n270_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT90), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT22), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n276_), .A2(G169gat), .ZN(new_n277_));
  INV_X1    g076(.A(G169gat), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n278_), .A2(KEYINPUT22), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n275_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(G176gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n278_), .A2(KEYINPUT22), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n276_), .A2(G169gat), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n282_), .A2(new_n283_), .A3(KEYINPUT90), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n280_), .A2(new_n281_), .A3(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT78), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n274_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT25), .B(G183gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT26), .B(G190gat), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT24), .ZN(new_n291_));
  NOR2_X1   g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292_));
  AOI22_X1  g091(.A1(new_n289_), .A2(new_n290_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n267_), .A2(new_n269_), .A3(KEYINPUT23), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT80), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n295_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n267_), .A2(new_n269_), .A3(new_n295_), .A4(KEYINPUT23), .ZN(new_n298_));
  INV_X1    g097(.A(new_n292_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n299_), .A2(KEYINPUT24), .A3(new_n286_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n293_), .A2(new_n297_), .A3(new_n298_), .A4(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n288_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT21), .ZN(new_n303_));
  AND2_X1   g102(.A1(G197gat), .A2(G204gat), .ZN(new_n304_));
  NOR2_X1   g103(.A1(G197gat), .A2(G204gat), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n303_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(G197gat), .ZN(new_n307_));
  INV_X1    g106(.A(G204gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G197gat), .A2(G204gat), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(KEYINPUT21), .A3(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G211gat), .B(G218gat), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n306_), .A2(new_n311_), .A3(KEYINPUT87), .A4(new_n312_), .ZN(new_n313_));
  AND3_X1   g112(.A1(new_n306_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT87), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n315_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n313_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n302_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n297_), .A2(new_n265_), .A3(new_n298_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT78), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n286_), .B(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n277_), .A2(new_n279_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n322_), .B1(new_n281_), .B2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n320_), .A2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n287_), .A2(KEYINPUT24), .A3(new_n299_), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n326_), .B(new_n293_), .C1(new_n273_), .C2(new_n270_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n325_), .A2(new_n327_), .A3(new_n317_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n319_), .A2(KEYINPUT20), .A3(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G226gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT19), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n325_), .A2(new_n327_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(new_n318_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n331_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n317_), .A2(new_n288_), .A3(new_n301_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n334_), .A2(KEYINPUT20), .A3(new_n335_), .A4(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n332_), .A2(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n338_), .A2(KEYINPUT95), .ZN(new_n339_));
  OR2_X1    g138(.A1(new_n329_), .A2(new_n331_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G8gat), .B(G36gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT92), .ZN(new_n344_));
  OR2_X1    g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n344_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G64gat), .B(G92gat), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n345_), .A2(new_n346_), .A3(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n348_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n342_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n351_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n353_), .A2(new_n341_), .A3(new_n349_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n355_), .A2(KEYINPUT32), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n334_), .A2(KEYINPUT20), .A3(new_n336_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(new_n331_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n340_), .A2(new_n356_), .A3(new_n358_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n332_), .A2(KEYINPUT95), .A3(new_n337_), .ZN(new_n360_));
  OAI22_X1  g159(.A1(new_n339_), .A2(new_n359_), .B1(new_n360_), .B2(new_n356_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n262_), .A2(new_n264_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT94), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT33), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n261_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n251_), .A2(new_n252_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n363_), .A2(new_n364_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n366_), .A2(new_n205_), .A3(new_n260_), .A4(new_n367_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n332_), .A2(new_n355_), .A3(new_n337_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n355_), .B1(new_n332_), .B2(new_n337_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n246_), .A2(new_n247_), .A3(new_n250_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n237_), .A2(new_n245_), .A3(new_n248_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(new_n206_), .A3(new_n373_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n365_), .A2(new_n368_), .A3(new_n371_), .A4(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n362_), .A2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G78gat), .B(G106gat), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT29), .B1(new_n235_), .B2(new_n236_), .ZN(new_n378_));
  INV_X1    g177(.A(G228gat), .ZN(new_n379_));
  INV_X1    g178(.A(G233gat), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n378_), .A2(new_n382_), .A3(new_n318_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n382_), .B1(new_n378_), .B2(new_n318_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n377_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n378_), .A2(new_n318_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(new_n381_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n378_), .A2(new_n382_), .A3(new_n318_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n377_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n387_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT88), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n385_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G22gat), .B(G50gat), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n243_), .A2(new_n244_), .A3(new_n221_), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT28), .B1(new_n394_), .B2(KEYINPUT29), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n235_), .A2(new_n236_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT28), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT29), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n396_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n393_), .B1(new_n395_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n395_), .A2(new_n399_), .A3(new_n393_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  OAI211_X1 g202(.A(KEYINPUT88), .B(new_n377_), .C1(new_n383_), .C2(new_n384_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n392_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n385_), .A2(KEYINPUT89), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n395_), .A2(new_n399_), .A3(new_n393_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n407_), .A2(new_n400_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT89), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n409_), .B(new_n377_), .C1(new_n383_), .C2(new_n384_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n406_), .A2(new_n408_), .A3(new_n410_), .A4(new_n390_), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n405_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n376_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT97), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n355_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n352_), .A2(new_n354_), .A3(KEYINPUT97), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n417_), .B1(new_n340_), .B2(new_n358_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT27), .ZN(new_n419_));
  NOR3_X1   g218(.A1(new_n418_), .A2(new_n369_), .A3(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n419_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT98), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  OAI211_X1 g222(.A(KEYINPUT98), .B(new_n419_), .C1(new_n369_), .C2(new_n370_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n420_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n405_), .A2(new_n411_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n262_), .A2(new_n264_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n425_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n413_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G227gat), .A2(G233gat), .ZN(new_n430_));
  INV_X1    g229(.A(G15gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G71gat), .B(G99gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(G43gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n433_), .A2(G43gat), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT30), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n433_), .A2(G43gat), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT30), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(new_n439_), .A3(new_n434_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n432_), .B1(new_n437_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n437_), .A2(new_n432_), .A3(new_n440_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n442_), .A2(new_n325_), .A3(new_n327_), .A4(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n443_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n333_), .B1(new_n445_), .B2(new_n441_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT82), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n444_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT31), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT31), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n444_), .A2(new_n446_), .A3(new_n447_), .A4(new_n450_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n449_), .A2(new_n213_), .A3(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n213_), .B1(new_n449_), .B2(new_n451_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  XOR2_X1   g253(.A(new_n454_), .B(KEYINPUT83), .Z(new_n455_));
  NAND4_X1  g254(.A1(new_n425_), .A2(new_n427_), .A3(new_n412_), .A4(new_n454_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT99), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n454_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n459_), .A2(new_n426_), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n460_), .A2(new_n425_), .A3(KEYINPUT99), .A4(new_n427_), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n429_), .A2(new_n455_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT13), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G230gat), .A2(G233gat), .ZN(new_n464_));
  INV_X1    g263(.A(G85gat), .ZN(new_n465_));
  INV_X1    g264(.A(G92gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G85gat), .A2(G92gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT8), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n471_), .A2(KEYINPUT64), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G99gat), .A2(G106gat), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT6), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT7), .ZN(new_n476_));
  INV_X1    g275(.A(G99gat), .ZN(new_n477_));
  INV_X1    g276(.A(G106gat), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n470_), .B(new_n472_), .C1(new_n475_), .C2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n473_), .B(KEYINPUT6), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n468_), .A2(KEYINPUT9), .ZN(new_n484_));
  OR2_X1    g283(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n478_), .A3(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n467_), .A2(KEYINPUT9), .A3(new_n468_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n483_), .A2(new_n484_), .A3(new_n487_), .A4(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n481_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n469_), .B1(new_n490_), .B2(new_n483_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT64), .B(KEYINPUT8), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n482_), .B(new_n489_), .C1(new_n491_), .C2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT66), .ZN(new_n496_));
  NAND2_X1  g295(.A1(KEYINPUT65), .A2(G71gat), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(KEYINPUT65), .A2(G71gat), .ZN(new_n499_));
  OAI21_X1  g298(.A(G78gat), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n499_), .ZN(new_n501_));
  INV_X1    g300(.A(G78gat), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n501_), .A2(new_n502_), .A3(new_n497_), .ZN(new_n503_));
  INV_X1    g302(.A(G64gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(G57gat), .ZN(new_n505_));
  INV_X1    g304(.A(G57gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(G64gat), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n505_), .A2(new_n507_), .A3(KEYINPUT11), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT11), .B1(new_n505_), .B2(new_n507_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n500_), .B(new_n503_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n505_), .A2(new_n507_), .A3(KEYINPUT11), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n502_), .B1(new_n501_), .B2(new_n497_), .ZN(new_n512_));
  NOR3_X1   g311(.A1(new_n498_), .A2(new_n499_), .A3(G78gat), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n511_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n496_), .B1(new_n510_), .B2(new_n514_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n510_), .A2(new_n514_), .A3(new_n496_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n495_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n510_), .A2(new_n514_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT66), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n510_), .A2(new_n514_), .A3(new_n496_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n519_), .A2(new_n494_), .A3(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n464_), .B1(new_n517_), .B2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G120gat), .B(G148gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT5), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G176gat), .B(G204gat), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n524_), .B(new_n525_), .Z(new_n526_));
  AOI21_X1  g325(.A(new_n494_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n464_), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT68), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT68), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n516_), .A2(new_n515_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n530_), .B(new_n464_), .C1(new_n531_), .C2(new_n494_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n494_), .A2(KEYINPUT67), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n470_), .B1(new_n475_), .B2(new_n481_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n492_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT67), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n536_), .A2(new_n537_), .A3(new_n482_), .A4(new_n489_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n534_), .A2(KEYINPUT12), .A3(new_n518_), .A4(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT12), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n521_), .A2(new_n540_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  AOI211_X1 g341(.A(new_n522_), .B(new_n526_), .C1(new_n533_), .C2(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(KEYINPUT70), .B1(new_n543_), .B2(KEYINPUT69), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n522_), .B1(new_n533_), .B2(new_n542_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n526_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT69), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT70), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n547_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n545_), .A2(new_n546_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n544_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n551_), .B1(new_n544_), .B2(new_n550_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n463_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NOR3_X1   g353(.A1(new_n543_), .A2(KEYINPUT69), .A3(KEYINPUT70), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n549_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n556_));
  OAI22_X1  g355(.A1(new_n555_), .A2(new_n556_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n544_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(KEYINPUT13), .A3(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n554_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G1gat), .B(G8gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT74), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G15gat), .B(G22gat), .ZN(new_n563_));
  INV_X1    g362(.A(G1gat), .ZN(new_n564_));
  INV_X1    g363(.A(G8gat), .ZN(new_n565_));
  OAI21_X1  g364(.A(KEYINPUT14), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n562_), .A2(new_n567_), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n561_), .A2(KEYINPUT74), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n561_), .A2(KEYINPUT74), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n569_), .A2(new_n566_), .A3(new_n563_), .A4(new_n570_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n568_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G29gat), .B(G36gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G43gat), .B(G50gat), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n574_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n572_), .B(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G229gat), .A2(G233gat), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n572_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT71), .B(KEYINPUT15), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n575_), .A2(new_n576_), .A3(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n583_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n582_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n572_), .A2(new_n577_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(new_n588_), .A3(new_n579_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n581_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G113gat), .B(G141gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT77), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G169gat), .B(G197gat), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n592_), .B(new_n593_), .Z(new_n594_));
  XNOR2_X1  g393(.A(new_n590_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G190gat), .B(G218gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G134gat), .B(G162gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT36), .Z(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n534_), .A2(new_n586_), .A3(new_n538_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n536_), .A2(new_n577_), .A3(new_n482_), .A4(new_n489_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G232gat), .A2(G233gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT34), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT35), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n602_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n601_), .A2(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n605_), .A2(new_n606_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n601_), .B(new_n608_), .C1(new_n606_), .C2(new_n605_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n600_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n598_), .A2(KEYINPUT36), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n611_), .A2(new_n614_), .A3(new_n612_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT72), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT72), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n611_), .A2(new_n617_), .A3(new_n612_), .A4(new_n614_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n613_), .B1(new_n616_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT37), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n616_), .A2(new_n618_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n599_), .B(KEYINPUT73), .ZN(new_n624_));
  INV_X1    g423(.A(new_n611_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n612_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n624_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n620_), .B1(new_n623_), .B2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n622_), .A2(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(G127gat), .B(G155gat), .Z(new_n630_));
  XNOR2_X1  g429(.A(G183gat), .B(G211gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT17), .ZN(new_n635_));
  AND2_X1   g434(.A1(G231gat), .A2(G233gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n572_), .B(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n531_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n637_), .A2(new_n638_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n635_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT17), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n634_), .A2(new_n642_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n518_), .B(KEYINPUT75), .Z(new_n644_));
  AOI21_X1  g443(.A(new_n643_), .B1(new_n637_), .B2(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n645_), .B1(new_n637_), .B2(new_n644_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n641_), .A2(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n629_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n560_), .A2(new_n595_), .A3(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n462_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n651_), .A2(KEYINPUT100), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(KEYINPUT100), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n427_), .A2(G1gat), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n652_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT38), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n652_), .A2(KEYINPUT38), .A3(new_n653_), .A4(new_n654_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n462_), .A2(new_n619_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n560_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n595_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n660_), .A2(new_n661_), .A3(new_n647_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n659_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n427_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(G1gat), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n657_), .A2(new_n658_), .A3(new_n666_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT101), .Z(G1324gat));
  INV_X1    g467(.A(KEYINPUT39), .ZN(new_n669_));
  INV_X1    g468(.A(new_n425_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n663_), .A2(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n669_), .B1(new_n671_), .B2(G8gat), .ZN(new_n672_));
  AOI211_X1 g471(.A(KEYINPUT39), .B(new_n565_), .C1(new_n663_), .C2(new_n670_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n652_), .A2(new_n653_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n670_), .A2(new_n565_), .ZN(new_n675_));
  OAI22_X1  g474(.A1(new_n672_), .A2(new_n673_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g476(.A(new_n455_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n431_), .B1(new_n663_), .B2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT41), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n650_), .A2(new_n431_), .A3(new_n678_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1326gat));
  INV_X1    g481(.A(G22gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n683_), .B1(new_n663_), .B2(new_n426_), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT42), .Z(new_n685_));
  NAND2_X1  g484(.A1(new_n426_), .A2(new_n683_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT102), .Z(new_n687_));
  OAI21_X1  g486(.A(new_n685_), .B1(new_n651_), .B2(new_n687_), .ZN(G1327gat));
  INV_X1    g487(.A(new_n613_), .ZN(new_n689_));
  AND4_X1   g488(.A1(KEYINPUT105), .A2(new_n623_), .A3(new_n647_), .A4(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT105), .B1(new_n619_), .B2(new_n647_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n552_), .A2(new_n553_), .A3(new_n463_), .ZN(new_n694_));
  AOI21_X1  g493(.A(KEYINPUT13), .B1(new_n557_), .B2(new_n558_), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n595_), .B(new_n693_), .C1(new_n694_), .C2(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(KEYINPUT106), .B1(new_n462_), .B2(new_n696_), .ZN(new_n697_));
  AOI211_X1 g496(.A(new_n661_), .B(new_n692_), .C1(new_n554_), .C2(new_n559_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n458_), .A2(new_n461_), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n425_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n426_), .B1(new_n362_), .B2(new_n375_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n455_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n699_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n698_), .A2(new_n703_), .A3(new_n704_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n697_), .A2(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G29gat), .B1(new_n706_), .B2(new_n664_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT104), .ZN(new_n708_));
  OAI21_X1  g507(.A(KEYINPUT103), .B1(new_n622_), .B2(new_n628_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT103), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n623_), .A2(new_n627_), .ZN(new_n711_));
  OAI211_X1 g510(.A(new_n710_), .B(new_n621_), .C1(new_n711_), .C2(new_n620_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n709_), .A2(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n713_), .B1(new_n699_), .B2(new_n702_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n629_), .A2(new_n715_), .ZN(new_n716_));
  OAI22_X1  g515(.A1(new_n714_), .A2(new_n715_), .B1(new_n462_), .B2(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n560_), .A2(new_n595_), .A3(new_n647_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n708_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT43), .B1(new_n462_), .B2(new_n713_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n703_), .A2(new_n715_), .A3(new_n629_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n718_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n725_), .A2(KEYINPUT104), .A3(KEYINPUT44), .ZN(new_n726_));
  AOI22_X1  g525(.A1(new_n722_), .A2(new_n726_), .B1(new_n721_), .B2(new_n720_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n664_), .A2(G29gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n707_), .B1(new_n727_), .B2(new_n728_), .ZN(G1328gat));
  AOI21_X1  g528(.A(KEYINPUT108), .B1(KEYINPUT109), .B2(KEYINPUT46), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n425_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n731_));
  AOI21_X1  g530(.A(KEYINPUT104), .B1(new_n725_), .B2(KEYINPUT44), .ZN(new_n732_));
  AND4_X1   g531(.A1(KEYINPUT104), .A2(new_n717_), .A3(KEYINPUT44), .A4(new_n719_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n731_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(G36gat), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n425_), .A2(G36gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n697_), .A2(new_n705_), .A3(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT107), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT107), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n697_), .A2(new_n705_), .A3(new_n739_), .A4(new_n736_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n738_), .A2(KEYINPUT45), .A3(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT45), .B1(new_n738_), .B2(new_n740_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n730_), .B1(new_n735_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n735_), .A2(new_n743_), .A3(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT109), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT46), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(G1329gat));
  AOI21_X1  g548(.A(G43gat), .B1(new_n706_), .B2(new_n678_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n454_), .A2(G43gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n727_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT47), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n752_), .B(new_n753_), .ZN(G1330gat));
  AOI21_X1  g553(.A(G50gat), .B1(new_n706_), .B2(new_n426_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n426_), .A2(G50gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n727_), .B2(new_n756_), .ZN(G1331gat));
  NOR3_X1   g556(.A1(new_n462_), .A2(new_n595_), .A3(new_n560_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n758_), .A2(new_n648_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n759_), .A2(new_n506_), .A3(new_n664_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n560_), .A2(new_n595_), .A3(new_n647_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n659_), .A2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(G57gat), .B1(new_n762_), .B2(new_n427_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n760_), .A2(new_n763_), .ZN(G1332gat));
  NAND3_X1  g563(.A1(new_n759_), .A2(new_n504_), .A3(new_n670_), .ZN(new_n765_));
  OAI21_X1  g564(.A(G64gat), .B1(new_n762_), .B2(new_n425_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n766_), .A2(KEYINPUT48), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(KEYINPUT48), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n765_), .B1(new_n767_), .B2(new_n768_), .ZN(G1333gat));
  INV_X1    g568(.A(G71gat), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n759_), .A2(new_n770_), .A3(new_n678_), .ZN(new_n771_));
  OAI21_X1  g570(.A(G71gat), .B1(new_n762_), .B2(new_n455_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n772_), .A2(KEYINPUT49), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(KEYINPUT49), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n771_), .B1(new_n773_), .B2(new_n774_), .ZN(G1334gat));
  NAND3_X1  g574(.A1(new_n759_), .A2(new_n502_), .A3(new_n426_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n659_), .A2(new_n426_), .A3(new_n761_), .ZN(new_n777_));
  XOR2_X1   g576(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n778_));
  AND3_X1   g577(.A1(new_n777_), .A2(G78gat), .A3(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n777_), .B2(G78gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n776_), .B1(new_n779_), .B2(new_n780_), .ZN(G1335gat));
  AND2_X1   g580(.A1(new_n758_), .A2(new_n693_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n782_), .A2(new_n465_), .A3(new_n664_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n717_), .A2(KEYINPUT111), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT111), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n723_), .A2(new_n786_), .A3(new_n724_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n647_), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n560_), .A2(new_n595_), .A3(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  OR3_X1    g589(.A1(new_n785_), .A2(new_n790_), .A3(KEYINPUT112), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT112), .B1(new_n785_), .B2(new_n790_), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n791_), .A2(new_n664_), .A3(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n783_), .B1(new_n793_), .B2(new_n465_), .ZN(G1336gat));
  NOR2_X1   g593(.A1(new_n425_), .A2(new_n466_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n791_), .A2(new_n792_), .A3(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(G92gat), .B1(new_n782_), .B2(new_n670_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n797_), .B(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n796_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT114), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT114), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n796_), .A2(new_n802_), .A3(new_n799_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n803_), .ZN(G1337gat));
  NAND4_X1  g603(.A1(new_n782_), .A2(new_n454_), .A3(new_n485_), .A4(new_n486_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n784_), .A2(new_n787_), .A3(new_n678_), .A4(new_n789_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n806_), .A2(KEYINPUT115), .A3(G99gat), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT115), .B1(new_n806_), .B2(G99gat), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n805_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g609(.A1(new_n717_), .A2(new_n426_), .A3(new_n789_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(G106gat), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(KEYINPUT52), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n782_), .A2(new_n478_), .A3(new_n426_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n815_), .B(new_n816_), .ZN(G1339gat));
  NAND3_X1  g616(.A1(new_n560_), .A2(new_n661_), .A3(new_n648_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n818_), .B(new_n819_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n661_), .A2(new_n543_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n533_), .A2(new_n542_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT117), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT55), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT117), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n825_), .B1(new_n533_), .B2(new_n542_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n542_), .A2(new_n517_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n528_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n824_), .A2(new_n828_), .A3(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(KEYINPUT56), .A3(new_n526_), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT56), .B1(new_n831_), .B2(new_n526_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n832_), .B1(new_n833_), .B2(KEYINPUT118), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n835_));
  AOI211_X1 g634(.A(new_n835_), .B(KEYINPUT56), .C1(new_n831_), .C2(new_n526_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n821_), .B1(new_n834_), .B2(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n590_), .A2(new_n594_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n587_), .A2(new_n588_), .A3(new_n580_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n594_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n840_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n838_), .B1(new_n839_), .B2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n557_), .A2(new_n558_), .A3(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n619_), .B1(new_n837_), .B2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT57), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846_));
  INV_X1    g645(.A(new_n843_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n828_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n830_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n526_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT56), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n835_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n833_), .A2(KEYINPUT118), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n854_), .A3(new_n832_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n847_), .B1(new_n855_), .B2(new_n821_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n846_), .B1(new_n856_), .B2(new_n619_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n842_), .A2(new_n547_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n858_), .B1(new_n852_), .B2(new_n832_), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n859_), .A2(KEYINPUT58), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(KEYINPUT58), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n629_), .A3(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n845_), .A2(new_n857_), .A3(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n820_), .B1(new_n863_), .B2(new_n647_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n670_), .A2(new_n427_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n460_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n864_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(G113gat), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n867_), .A2(new_n868_), .A3(new_n595_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n870_), .B1(new_n864_), .B2(new_n866_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n862_), .B1(new_n844_), .B2(KEYINPUT57), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n856_), .A2(new_n846_), .A3(new_n619_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n647_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n820_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n866_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n876_), .A2(KEYINPUT59), .A3(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n661_), .B1(new_n871_), .B2(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n869_), .B1(new_n879_), .B2(new_n868_), .ZN(G1340gat));
  INV_X1    g679(.A(KEYINPUT60), .ZN(new_n881_));
  AOI21_X1  g680(.A(KEYINPUT119), .B1(new_n881_), .B2(G120gat), .ZN(new_n882_));
  AOI21_X1  g681(.A(G120gat), .B1(new_n660_), .B2(new_n881_), .ZN(new_n883_));
  MUX2_X1   g682(.A(new_n882_), .B(KEYINPUT119), .S(new_n883_), .Z(new_n884_));
  NAND2_X1  g683(.A1(new_n867_), .A2(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n560_), .B1(new_n871_), .B2(new_n878_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n887_));
  OAI21_X1  g686(.A(G120gat), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  AOI211_X1 g687(.A(KEYINPUT120), .B(new_n560_), .C1(new_n871_), .C2(new_n878_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n885_), .B1(new_n888_), .B2(new_n889_), .ZN(G1341gat));
  INV_X1    g689(.A(G127gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n867_), .A2(new_n891_), .A3(new_n788_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n647_), .B1(new_n871_), .B2(new_n878_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n891_), .ZN(G1342gat));
  INV_X1    g693(.A(G134gat), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n867_), .A2(new_n895_), .A3(new_n619_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n629_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n897_), .B1(new_n871_), .B2(new_n878_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n896_), .B1(new_n898_), .B2(new_n895_), .ZN(G1343gat));
  NOR2_X1   g698(.A1(new_n678_), .A2(new_n412_), .ZN(new_n900_));
  AND3_X1   g699(.A1(new_n876_), .A2(new_n865_), .A3(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n595_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n660_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(KEYINPUT121), .B(G148gat), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n904_), .B(new_n905_), .ZN(G1345gat));
  XNOR2_X1  g705(.A(KEYINPUT61), .B(G155gat), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n909_), .B1(new_n901_), .B2(new_n788_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n900_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n864_), .A2(new_n911_), .ZN(new_n912_));
  AND4_X1   g711(.A1(new_n909_), .A2(new_n912_), .A3(new_n788_), .A4(new_n865_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n908_), .B1(new_n910_), .B2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n912_), .A2(new_n865_), .ZN(new_n915_));
  OAI21_X1  g714(.A(KEYINPUT122), .B1(new_n915_), .B2(new_n647_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n901_), .A2(new_n909_), .A3(new_n788_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n916_), .A2(new_n917_), .A3(new_n907_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n914_), .A2(new_n918_), .ZN(G1346gat));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n920_));
  AOI21_X1  g719(.A(G162gat), .B1(new_n901_), .B2(new_n619_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n713_), .ZN(new_n922_));
  AND4_X1   g721(.A1(G162gat), .A2(new_n912_), .A3(new_n922_), .A4(new_n865_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n920_), .B1(new_n921_), .B2(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(G162gat), .ZN(new_n925_));
  INV_X1    g724(.A(new_n619_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n925_), .B1(new_n915_), .B2(new_n926_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n901_), .A2(G162gat), .A3(new_n922_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n927_), .A2(KEYINPUT123), .A3(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n924_), .A2(new_n929_), .ZN(G1347gat));
  NOR2_X1   g729(.A1(new_n664_), .A2(new_n425_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n678_), .A2(new_n931_), .ZN(new_n932_));
  INV_X1    g731(.A(new_n932_), .ZN(new_n933_));
  NAND4_X1  g732(.A1(new_n876_), .A2(new_n412_), .A3(new_n595_), .A4(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(KEYINPUT124), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n426_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n937_));
  NAND4_X1  g736(.A1(new_n936_), .A2(new_n937_), .A3(new_n595_), .A4(new_n933_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n935_), .A2(G169gat), .A3(new_n938_), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n936_), .A2(new_n933_), .ZN(new_n942_));
  INV_X1    g741(.A(new_n942_), .ZN(new_n943_));
  NAND4_X1  g742(.A1(new_n943_), .A2(new_n280_), .A3(new_n284_), .A4(new_n595_), .ZN(new_n944_));
  NAND4_X1  g743(.A1(new_n935_), .A2(KEYINPUT62), .A3(G169gat), .A4(new_n938_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n941_), .A2(new_n944_), .A3(new_n945_), .ZN(G1348gat));
  AOI21_X1  g745(.A(G176gat), .B1(new_n943_), .B2(new_n660_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT125), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n936_), .A2(new_n948_), .ZN(new_n949_));
  OAI21_X1  g748(.A(KEYINPUT125), .B1(new_n864_), .B2(new_n426_), .ZN(new_n950_));
  AND2_X1   g749(.A1(new_n949_), .A2(new_n950_), .ZN(new_n951_));
  NOR3_X1   g750(.A1(new_n932_), .A2(new_n560_), .A3(new_n281_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n947_), .B1(new_n951_), .B2(new_n952_), .ZN(G1349gat));
  NOR3_X1   g752(.A1(new_n942_), .A2(new_n289_), .A3(new_n647_), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n951_), .A2(new_n788_), .A3(new_n933_), .ZN(new_n955_));
  INV_X1    g754(.A(G183gat), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n954_), .B1(new_n955_), .B2(new_n956_), .ZN(G1350gat));
  OAI21_X1  g756(.A(G190gat), .B1(new_n942_), .B2(new_n897_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n619_), .A2(new_n290_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n958_), .B1(new_n942_), .B2(new_n959_), .ZN(G1351gat));
  NAND2_X1  g759(.A1(new_n912_), .A2(new_n931_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n961_), .A2(new_n661_), .ZN(new_n962_));
  XNOR2_X1  g761(.A(new_n962_), .B(new_n307_), .ZN(G1352gat));
  NOR2_X1   g762(.A1(new_n961_), .A2(new_n560_), .ZN(new_n964_));
  OAI21_X1  g763(.A(new_n964_), .B1(KEYINPUT126), .B2(new_n308_), .ZN(new_n965_));
  XNOR2_X1  g764(.A(KEYINPUT126), .B(G204gat), .ZN(new_n966_));
  OAI21_X1  g765(.A(new_n965_), .B1(new_n964_), .B2(new_n966_), .ZN(G1353gat));
  INV_X1    g766(.A(KEYINPUT63), .ZN(new_n968_));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n969_));
  AOI21_X1  g768(.A(new_n647_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n970_));
  NAND4_X1  g769(.A1(new_n912_), .A2(new_n969_), .A3(new_n931_), .A4(new_n970_), .ZN(new_n971_));
  NAND4_X1  g770(.A1(new_n876_), .A2(new_n900_), .A3(new_n931_), .A4(new_n970_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n972_), .A2(KEYINPUT127), .ZN(new_n973_));
  INV_X1    g772(.A(G211gat), .ZN(new_n974_));
  AND4_X1   g773(.A1(new_n968_), .A2(new_n971_), .A3(new_n973_), .A4(new_n974_), .ZN(new_n975_));
  AOI22_X1  g774(.A1(new_n971_), .A2(new_n973_), .B1(new_n968_), .B2(new_n974_), .ZN(new_n976_));
  NOR2_X1   g775(.A1(new_n975_), .A2(new_n976_), .ZN(G1354gat));
  OAI21_X1  g776(.A(G218gat), .B1(new_n961_), .B2(new_n897_), .ZN(new_n978_));
  OR2_X1    g777(.A1(new_n926_), .A2(G218gat), .ZN(new_n979_));
  OAI21_X1  g778(.A(new_n978_), .B1(new_n961_), .B2(new_n979_), .ZN(G1355gat));
endmodule


