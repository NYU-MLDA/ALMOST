//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n620_, new_n621_, new_n622_, new_n623_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n827_, new_n828_, new_n829_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n841_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT15), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206_));
  INV_X1    g005(.A(G1gat), .ZN(new_n207_));
  INV_X1    g006(.A(G8gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n206_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G1gat), .B(G8gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n205_), .A2(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(new_n213_), .B(KEYINPUT77), .Z(new_n214_));
  NAND2_X1  g013(.A1(G229gat), .A2(G233gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n212_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n216_), .B1(new_n217_), .B2(new_n204_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  XOR2_X1   g018(.A(new_n212_), .B(new_n204_), .Z(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT76), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n219_), .B1(new_n221_), .B2(new_n215_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G113gat), .B(G141gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G169gat), .B(G197gat), .ZN(new_n224_));
  XOR2_X1   g023(.A(new_n223_), .B(new_n224_), .Z(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n222_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n222_), .A2(new_n226_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  XOR2_X1   g028(.A(new_n229_), .B(KEYINPUT78), .Z(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT89), .B(G106gat), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT21), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT88), .B(G204gat), .ZN(new_n235_));
  INV_X1    g034(.A(G197gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(G197gat), .A2(G204gat), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n234_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G211gat), .B(G218gat), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n235_), .A2(new_n236_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n234_), .B1(G197gat), .B2(G204gat), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n241_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n239_), .A2(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n237_), .A2(new_n238_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n240_), .A2(new_n234_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n245_), .A2(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(G155gat), .A2(G162gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G155gat), .A2(G162gat), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n250_), .B1(KEYINPUT1), .B2(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n252_), .B1(KEYINPUT1), .B2(new_n251_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G141gat), .A2(G148gat), .ZN(new_n254_));
  INV_X1    g053(.A(G141gat), .ZN(new_n255_));
  INV_X1    g054(.A(G148gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n253_), .A2(new_n254_), .A3(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(G155gat), .B(G162gat), .Z(new_n260_));
  INV_X1    g059(.A(KEYINPUT3), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT84), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n261_), .A2(new_n255_), .A3(new_n256_), .A4(KEYINPUT84), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(KEYINPUT85), .A2(KEYINPUT2), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(new_n254_), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT2), .ZN(new_n270_));
  AOI21_X1  g069(.A(KEYINPUT85), .B1(G141gat), .B2(G148gat), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n268_), .B(new_n269_), .C1(new_n270_), .C2(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n260_), .B1(new_n266_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT86), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  AOI22_X1  g074(.A1(new_n257_), .A2(KEYINPUT3), .B1(new_n267_), .B2(new_n254_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT85), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n254_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT2), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n276_), .A2(new_n264_), .A3(new_n279_), .A4(new_n265_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n280_), .A2(KEYINPUT86), .A3(new_n260_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n259_), .B1(new_n275_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT29), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n249_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(G22gat), .B(G50gat), .Z(new_n285_));
  OR2_X1    g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n285_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n282_), .A2(new_n283_), .ZN(new_n289_));
  XOR2_X1   g088(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n288_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n290_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n289_), .B(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n294_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G228gat), .A2(G233gat), .ZN(new_n296_));
  INV_X1    g095(.A(G78gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n292_), .A2(new_n295_), .A3(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n299_), .B1(new_n292_), .B2(new_n295_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n233_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n295_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n294_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n298_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n292_), .A2(new_n295_), .A3(new_n299_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n305_), .A2(new_n232_), .A3(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n302_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G127gat), .B(G134gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G113gat), .B(G120gat), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n311_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT83), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(KEYINPUT83), .B1(new_n312_), .B2(new_n313_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT31), .ZN(new_n319_));
  XOR2_X1   g118(.A(G71gat), .B(G99gat), .Z(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n322_));
  INV_X1    g121(.A(G169gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(G183gat), .ZN(new_n325_));
  INV_X1    g124(.A(G190gat), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT23), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT23), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n328_), .A2(G183gat), .A3(G190gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(G183gat), .A2(G190gat), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n324_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT79), .ZN(new_n334_));
  INV_X1    g133(.A(G176gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(new_n323_), .A3(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT79), .B1(G169gat), .B2(G176gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT24), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT25), .B(G183gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT26), .B(G190gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n329_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n327_), .A2(KEYINPUT81), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT81), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n347_), .B(KEYINPUT23), .C1(new_n325_), .C2(new_n326_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n345_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n344_), .A2(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n339_), .B1(G169gat), .B2(G176gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT80), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n333_), .B1(new_n350_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G227gat), .A2(G233gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(G15gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT30), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n355_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT82), .B(G43gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n321_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n321_), .A2(new_n361_), .ZN(new_n363_));
  AND2_X1   g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n309_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n351_), .A2(KEYINPUT90), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n367_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n351_), .A2(KEYINPUT90), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n343_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n340_), .A2(new_n330_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT91), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n340_), .A2(KEYINPUT91), .A3(new_n330_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n370_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n349_), .A2(new_n331_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n376_), .A2(new_n324_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n249_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT20), .ZN(new_n379_));
  AOI22_X1  g178(.A1(new_n239_), .A2(new_n244_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n379_), .B1(new_n355_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n378_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G226gat), .A2(G233gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT19), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT20), .B1(new_n355_), .B2(new_n380_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n373_), .A2(new_n374_), .ZN(new_n388_));
  OAI221_X1 g187(.A(new_n380_), .B1(new_n324_), .B2(new_n376_), .C1(new_n388_), .C2(new_n370_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n384_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n387_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(G8gat), .B(G36gat), .Z(new_n392_));
  XNOR2_X1  g191(.A(G64gat), .B(G92gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n385_), .A2(new_n391_), .A3(new_n396_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n397_), .A2(KEYINPUT27), .ZN(new_n398_));
  INV_X1    g197(.A(new_n396_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n382_), .A2(new_n384_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n390_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n399_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  NOR3_X1   g201(.A1(new_n375_), .A2(new_n377_), .A3(new_n249_), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n403_), .A2(new_n386_), .A3(new_n384_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n390_), .B1(new_n378_), .B2(new_n381_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n399_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n397_), .ZN(new_n407_));
  XOR2_X1   g206(.A(KEYINPUT98), .B(KEYINPUT27), .Z(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  AOI22_X1  g208(.A1(new_n398_), .A2(new_n402_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT100), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n366_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G1gat), .B(G29gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(G85gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT0), .B(G57gat), .ZN(new_n416_));
  XOR2_X1   g215(.A(new_n415_), .B(new_n416_), .Z(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n280_), .A2(KEYINPUT86), .A3(new_n260_), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT86), .B1(new_n280_), .B2(new_n260_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n258_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n314_), .B(new_n315_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT95), .B1(new_n423_), .B2(KEYINPUT4), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT95), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT4), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n421_), .A2(new_n422_), .A3(new_n425_), .A4(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n424_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G225gat), .A2(G233gat), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n314_), .B(new_n258_), .C1(new_n419_), .C2(new_n420_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n432_), .B(KEYINPUT93), .C1(new_n282_), .C2(new_n318_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT93), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n421_), .A2(new_n422_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT4), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT94), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n436_), .A2(KEYINPUT94), .A3(KEYINPUT4), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n431_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n436_), .A2(new_n429_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n418_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n429_), .B1(new_n424_), .B2(new_n427_), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT94), .B1(new_n436_), .B2(KEYINPUT4), .ZN(new_n446_));
  AOI211_X1 g245(.A(new_n438_), .B(new_n426_), .C1(new_n433_), .C2(new_n435_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n445_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n448_), .A2(new_n442_), .A3(new_n417_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n444_), .A2(KEYINPUT97), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT97), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n452_), .B(new_n418_), .C1(new_n441_), .C2(new_n443_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n451_), .A2(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n413_), .A2(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n400_), .A2(new_n401_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n385_), .A2(new_n391_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n396_), .A2(KEYINPUT32), .ZN(new_n459_));
  MUX2_X1   g258(.A(new_n457_), .B(new_n458_), .S(new_n459_), .Z(new_n460_));
  NAND3_X1  g259(.A1(new_n450_), .A2(new_n453_), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT33), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n449_), .A2(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n430_), .B1(new_n424_), .B2(new_n427_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n464_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n417_), .B1(new_n436_), .B2(new_n430_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n407_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n418_), .A2(new_n462_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n448_), .A2(new_n442_), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT96), .B1(new_n463_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n449_), .A2(new_n462_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT96), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n472_), .A2(new_n473_), .A3(new_n469_), .A4(new_n467_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n461_), .A2(new_n471_), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(new_n308_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n302_), .A2(new_n307_), .A3(new_n410_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n477_), .B1(new_n453_), .B2(new_n450_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n364_), .B1(new_n476_), .B2(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n456_), .B1(new_n480_), .B2(KEYINPUT99), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT99), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n478_), .B1(new_n475_), .B2(new_n308_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n482_), .B1(new_n483_), .B2(new_n364_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n231_), .B1(new_n481_), .B2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT8), .ZN(new_n486_));
  NOR2_X1   g285(.A1(G99gat), .A2(G106gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT7), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G99gat), .A2(G106gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT6), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT6), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n491_), .A2(G99gat), .A3(G106gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n488_), .A2(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(G85gat), .B(G92gat), .Z(new_n495_));
  AOI21_X1  g294(.A(new_n486_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT66), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n493_), .B(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n488_), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n495_), .A2(new_n486_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n496_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(KEYINPUT10), .B(G99gat), .Z(new_n502_));
  INV_X1    g301(.A(G106gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT65), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(G85gat), .ZN(new_n507_));
  INV_X1    g306(.A(G92gat), .ZN(new_n508_));
  NOR3_X1   g307(.A1(new_n507_), .A2(new_n508_), .A3(KEYINPUT9), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n509_), .B1(new_n495_), .B2(KEYINPUT9), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n506_), .A2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n501_), .B1(new_n511_), .B2(new_n498_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n204_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n506_), .A2(new_n498_), .A3(new_n510_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n499_), .A2(new_n500_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n514_), .B1(new_n515_), .B2(new_n496_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n205_), .ZN(new_n517_));
  XOR2_X1   g316(.A(KEYINPUT69), .B(KEYINPUT34), .Z(new_n518_));
  NAND2_X1  g317(.A1(G232gat), .A2(G233gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n513_), .B(new_n517_), .C1(KEYINPUT35), .C2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(KEYINPUT35), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(G190gat), .B(G218gat), .Z(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT70), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G134gat), .B(G162gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT36), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  XOR2_X1   g328(.A(new_n529_), .B(KEYINPUT71), .Z(new_n530_));
  AND2_X1   g329(.A1(new_n523_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n527_), .B(new_n528_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n523_), .A2(new_n532_), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT37), .B1(new_n533_), .B2(KEYINPUT72), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n212_), .B(KEYINPUT73), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G231gat), .A2(G233gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G57gat), .B(G64gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT11), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n542_), .B(KEYINPUT67), .Z(new_n543_));
  XOR2_X1   g342(.A(G71gat), .B(G78gat), .Z(new_n544_));
  OAI21_X1  g343(.A(new_n544_), .B1(KEYINPUT11), .B2(new_n541_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n543_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n540_), .B(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT74), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G127gat), .B(G155gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT16), .ZN(new_n550_));
  XOR2_X1   g349(.A(G183gat), .B(G211gat), .Z(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT17), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n548_), .B(new_n554_), .ZN(new_n555_));
  OR3_X1    g354(.A1(new_n547_), .A2(KEYINPUT17), .A3(new_n553_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT75), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n537_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G230gat), .A2(G233gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT64), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n543_), .B(new_n545_), .Z(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n516_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n512_), .A2(new_n546_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n563_), .A2(new_n564_), .A3(KEYINPUT12), .ZN(new_n565_));
  OR3_X1    g364(.A1(new_n512_), .A2(KEYINPUT12), .A3(new_n546_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n561_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT68), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n563_), .A2(new_n564_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(new_n561_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G120gat), .B(G148gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT5), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G176gat), .B(G204gat), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n573_), .B(new_n574_), .Z(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n569_), .A2(new_n571_), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n576_), .B1(new_n569_), .B2(new_n571_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n580_), .A2(KEYINPUT13), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(KEYINPUT13), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n559_), .A2(new_n583_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n485_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n585_), .A2(new_n207_), .A3(new_n455_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT38), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n588_), .B(KEYINPUT101), .Z(new_n589_));
  NAND2_X1  g388(.A1(new_n586_), .A2(new_n587_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT104), .ZN(new_n591_));
  INV_X1    g390(.A(new_n229_), .ZN(new_n592_));
  OAI21_X1  g391(.A(KEYINPUT102), .B1(new_n583_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT102), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n581_), .A2(new_n594_), .A3(new_n229_), .A4(new_n582_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n593_), .A2(new_n557_), .A3(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT103), .ZN(new_n597_));
  INV_X1    g396(.A(new_n534_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n598_), .B1(new_n481_), .B2(new_n484_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n455_), .ZN(new_n601_));
  OAI21_X1  g400(.A(G1gat), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n589_), .A2(new_n591_), .A3(new_n602_), .ZN(G1324gat));
  INV_X1    g402(.A(new_n412_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n597_), .A2(new_n604_), .A3(new_n599_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(G8gat), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT39), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT39), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n605_), .A2(new_n608_), .A3(G8gat), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n585_), .A2(new_n208_), .A3(new_n604_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(G1325gat));
  OAI21_X1  g413(.A(G15gat), .B1(new_n600_), .B2(new_n365_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT41), .Z(new_n616_));
  INV_X1    g415(.A(G15gat), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n585_), .A2(new_n617_), .A3(new_n364_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(G1326gat));
  OAI21_X1  g418(.A(G22gat), .B1(new_n600_), .B2(new_n308_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT42), .ZN(new_n621_));
  INV_X1    g420(.A(G22gat), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n585_), .A2(new_n622_), .A3(new_n309_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(G1327gat));
  NAND2_X1  g423(.A1(new_n455_), .A2(G29gat), .ZN(new_n625_));
  AOI211_X1 g424(.A(KEYINPUT43), .B(new_n537_), .C1(new_n481_), .C2(new_n484_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n476_), .A2(new_n479_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(KEYINPUT99), .A3(new_n365_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n456_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(new_n484_), .A3(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n627_), .B1(new_n631_), .B2(new_n536_), .ZN(new_n632_));
  OAI21_X1  g431(.A(KEYINPUT107), .B1(new_n626_), .B2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n536_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n627_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT107), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n633_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n558_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n593_), .A2(new_n640_), .A3(new_n595_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT44), .B1(new_n639_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT43), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n631_), .A2(new_n644_), .A3(new_n536_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n637_), .B1(new_n636_), .B2(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n632_), .A2(KEYINPUT107), .ZN(new_n647_));
  OAI211_X1 g446(.A(KEYINPUT44), .B(new_n642_), .C1(new_n646_), .C2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT108), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n641_), .B1(new_n633_), .B2(new_n638_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT108), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(new_n651_), .A3(KEYINPUT44), .ZN(new_n652_));
  AOI211_X1 g451(.A(new_n625_), .B(new_n643_), .C1(new_n649_), .C2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n583_), .ZN(new_n654_));
  AND4_X1   g453(.A1(new_n485_), .A2(new_n598_), .A3(new_n640_), .A4(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(new_n455_), .ZN(new_n656_));
  INV_X1    g455(.A(G29gat), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(KEYINPUT109), .B1(new_n653_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT109), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n649_), .A2(new_n652_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n643_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  OAI211_X1 g463(.A(new_n661_), .B(new_n658_), .C1(new_n664_), .C2(new_n625_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n660_), .A2(new_n665_), .ZN(G1328gat));
  INV_X1    g465(.A(KEYINPUT46), .ZN(new_n667_));
  INV_X1    g466(.A(G36gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n604_), .B1(new_n650_), .B2(KEYINPUT44), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n668_), .B1(new_n662_), .B2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n655_), .A2(new_n668_), .A3(new_n604_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT45), .Z(new_n673_));
  OAI21_X1  g472(.A(new_n667_), .B1(new_n671_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n673_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n669_), .B1(new_n649_), .B2(new_n652_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n675_), .B(KEYINPUT46), .C1(new_n676_), .C2(new_n668_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n674_), .A2(new_n677_), .ZN(G1329gat));
  NAND2_X1  g477(.A1(new_n364_), .A2(G43gat), .ZN(new_n679_));
  AOI211_X1 g478(.A(new_n679_), .B(new_n643_), .C1(new_n649_), .C2(new_n652_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n655_), .A2(new_n364_), .ZN(new_n681_));
  INV_X1    g480(.A(G43gat), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(KEYINPUT47), .B1(new_n680_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT47), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n686_), .B(new_n683_), .C1(new_n664_), .C2(new_n679_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(G1330gat));
  INV_X1    g487(.A(KEYINPUT110), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n309_), .A2(G50gat), .ZN(new_n690_));
  AOI211_X1 g489(.A(new_n690_), .B(new_n643_), .C1(new_n649_), .C2(new_n652_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n655_), .A2(new_n309_), .ZN(new_n692_));
  INV_X1    g491(.A(G50gat), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n689_), .B1(new_n691_), .B2(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(KEYINPUT110), .B(new_n694_), .C1(new_n664_), .C2(new_n690_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1331gat));
  NAND2_X1  g497(.A1(new_n631_), .A2(new_n592_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n699_), .A2(new_n559_), .A3(new_n654_), .ZN(new_n700_));
  INV_X1    g499(.A(G57gat), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n700_), .A2(new_n701_), .A3(new_n455_), .ZN(new_n702_));
  AND4_X1   g501(.A1(new_n231_), .A2(new_n599_), .A3(new_n558_), .A4(new_n583_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n703_), .A2(new_n455_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n702_), .B1(new_n704_), .B2(new_n701_), .ZN(G1332gat));
  INV_X1    g504(.A(G64gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n703_), .B2(new_n604_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT48), .Z(new_n708_));
  NAND3_X1  g507(.A1(new_n700_), .A2(new_n706_), .A3(new_n604_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1333gat));
  INV_X1    g509(.A(G71gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n711_), .B1(new_n703_), .B2(new_n364_), .ZN(new_n712_));
  XOR2_X1   g511(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n713_));
  XNOR2_X1  g512(.A(new_n712_), .B(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n364_), .A2(new_n711_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT112), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n700_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n714_), .A2(new_n717_), .ZN(G1334gat));
  AOI21_X1  g517(.A(new_n297_), .B1(new_n703_), .B2(new_n309_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n719_), .B(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n700_), .A2(new_n297_), .A3(new_n309_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1335gat));
  NOR4_X1   g522(.A1(new_n699_), .A2(new_n534_), .A3(new_n558_), .A4(new_n654_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n724_), .A2(new_n507_), .A3(new_n455_), .ZN(new_n725_));
  OAI21_X1  g524(.A(KEYINPUT114), .B1(new_n646_), .B2(new_n647_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT114), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n633_), .A2(new_n727_), .A3(new_n638_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n583_), .A2(new_n592_), .A3(new_n640_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT115), .Z(new_n730_));
  AND3_X1   g529(.A1(new_n726_), .A2(new_n728_), .A3(new_n730_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n731_), .A2(new_n455_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n725_), .B1(new_n732_), .B2(new_n507_), .ZN(G1336gat));
  NAND3_X1  g532(.A1(new_n724_), .A2(new_n508_), .A3(new_n604_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n731_), .A2(new_n604_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n735_), .B2(new_n508_), .ZN(G1337gat));
  NAND4_X1  g535(.A1(new_n726_), .A2(new_n364_), .A3(new_n728_), .A4(new_n730_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(G99gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n724_), .A2(new_n364_), .A3(new_n502_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  XOR2_X1   g539(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n741_));
  XNOR2_X1  g540(.A(new_n740_), .B(new_n741_), .ZN(G1338gat));
  NAND3_X1  g541(.A1(new_n724_), .A2(new_n503_), .A3(new_n309_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n639_), .A2(new_n309_), .A3(new_n730_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT52), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n744_), .A2(new_n745_), .A3(G106gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n744_), .B2(G106gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n743_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT53), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT53), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n750_), .B(new_n743_), .C1(new_n746_), .C2(new_n747_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(G1339gat));
  OAI21_X1  g551(.A(KEYINPUT117), .B1(new_n578_), .B2(new_n592_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT117), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n577_), .A2(new_n754_), .A3(new_n229_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT118), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT55), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n569_), .A2(new_n757_), .A3(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n565_), .A2(new_n566_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n561_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n568_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n567_), .A2(KEYINPUT68), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n763_), .A2(new_n758_), .A3(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT118), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n759_), .A2(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n760_), .A2(new_n761_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n768_), .B1(new_n567_), .B2(KEYINPUT55), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n770_), .A2(KEYINPUT56), .A3(new_n575_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT56), .ZN(new_n772_));
  INV_X1    g571(.A(new_n769_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n773_), .B1(new_n759_), .B2(new_n766_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n772_), .B1(new_n774_), .B2(new_n576_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n756_), .B1(new_n771_), .B2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n226_), .B1(new_n221_), .B2(new_n216_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n215_), .B1(new_n217_), .B2(new_n204_), .ZN(new_n778_));
  AOI22_X1  g577(.A1(new_n777_), .A2(KEYINPUT119), .B1(new_n214_), .B2(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n779_), .B1(KEYINPUT119), .B2(new_n777_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n227_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n580_), .A2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n534_), .B1(new_n776_), .B2(new_n782_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT57), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n771_), .A2(KEYINPUT120), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT120), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n770_), .A2(new_n786_), .A3(KEYINPUT56), .A4(new_n575_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n785_), .A2(new_n787_), .A3(new_n775_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n578_), .A2(new_n781_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT58), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n788_), .A2(KEYINPUT58), .A3(new_n789_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(new_n536_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n784_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n640_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n584_), .A2(new_n231_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n797_), .B(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n796_), .A2(new_n800_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n413_), .A2(KEYINPUT59), .A3(new_n601_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n413_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n557_), .B1(new_n784_), .B2(new_n794_), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n455_), .B(new_n804_), .C1(new_n805_), .C2(new_n799_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n806_), .A2(KEYINPUT121), .A3(KEYINPUT59), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT121), .B1(new_n806_), .B2(KEYINPUT59), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n230_), .B(new_n803_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(G113gat), .ZN(new_n810_));
  OR3_X1    g609(.A1(new_n806_), .A2(G113gat), .A3(new_n592_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(G1340gat));
  OAI211_X1 g611(.A(new_n583_), .B(new_n803_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(G120gat), .ZN(new_n814_));
  INV_X1    g613(.A(new_n806_), .ZN(new_n815_));
  INV_X1    g614(.A(G120gat), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(new_n654_), .B2(KEYINPUT60), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n815_), .B(new_n817_), .C1(KEYINPUT60), .C2(new_n816_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n814_), .A2(new_n818_), .ZN(G1341gat));
  AOI21_X1  g618(.A(G127gat), .B1(new_n815_), .B2(new_n558_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n808_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n806_), .A2(KEYINPUT121), .A3(KEYINPUT59), .ZN(new_n822_));
  AOI22_X1  g621(.A1(new_n821_), .A2(new_n822_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n823_));
  XOR2_X1   g622(.A(KEYINPUT122), .B(G127gat), .Z(new_n824_));
  AOI21_X1  g623(.A(new_n824_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n820_), .B1(new_n823_), .B2(new_n825_), .ZN(G1342gat));
  OAI211_X1 g625(.A(new_n536_), .B(new_n803_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(G134gat), .ZN(new_n828_));
  OR3_X1    g627(.A1(new_n806_), .A2(G134gat), .A3(new_n534_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(G1343gat));
  OR2_X1    g629(.A1(new_n805_), .A2(new_n799_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n831_), .A2(new_n455_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n308_), .A2(new_n364_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n833_), .A2(new_n412_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n836_), .A2(new_n255_), .A3(new_n229_), .ZN(new_n837_));
  OAI21_X1  g636(.A(G141gat), .B1(new_n835_), .B2(new_n592_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(G1344gat));
  NAND3_X1  g638(.A1(new_n836_), .A2(new_n256_), .A3(new_n583_), .ZN(new_n840_));
  OAI21_X1  g639(.A(G148gat), .B1(new_n835_), .B2(new_n654_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(G1345gat));
  XNOR2_X1  g641(.A(KEYINPUT61), .B(G155gat), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n836_), .A2(new_n558_), .A3(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n843_), .B1(new_n835_), .B2(new_n640_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(G1346gat));
  OAI21_X1  g646(.A(G162gat), .B1(new_n835_), .B2(new_n537_), .ZN(new_n848_));
  INV_X1    g647(.A(G162gat), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n598_), .A2(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n848_), .B1(new_n835_), .B2(new_n850_), .ZN(G1347gat));
  NAND3_X1  g650(.A1(new_n601_), .A2(new_n366_), .A3(new_n604_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n796_), .B2(new_n800_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n229_), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT62), .B1(new_n854_), .B2(KEYINPUT22), .ZN(new_n855_));
  OAI21_X1  g654(.A(G169gat), .B1(new_n854_), .B2(KEYINPUT62), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n323_), .B2(new_n855_), .ZN(G1348gat));
  INV_X1    g657(.A(new_n853_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n335_), .B1(new_n859_), .B2(new_n654_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n861_));
  INV_X1    g660(.A(new_n852_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n831_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n583_), .A2(G176gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n861_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n860_), .A2(new_n865_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n863_), .A2(new_n861_), .A3(new_n864_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1349gat));
  AND2_X1   g667(.A1(new_n831_), .A2(new_n862_), .ZN(new_n869_));
  AOI21_X1  g668(.A(G183gat), .B1(new_n869_), .B2(new_n558_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n341_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n557_), .A2(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n859_), .A2(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(KEYINPUT124), .B1(new_n870_), .B2(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n325_), .B1(new_n863_), .B2(new_n640_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT124), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n875_), .B(new_n876_), .C1(new_n859_), .C2(new_n872_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n874_), .A2(new_n877_), .ZN(G1350gat));
  AND3_X1   g677(.A1(new_n853_), .A2(new_n342_), .A3(new_n598_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n326_), .B1(new_n853_), .B2(new_n536_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT125), .ZN(new_n881_));
  OR3_X1    g680(.A1(new_n879_), .A2(new_n880_), .A3(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1351gat));
  NAND2_X1  g683(.A1(new_n601_), .A2(new_n833_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(KEYINPUT126), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n886_), .A2(new_n412_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n831_), .A2(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(new_n592_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(new_n236_), .ZN(G1352gat));
  AND2_X1   g689(.A1(new_n831_), .A2(new_n887_), .ZN(new_n891_));
  AOI21_X1  g690(.A(G204gat), .B1(new_n891_), .B2(new_n583_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n888_), .A2(new_n235_), .A3(new_n654_), .ZN(new_n893_));
  OAI21_X1  g692(.A(KEYINPUT127), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n235_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n891_), .A2(new_n895_), .A3(new_n583_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT127), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n888_), .A2(new_n654_), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n896_), .B(new_n897_), .C1(G204gat), .C2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n894_), .A2(new_n899_), .ZN(G1353gat));
  AOI211_X1 g699(.A(KEYINPUT63), .B(G211gat), .C1(new_n891_), .C2(new_n557_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n888_), .B1(new_n556_), .B2(new_n555_), .ZN(new_n902_));
  XOR2_X1   g701(.A(KEYINPUT63), .B(G211gat), .Z(new_n903_));
  AOI21_X1  g702(.A(new_n901_), .B1(new_n902_), .B2(new_n903_), .ZN(G1354gat));
  OAI21_X1  g703(.A(G218gat), .B1(new_n888_), .B2(new_n537_), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n534_), .A2(G218gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n888_), .B2(new_n906_), .ZN(G1355gat));
endmodule


