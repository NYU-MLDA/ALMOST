//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 1 1 0 1 1 0 1 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n920_, new_n922_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_;
  XOR2_X1   g000(.A(G1gat), .B(G8gat), .Z(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G15gat), .B(G22gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G1gat), .A2(G8gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT14), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT79), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT80), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT79), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n204_), .A2(new_n210_), .A3(new_n206_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n208_), .A2(new_n209_), .A3(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n209_), .B1(new_n208_), .B2(new_n211_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n203_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n208_), .A2(new_n211_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT80), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(new_n202_), .A3(new_n212_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n215_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G231gat), .A2(G233gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G57gat), .B(G64gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT11), .ZN(new_n222_));
  XOR2_X1   g021(.A(G71gat), .B(G78gat), .Z(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n221_), .A2(KEYINPUT11), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n222_), .A2(new_n223_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n220_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n220_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  OR3_X1    g029(.A1(new_n219_), .A2(new_n228_), .A3(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n219_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT17), .ZN(new_n234_));
  XOR2_X1   g033(.A(G127gat), .B(G155gat), .Z(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT16), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G183gat), .B(G211gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n233_), .A2(new_n234_), .A3(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n231_), .A2(new_n232_), .A3(KEYINPUT81), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n238_), .A2(new_n234_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  AND2_X1   g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n240_), .A2(new_n242_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n239_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT82), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G190gat), .B(G218gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G134gat), .B(G162gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT72), .ZN(new_n251_));
  INV_X1    g050(.A(G99gat), .ZN(new_n252_));
  INV_X1    g051(.A(G106gat), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(new_n253_), .A3(KEYINPUT70), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT70), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n255_), .B1(G99gat), .B2(G106gat), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT7), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n254_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G99gat), .A2(G106gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT6), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT6), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n264_), .A2(G99gat), .A3(G106gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  OAI211_X1 g065(.A(KEYINPUT69), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n258_), .A2(new_n261_), .A3(new_n266_), .A4(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT8), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n270_));
  INV_X1    g069(.A(G92gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(G85gat), .ZN(new_n272_));
  INV_X1    g071(.A(G85gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(G92gat), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n270_), .B1(new_n272_), .B2(new_n274_), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n268_), .A2(new_n269_), .A3(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n269_), .B1(new_n268_), .B2(new_n275_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT9), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n279_), .A2(new_n273_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n273_), .A2(KEYINPUT67), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT67), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(G85gat), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n281_), .A2(new_n283_), .A3(new_n279_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n280_), .B1(new_n284_), .B2(G92gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT68), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n266_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n288_));
  AND2_X1   g087(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT64), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT10), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(new_n252_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT64), .ZN(new_n294_));
  NAND2_X1  g093(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n291_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n253_), .A2(KEYINPUT65), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT65), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(G106gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT66), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT66), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n297_), .A2(new_n305_), .A3(new_n302_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n288_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n251_), .B1(new_n278_), .B2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G29gat), .B(G36gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G43gat), .B(G50gat), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n310_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT15), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n266_), .A2(new_n261_), .A3(new_n267_), .ZN(new_n315_));
  AND3_X1   g114(.A1(new_n254_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n275_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT8), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n268_), .A2(new_n269_), .A3(new_n275_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n286_), .B(KEYINPUT68), .Z(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT67), .B(G85gat), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n271_), .B1(new_n322_), .B2(new_n279_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n321_), .B1(new_n323_), .B2(new_n280_), .ZN(new_n324_));
  AOI211_X1 g123(.A(KEYINPUT66), .B(new_n301_), .C1(new_n296_), .C2(new_n291_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n305_), .B1(new_n297_), .B2(new_n302_), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n266_), .B(new_n324_), .C1(new_n325_), .C2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n320_), .A2(new_n327_), .A3(KEYINPUT72), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n308_), .A2(new_n314_), .A3(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G232gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT34), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT35), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT76), .ZN(new_n333_));
  OAI22_X1  g132(.A1(new_n333_), .A2(KEYINPUT78), .B1(KEYINPUT35), .B2(new_n331_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n278_), .A2(new_n307_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n334_), .B1(new_n335_), .B2(new_n313_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n333_), .A2(KEYINPUT78), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n329_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n337_), .B1(new_n329_), .B2(new_n336_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n250_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT36), .ZN(new_n342_));
  INV_X1    g141(.A(new_n340_), .ZN(new_n343_));
  AOI21_X1  g142(.A(KEYINPUT77), .B1(new_n343_), .B2(new_n338_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n341_), .B(new_n342_), .C1(new_n344_), .C2(new_n250_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n250_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n339_), .A2(new_n340_), .ZN(new_n347_));
  OAI211_X1 g146(.A(KEYINPUT36), .B(new_n346_), .C1(new_n347_), .C2(KEYINPUT77), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n247_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G226gat), .A2(G233gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT19), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT94), .ZN(new_n354_));
  INV_X1    g153(.A(G169gat), .ZN(new_n355_));
  INV_X1    g154(.A(G176gat), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT22), .B(G169gat), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n357_), .B1(new_n358_), .B2(new_n356_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n359_), .A2(KEYINPUT87), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G183gat), .A2(G190gat), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT23), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n363_), .B(new_n364_), .C1(G183gat), .C2(G190gat), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n360_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n359_), .A2(KEYINPUT87), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(G204gat), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n370_), .A2(G197gat), .ZN(new_n371_));
  INV_X1    g170(.A(G197gat), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n372_), .A2(G204gat), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT21), .B1(new_n371_), .B2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G211gat), .B(G218gat), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT92), .B1(new_n370_), .B2(G197gat), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT92), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n377_), .A2(new_n372_), .A3(G204gat), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n376_), .B(new_n378_), .C1(new_n372_), .C2(G204gat), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n374_), .B(new_n375_), .C1(new_n379_), .C2(KEYINPUT21), .ZN(new_n380_));
  INV_X1    g179(.A(new_n375_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(KEYINPUT21), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT24), .ZN(new_n385_));
  NOR2_X1   g184(.A1(G169gat), .A2(G176gat), .ZN(new_n386_));
  NOR3_X1   g185(.A1(new_n357_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n385_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n388_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT25), .B(G183gat), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT86), .ZN(new_n392_));
  INV_X1    g191(.A(G190gat), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n392_), .B1(new_n393_), .B2(KEYINPUT26), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT26), .B(G190gat), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n391_), .B(new_n394_), .C1(new_n395_), .C2(new_n392_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n390_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n369_), .A2(new_n384_), .A3(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n387_), .B1(new_n395_), .B2(new_n391_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT95), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n389_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n389_), .A2(new_n400_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n399_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n365_), .A2(KEYINPUT96), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n365_), .A2(KEYINPUT96), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n404_), .A2(new_n359_), .A3(new_n405_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n403_), .A2(new_n406_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n398_), .B(KEYINPUT20), .C1(new_n407_), .C2(KEYINPUT97), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(KEYINPUT97), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n354_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n384_), .A2(new_n403_), .A3(new_n406_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n412_), .A2(KEYINPUT98), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT20), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n369_), .A2(new_n397_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n414_), .B1(new_n415_), .B2(new_n383_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n353_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n412_), .A2(KEYINPUT98), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n413_), .A2(new_n416_), .A3(new_n417_), .A4(new_n418_), .ZN(new_n419_));
  XOR2_X1   g218(.A(G8gat), .B(G36gat), .Z(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G64gat), .B(G92gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT32), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n411_), .A2(new_n419_), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT102), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G155gat), .A2(G162gat), .ZN(new_n429_));
  OR2_X1    g228(.A1(G155gat), .A2(G162gat), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT89), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G141gat), .A2(G148gat), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT2), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n437_));
  INV_X1    g236(.A(G141gat), .ZN(new_n438_));
  INV_X1    g237(.A(G148gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n436_), .B(new_n437_), .C1(new_n440_), .C2(KEYINPUT3), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n429_), .B(new_n430_), .C1(new_n433_), .C2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT88), .B1(new_n429_), .B2(KEYINPUT1), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n429_), .A2(KEYINPUT1), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(new_n444_), .A3(new_n430_), .ZN(new_n445_));
  NOR3_X1   g244(.A1(new_n429_), .A2(KEYINPUT88), .A3(KEYINPUT1), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n434_), .B(new_n440_), .C1(new_n445_), .C2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n442_), .A2(new_n447_), .ZN(new_n448_));
  XOR2_X1   g247(.A(G127gat), .B(G134gat), .Z(new_n449_));
  XOR2_X1   g248(.A(G113gat), .B(G120gat), .Z(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n448_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n451_), .A2(new_n442_), .A3(new_n447_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G225gat), .A2(G233gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n453_), .A2(KEYINPUT4), .A3(new_n454_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n456_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT4), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n448_), .A2(new_n452_), .A3(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n458_), .A2(new_n459_), .A3(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n457_), .A2(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(G1gat), .B(G29gat), .Z(new_n464_));
  XNOR2_X1  g263(.A(G57gat), .B(G85gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT100), .B(KEYINPUT0), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n463_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n457_), .A2(new_n462_), .A3(new_n468_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n367_), .A2(new_n368_), .B1(new_n396_), .B2(new_n390_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT20), .B1(new_n473_), .B2(new_n384_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n412_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n353_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n403_), .A2(new_n406_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(new_n383_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT97), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n480_), .A2(KEYINPUT20), .A3(new_n409_), .A4(new_n398_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n476_), .B1(new_n481_), .B2(new_n354_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n425_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n411_), .A2(new_n419_), .A3(KEYINPUT102), .A4(new_n425_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n428_), .A2(new_n472_), .A3(new_n484_), .A4(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n411_), .A2(new_n419_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n424_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n471_), .A2(KEYINPUT33), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT33), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n457_), .A2(new_n462_), .A3(new_n491_), .A4(new_n468_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n411_), .A2(new_n419_), .A3(new_n424_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n458_), .A2(new_n456_), .A3(new_n461_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT101), .ZN(new_n496_));
  OR2_X1    g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n496_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n468_), .B1(new_n455_), .B2(new_n459_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n497_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n489_), .A2(new_n493_), .A3(new_n494_), .A4(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n486_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G227gat), .A2(G233gat), .ZN(new_n503_));
  INV_X1    g302(.A(G15gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT30), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT31), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G71gat), .B(G99gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(G43gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n415_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n473_), .A2(new_n510_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(new_n451_), .A3(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n451_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n508_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n512_), .A2(new_n513_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(new_n452_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n519_), .A2(new_n514_), .A3(new_n507_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n517_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G78gat), .B(G106gat), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT91), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n383_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT29), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n527_), .B1(new_n442_), .B2(new_n447_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G228gat), .A2(G233gat), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n526_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  OAI211_X1 g331(.A(G228gat), .B(G233gat), .C1(new_n525_), .C2(new_n528_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n523_), .B1(new_n532_), .B2(new_n534_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n442_), .A2(new_n447_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(new_n527_), .A3(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(G22gat), .B(G50gat), .Z(new_n540_));
  OAI21_X1  g339(.A(new_n537_), .B1(new_n448_), .B2(KEYINPUT29), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n540_), .B1(new_n539_), .B2(new_n541_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n523_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n531_), .A2(new_n533_), .A3(new_n545_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n535_), .A2(new_n544_), .A3(KEYINPUT93), .A4(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n535_), .A2(new_n546_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n544_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT93), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n546_), .A2(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n548_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n522_), .B1(new_n547_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n502_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n472_), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n552_), .A2(new_n521_), .A3(new_n547_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n521_), .B1(new_n552_), .B2(new_n547_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n555_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT103), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n494_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n494_), .A2(new_n559_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT27), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n562_), .B1(new_n482_), .B2(new_n488_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n560_), .A2(new_n561_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n489_), .A2(new_n494_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(new_n562_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n554_), .B1(new_n558_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT13), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n226_), .A2(new_n227_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n320_), .A2(new_n327_), .A3(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT73), .B(KEYINPUT12), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n227_), .B(new_n226_), .C1(new_n278_), .C2(new_n307_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G230gat), .A2(G233gat), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n226_), .A2(KEYINPUT12), .A3(new_n227_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n308_), .A2(new_n328_), .A3(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n575_), .A2(new_n576_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n574_), .A2(new_n571_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n576_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(G120gat), .B(G148gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(G176gat), .B(G204gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT74), .B(KEYINPUT5), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n580_), .A2(new_n583_), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n588_), .B1(new_n580_), .B2(new_n583_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n569_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n591_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n593_), .A2(KEYINPUT13), .A3(new_n589_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT83), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n313_), .A2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n311_), .A2(KEYINPUT83), .A3(new_n312_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n215_), .A2(new_n218_), .A3(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G229gat), .A2(G233gat), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n600_), .B1(new_n215_), .B2(new_n218_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n604_), .A2(KEYINPUT84), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT84), .ZN(new_n606_));
  AOI211_X1 g405(.A(new_n606_), .B(new_n600_), .C1(new_n215_), .C2(new_n218_), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n601_), .B(new_n603_), .C1(new_n605_), .C2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G113gat), .B(G141gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G169gat), .B(G197gat), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n609_), .B(new_n610_), .Z(new_n611_));
  NOR2_X1   g410(.A1(new_n611_), .A2(KEYINPUT85), .ZN(new_n612_));
  INV_X1    g411(.A(new_n314_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n219_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n600_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n219_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n606_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n604_), .A2(KEYINPUT84), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n614_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n608_), .B(new_n612_), .C1(new_n619_), .C2(new_n603_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  OAI22_X1  g420(.A1(new_n605_), .A2(new_n607_), .B1(new_n219_), .B2(new_n613_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(new_n602_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n612_), .B1(new_n623_), .B2(new_n608_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n621_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n596_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n351_), .A2(new_n568_), .A3(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(G1gat), .B1(new_n629_), .B2(new_n555_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT106), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n568_), .A2(new_n626_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT104), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n595_), .B(KEYINPUT75), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n345_), .A2(new_n348_), .A3(KEYINPUT37), .ZN(new_n637_));
  AOI21_X1  g436(.A(KEYINPUT37), .B1(new_n345_), .B2(new_n348_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(new_n246_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n634_), .A2(new_n636_), .A3(new_n641_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n642_), .A2(G1gat), .A3(new_n555_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(KEYINPUT38), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n644_), .A2(KEYINPUT105), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n644_), .A2(KEYINPUT105), .ZN(new_n646_));
  OAI221_X1 g445(.A(new_n631_), .B1(KEYINPUT38), .B2(new_n643_), .C1(new_n645_), .C2(new_n646_), .ZN(G1324gat));
  INV_X1    g446(.A(new_n567_), .ZN(new_n648_));
  OAI21_X1  g447(.A(G8gat), .B1(new_n629_), .B2(new_n648_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT39), .Z(new_n650_));
  NOR3_X1   g449(.A1(new_n642_), .A2(G8gat), .A3(new_n648_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT40), .ZN(G1325gat));
  OAI21_X1  g452(.A(G15gat), .B1(new_n629_), .B2(new_n521_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT41), .Z(new_n655_));
  NAND2_X1  g454(.A1(new_n522_), .A2(new_n504_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n655_), .B1(new_n642_), .B2(new_n656_), .ZN(G1326gat));
  INV_X1    g456(.A(new_n552_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n547_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G22gat), .B1(new_n629_), .B2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT42), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n661_), .A2(G22gat), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n663_), .B1(new_n642_), .B2(new_n664_), .ZN(G1327gat));
  NOR2_X1   g464(.A1(new_n246_), .A2(new_n349_), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n634_), .A2(new_n596_), .A3(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(G29gat), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n667_), .A2(new_n668_), .A3(new_n472_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT37), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n349_), .A2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n345_), .A2(new_n348_), .A3(KEYINPUT37), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(new_n568_), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n674_), .B1(new_n673_), .B2(new_n568_), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n247_), .B(new_n628_), .C1(new_n676_), .C2(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT44), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(new_n472_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n680_), .A2(KEYINPUT107), .A3(G29gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT107), .B1(new_n680_), .B2(G29gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n669_), .B1(new_n681_), .B2(new_n682_), .ZN(G1328gat));
  NOR2_X1   g482(.A1(new_n648_), .A2(G36gat), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n667_), .A2(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT45), .ZN(new_n686_));
  INV_X1    g485(.A(G36gat), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n679_), .A2(new_n567_), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n686_), .B(KEYINPUT46), .C1(new_n687_), .C2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT46), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT45), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n685_), .B(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n687_), .B1(new_n679_), .B2(new_n567_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n690_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n689_), .A2(new_n694_), .ZN(G1329gat));
  XOR2_X1   g494(.A(KEYINPUT108), .B(G43gat), .Z(new_n696_));
  AOI21_X1  g495(.A(new_n696_), .B1(new_n667_), .B2(new_n522_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n522_), .A2(G43gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n679_), .B2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT47), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n699_), .B(new_n700_), .ZN(G1330gat));
  AOI21_X1  g500(.A(G50gat), .B1(new_n667_), .B2(new_n660_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n660_), .A2(G50gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n679_), .B2(new_n703_), .ZN(G1331gat));
  AND2_X1   g503(.A1(new_n568_), .A2(new_n625_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n705_), .A2(new_n635_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(new_n351_), .ZN(new_n707_));
  OAI21_X1  g506(.A(G57gat), .B1(new_n707_), .B2(new_n555_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n641_), .A2(new_n595_), .A3(new_n705_), .ZN(new_n709_));
  INV_X1    g508(.A(G57gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n709_), .A2(new_n710_), .A3(new_n472_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n708_), .A2(new_n711_), .ZN(G1332gat));
  OAI21_X1  g511(.A(G64gat), .B1(new_n707_), .B2(new_n648_), .ZN(new_n713_));
  XOR2_X1   g512(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n714_));
  XNOR2_X1  g513(.A(new_n713_), .B(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(G64gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n709_), .A2(new_n716_), .A3(new_n567_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(G1333gat));
  OAI21_X1  g517(.A(G71gat), .B1(new_n707_), .B2(new_n521_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT49), .ZN(new_n720_));
  INV_X1    g519(.A(G71gat), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n709_), .A2(new_n721_), .A3(new_n522_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1334gat));
  INV_X1    g522(.A(G78gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n709_), .A2(new_n724_), .A3(new_n660_), .ZN(new_n725_));
  OAI21_X1  g524(.A(G78gat), .B1(new_n707_), .B2(new_n661_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(KEYINPUT50), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n726_), .A2(KEYINPUT50), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n725_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT110), .ZN(G1335gat));
  AND2_X1   g529(.A1(new_n706_), .A2(new_n666_), .ZN(new_n731_));
  AOI21_X1  g530(.A(G85gat), .B1(new_n731_), .B2(new_n472_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT111), .Z(new_n733_));
  NOR3_X1   g532(.A1(new_n246_), .A2(new_n626_), .A3(new_n596_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n673_), .A2(new_n568_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT43), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n735_), .B1(new_n737_), .B2(new_n675_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n739_), .A2(new_n555_), .A3(new_n322_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n733_), .A2(new_n740_), .ZN(G1336gat));
  OAI21_X1  g540(.A(G92gat), .B1(new_n739_), .B2(new_n648_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n731_), .A2(new_n271_), .A3(new_n567_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1337gat));
  AOI21_X1  g543(.A(new_n252_), .B1(new_n738_), .B2(new_n522_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n521_), .B1(new_n296_), .B2(new_n291_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n731_), .B2(new_n746_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n747_), .B(new_n748_), .ZN(G1338gat));
  OAI211_X1 g548(.A(new_n660_), .B(new_n734_), .C1(new_n676_), .C2(new_n677_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT114), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT114), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n738_), .A2(new_n752_), .A3(new_n660_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT115), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n751_), .A2(new_n753_), .A3(new_n754_), .A4(G106gat), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT52), .ZN(new_n756_));
  AOI211_X1 g555(.A(new_n661_), .B(new_n735_), .C1(new_n737_), .C2(new_n675_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n253_), .B1(new_n757_), .B2(new_n752_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n754_), .B1(new_n758_), .B2(new_n751_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n756_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n753_), .A2(G106gat), .ZN(new_n762_));
  INV_X1    g561(.A(new_n751_), .ZN(new_n763_));
  OAI211_X1 g562(.A(KEYINPUT115), .B(new_n761_), .C1(new_n762_), .C2(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n661_), .A2(new_n301_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n731_), .A2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT113), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n731_), .A2(new_n768_), .A3(new_n765_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n764_), .A2(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(KEYINPUT53), .B1(new_n760_), .B2(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT115), .B1(new_n762_), .B2(new_n763_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n773_), .A2(KEYINPUT52), .A3(new_n755_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n774_), .A2(new_n775_), .A3(new_n764_), .A4(new_n770_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n772_), .A2(new_n776_), .ZN(G1339gat));
  NOR2_X1   g576(.A1(new_n567_), .A2(new_n555_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n589_), .B1(new_n621_), .B2(new_n624_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT56), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n580_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n308_), .A2(new_n328_), .A3(new_n578_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n570_), .B1(new_n320_), .B2(new_n327_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n786_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n582_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n575_), .A2(new_n579_), .A3(KEYINPUT55), .A4(new_n576_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n782_), .B1(new_n580_), .B2(new_n783_), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n784_), .A2(new_n790_), .A3(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n781_), .B1(new_n792_), .B2(new_n588_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n788_), .A2(new_n789_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n580_), .A2(new_n783_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT117), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n580_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n794_), .A2(new_n796_), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n588_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(KEYINPUT56), .A3(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n780_), .B1(new_n793_), .B2(new_n800_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n601_), .B(new_n602_), .C1(new_n605_), .C2(new_n607_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n802_), .B1(new_n619_), .B2(new_n602_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n611_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n608_), .B1(new_n619_), .B2(new_n603_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n611_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n805_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n593_), .A2(new_n589_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  OAI211_X1 g610(.A(KEYINPUT57), .B(new_n349_), .C1(new_n801_), .C2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT118), .ZN(new_n813_));
  INV_X1    g612(.A(new_n780_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n798_), .A2(KEYINPUT56), .A3(new_n799_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT56), .B1(new_n798_), .B2(new_n799_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n814_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n810_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n818_), .A2(new_n819_), .A3(KEYINPUT57), .A4(new_n349_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n349_), .B1(new_n801_), .B2(new_n811_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n805_), .A2(new_n807_), .A3(new_n589_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n824_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT58), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  OAI211_X1 g626(.A(KEYINPUT58), .B(new_n824_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n827_), .A2(new_n673_), .A3(new_n828_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n813_), .A2(new_n820_), .A3(new_n823_), .A4(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n247_), .ZN(new_n831_));
  AND3_X1   g630(.A1(new_n625_), .A2(new_n592_), .A3(new_n594_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n671_), .A2(new_n246_), .A3(new_n832_), .A4(new_n672_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT116), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n639_), .A2(new_n835_), .A3(new_n246_), .A4(new_n832_), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n834_), .A2(new_n836_), .A3(KEYINPUT54), .ZN(new_n837_));
  AOI21_X1  g636(.A(KEYINPUT54), .B1(new_n834_), .B2(new_n836_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n779_), .B1(new_n831_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n557_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(G113gat), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n843_), .A3(new_n626_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n841_), .A2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n840_), .A2(KEYINPUT59), .A3(new_n557_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n625_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n844_), .B1(new_n848_), .B2(new_n843_), .ZN(G1340gat));
  INV_X1    g648(.A(G120gat), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n850_), .B1(new_n596_), .B2(KEYINPUT60), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n842_), .B(new_n851_), .C1(KEYINPUT60), .C2(new_n850_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n636_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n850_), .ZN(G1341gat));
  AOI21_X1  g653(.A(G127gat), .B1(new_n842_), .B2(new_n246_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n846_), .A2(new_n847_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(G127gat), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n246_), .A2(KEYINPUT119), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n858_), .B1(new_n859_), .B2(G127gat), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n855_), .B1(new_n856_), .B2(new_n860_), .ZN(G1342gat));
  AOI21_X1  g660(.A(G134gat), .B1(new_n842_), .B2(new_n350_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n673_), .A2(G134gat), .ZN(new_n863_));
  XOR2_X1   g662(.A(new_n863_), .B(KEYINPUT120), .Z(new_n864_));
  AOI21_X1  g663(.A(new_n862_), .B1(new_n856_), .B2(new_n864_), .ZN(G1343gat));
  NAND2_X1  g664(.A1(new_n831_), .A2(new_n839_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n778_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n556_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n867_), .A2(new_n625_), .A3(new_n868_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(new_n438_), .ZN(G1344gat));
  NOR3_X1   g669(.A1(new_n867_), .A2(new_n868_), .A3(new_n636_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(new_n439_), .ZN(G1345gat));
  NAND4_X1  g671(.A1(new_n866_), .A2(new_n556_), .A3(new_n246_), .A4(new_n778_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT121), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n840_), .A2(KEYINPUT121), .A3(new_n556_), .A4(new_n246_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(KEYINPUT61), .B(G155gat), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n875_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1346gat));
  NAND3_X1  g679(.A1(new_n840_), .A2(new_n556_), .A3(new_n350_), .ZN(new_n881_));
  INV_X1    g680(.A(G162gat), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n881_), .A2(KEYINPUT122), .A3(new_n882_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n867_), .A2(new_n868_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n639_), .A2(new_n882_), .ZN(new_n888_));
  AOI22_X1  g687(.A1(new_n885_), .A2(new_n886_), .B1(new_n887_), .B2(new_n888_), .ZN(G1347gat));
  NOR2_X1   g688(.A1(new_n648_), .A2(new_n472_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n891_), .B1(new_n831_), .B2(new_n839_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n892_), .A2(new_n626_), .A3(new_n557_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(G169gat), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT62), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n893_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n897_));
  INV_X1    g696(.A(new_n358_), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n896_), .B(new_n897_), .C1(new_n898_), .C2(new_n893_), .ZN(G1348gat));
  INV_X1    g698(.A(new_n557_), .ZN(new_n900_));
  AOI211_X1 g699(.A(new_n900_), .B(new_n891_), .C1(new_n831_), .C2(new_n839_), .ZN(new_n901_));
  AOI21_X1  g700(.A(G176gat), .B1(new_n901_), .B2(new_n595_), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n892_), .A2(G176gat), .A3(new_n557_), .A4(new_n635_), .ZN(new_n903_));
  OR2_X1    g702(.A1(new_n903_), .A2(KEYINPUT123), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(KEYINPUT123), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n902_), .B1(new_n904_), .B2(new_n905_), .ZN(G1349gat));
  NAND2_X1  g705(.A1(new_n901_), .A2(new_n246_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n391_), .ZN(new_n908_));
  INV_X1    g707(.A(G183gat), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n908_), .B1(new_n909_), .B2(new_n907_), .ZN(G1350gat));
  AOI21_X1  g709(.A(new_n393_), .B1(new_n901_), .B2(new_n673_), .ZN(new_n911_));
  AND4_X1   g710(.A1(new_n395_), .A2(new_n892_), .A3(new_n557_), .A4(new_n350_), .ZN(new_n912_));
  OAI21_X1  g711(.A(KEYINPUT124), .B1(new_n911_), .B2(new_n912_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n892_), .A2(new_n557_), .A3(new_n673_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(G190gat), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n901_), .A2(new_n395_), .A3(new_n350_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n915_), .A2(new_n916_), .A3(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n913_), .A2(new_n918_), .ZN(G1351gat));
  NAND3_X1  g718(.A1(new_n892_), .A2(new_n626_), .A3(new_n556_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g720(.A1(new_n866_), .A2(new_n890_), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n922_), .A2(new_n868_), .A3(new_n636_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(new_n370_), .ZN(G1353gat));
  NOR2_X1   g723(.A1(new_n922_), .A2(new_n868_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n925_), .A2(new_n246_), .A3(new_n926_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n928_));
  XOR2_X1   g727(.A(new_n928_), .B(KEYINPUT125), .Z(new_n929_));
  XOR2_X1   g728(.A(new_n929_), .B(KEYINPUT126), .Z(new_n930_));
  INV_X1    g729(.A(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n927_), .A2(new_n931_), .ZN(new_n932_));
  NAND4_X1  g731(.A1(new_n925_), .A2(new_n246_), .A3(new_n926_), .A4(new_n930_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1354gat));
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n935_));
  NAND4_X1  g734(.A1(new_n892_), .A2(new_n935_), .A3(new_n556_), .A4(new_n350_), .ZN(new_n936_));
  INV_X1    g735(.A(G218gat), .ZN(new_n937_));
  AND2_X1   g736(.A1(new_n936_), .A2(new_n937_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n892_), .A2(new_n556_), .A3(new_n350_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(KEYINPUT127), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n639_), .A2(new_n937_), .ZN(new_n941_));
  AOI22_X1  g740(.A1(new_n938_), .A2(new_n940_), .B1(new_n925_), .B2(new_n941_), .ZN(G1355gat));
endmodule


