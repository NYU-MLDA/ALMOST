//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 0 0 0 0 0 1 0 0 0 1 1 1 0 1 0 0 1 1 0 0 0 1 0 0 0 1 0 1 1 1 1 0 0 0 1 1 0 1 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n787_, new_n788_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n927_, new_n928_, new_n929_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n941_, new_n942_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_, new_n952_;
  INV_X1    g000(.A(KEYINPUT86), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT23), .ZN(new_n204_));
  INV_X1    g003(.A(G169gat), .ZN(new_n205_));
  INV_X1    g004(.A(G176gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n204_), .B1(KEYINPUT24), .B2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209_));
  AND3_X1   g008(.A1(new_n207_), .A2(KEYINPUT24), .A3(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  AND2_X1   g010(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT25), .ZN(new_n215_));
  INV_X1    g014(.A(G183gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT84), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT84), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(G183gat), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n215_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n221_));
  OAI211_X1 g020(.A(KEYINPUT85), .B(new_n214_), .C1(new_n220_), .C2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n221_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT84), .B(G183gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n224_), .B1(new_n225_), .B2(new_n215_), .ZN(new_n226_));
  AOI21_X1  g025(.A(KEYINPUT85), .B1(new_n226_), .B2(new_n214_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n211_), .B1(new_n223_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n225_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n204_), .B1(new_n229_), .B2(G190gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n205_), .A2(new_n206_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT22), .B(G169gat), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n231_), .B1(new_n232_), .B2(new_n206_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n230_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n228_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G71gat), .B(G99gat), .ZN(new_n236_));
  INV_X1    g035(.A(G43gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n235_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n235_), .A2(new_n238_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G227gat), .A2(G233gat), .ZN(new_n242_));
  INV_X1    g041(.A(G15gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT30), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT31), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n241_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n239_), .A2(new_n240_), .A3(new_n246_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n202_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G127gat), .B(G134gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G113gat), .B(G120gat), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n252_), .B(new_n253_), .Z(new_n254_));
  NAND3_X1  g053(.A1(new_n248_), .A2(new_n202_), .A3(new_n249_), .ZN(new_n255_));
  AND3_X1   g054(.A1(new_n251_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n254_), .B1(new_n251_), .B2(new_n255_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G141gat), .A2(G148gat), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(G141gat), .A2(G148gat), .ZN(new_n261_));
  NOR2_X1   g060(.A1(G155gat), .A2(G162gat), .ZN(new_n262_));
  INV_X1    g061(.A(G155gat), .ZN(new_n263_));
  INV_X1    g062(.A(G162gat), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT1), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n262_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT1), .B1(new_n263_), .B2(new_n264_), .ZN(new_n268_));
  AOI211_X1 g067(.A(new_n260_), .B(new_n261_), .C1(new_n267_), .C2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT87), .B(KEYINPUT2), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT88), .B1(new_n271_), .B2(new_n260_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT88), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT2), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n274_), .A2(KEYINPUT87), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n274_), .A2(KEYINPUT87), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n273_), .B(new_n259_), .C1(new_n275_), .C2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n261_), .A2(KEYINPUT3), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT3), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n279_), .B1(G141gat), .B2(G148gat), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n278_), .A2(new_n280_), .B1(new_n260_), .B2(KEYINPUT2), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n272_), .A2(new_n277_), .A3(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n265_), .A2(new_n262_), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n282_), .A2(KEYINPUT89), .A3(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(KEYINPUT89), .B1(new_n282_), .B2(new_n283_), .ZN(new_n285_));
  OAI211_X1 g084(.A(KEYINPUT98), .B(new_n270_), .C1(new_n284_), .C2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT97), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n254_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n286_), .A2(new_n287_), .A3(new_n254_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n282_), .A2(new_n283_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT89), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n282_), .A2(KEYINPUT89), .A3(new_n283_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n269_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT97), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n290_), .A2(KEYINPUT4), .A3(new_n291_), .A4(new_n297_), .ZN(new_n298_));
  NOR3_X1   g097(.A1(new_n296_), .A2(KEYINPUT4), .A3(new_n289_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G225gat), .A2(G233gat), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n290_), .A2(new_n291_), .A3(new_n297_), .A4(new_n300_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G1gat), .B(G29gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(G85gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT0), .B(G57gat), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n305_), .B(new_n306_), .Z(new_n307_));
  AND3_X1   g106(.A1(new_n302_), .A2(new_n303_), .A3(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n307_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n258_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT92), .B(G106gat), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  XOR2_X1   g112(.A(G197gat), .B(G204gat), .Z(new_n314_));
  AND2_X1   g113(.A1(KEYINPUT91), .A2(KEYINPUT21), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G211gat), .B(G218gat), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n314_), .A2(KEYINPUT21), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n314_), .A2(new_n315_), .A3(new_n317_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n270_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n322_), .B1(new_n323_), .B2(KEYINPUT29), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT28), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT29), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n325_), .B1(new_n296_), .B2(new_n326_), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n326_), .B(new_n270_), .C1(new_n284_), .C2(new_n285_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n328_), .A2(KEYINPUT28), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n324_), .B1(new_n327_), .B2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G22gat), .B(G50gat), .ZN(new_n331_));
  INV_X1    g130(.A(new_n322_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n332_), .B1(new_n296_), .B2(new_n326_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n328_), .A2(KEYINPUT28), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n296_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n333_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n330_), .A2(new_n331_), .A3(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n331_), .B1(new_n330_), .B2(new_n336_), .ZN(new_n338_));
  INV_X1    g137(.A(G228gat), .ZN(new_n339_));
  INV_X1    g138(.A(G233gat), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n340_), .A2(KEYINPUT90), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(KEYINPUT90), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n339_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(G78gat), .ZN(new_n344_));
  NOR3_X1   g143(.A1(new_n337_), .A2(new_n338_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n344_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n331_), .ZN(new_n347_));
  NOR3_X1   g146(.A1(new_n327_), .A2(new_n324_), .A3(new_n329_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n333_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n347_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n330_), .A2(new_n331_), .A3(new_n336_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n346_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n313_), .B1(new_n345_), .B2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n344_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n350_), .A2(new_n351_), .A3(new_n346_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(new_n355_), .A3(new_n312_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n353_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT27), .ZN(new_n358_));
  XOR2_X1   g157(.A(G8gat), .B(G36gat), .Z(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G64gat), .B(G92gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  AND2_X1   g163(.A1(KEYINPUT93), .A2(KEYINPUT24), .ZN(new_n365_));
  NOR2_X1   g164(.A1(KEYINPUT93), .A2(KEYINPUT24), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n207_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(new_n204_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  AND2_X1   g170(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n372_));
  OAI22_X1  g171(.A1(new_n213_), .A2(new_n212_), .B1(new_n372_), .B2(new_n221_), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n207_), .B(new_n209_), .C1(new_n365_), .C2(new_n366_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT94), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n373_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n375_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n371_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n204_), .B1(G183gat), .B2(G190gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(new_n233_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n378_), .A2(new_n322_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT20), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n322_), .B1(new_n228_), .B2(new_n234_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G226gat), .A2(G233gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT19), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n382_), .A2(new_n383_), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT95), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n228_), .A2(new_n322_), .A3(new_n234_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n373_), .A2(new_n374_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT94), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n373_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n370_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n380_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n332_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n388_), .A2(new_n394_), .A3(KEYINPUT20), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n385_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n386_), .B1(new_n387_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n385_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT20), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n378_), .A2(new_n380_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n399_), .B1(new_n400_), .B2(new_n332_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n398_), .B1(new_n401_), .B2(new_n388_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT95), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n364_), .B1(new_n397_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n235_), .A2(new_n332_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n405_), .A2(KEYINPUT20), .A3(new_n398_), .A4(new_n381_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n406_), .B1(new_n402_), .B2(KEYINPUT95), .ZN(new_n407_));
  AOI211_X1 g206(.A(new_n387_), .B(new_n398_), .C1(new_n401_), .C2(new_n388_), .ZN(new_n408_));
  NOR3_X1   g207(.A1(new_n407_), .A2(new_n408_), .A3(new_n363_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n358_), .B1(new_n404_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n396_), .A2(new_n387_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n411_), .A2(new_n403_), .A3(new_n364_), .A4(new_n406_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n385_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n401_), .A2(new_n398_), .A3(new_n388_), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n412_), .B(KEYINPUT27), .C1(new_n364_), .C2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n410_), .A2(new_n416_), .ZN(new_n417_));
  NOR3_X1   g216(.A1(new_n311_), .A2(new_n357_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT102), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n290_), .A2(new_n291_), .A3(new_n297_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT101), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n300_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n290_), .A2(KEYINPUT101), .A3(new_n291_), .A4(new_n297_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n422_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n299_), .A2(new_n423_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n307_), .B1(new_n298_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n363_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n429_), .A2(new_n412_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n302_), .A2(KEYINPUT33), .A3(new_n303_), .A4(new_n307_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n428_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n302_), .A2(new_n303_), .A3(new_n307_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT99), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT100), .B(KEYINPUT33), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n437_), .B1(new_n308_), .B2(KEYINPUT99), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n432_), .B1(new_n435_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n364_), .A2(KEYINPUT32), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n440_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n407_), .A2(new_n408_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n441_), .B1(new_n442_), .B2(new_n440_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n443_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n353_), .A2(new_n356_), .A3(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n439_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n302_), .A2(new_n303_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n307_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n410_), .A2(new_n449_), .A3(new_n433_), .A4(new_n416_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n354_), .A2(new_n355_), .A3(new_n312_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n312_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n450_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n258_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n419_), .B1(new_n446_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n429_), .A2(new_n412_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n457_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n435_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n436_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n458_), .B(new_n431_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n461_), .A2(new_n356_), .A3(new_n353_), .A4(new_n444_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n258_), .B1(new_n357_), .B2(new_n450_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(new_n463_), .A3(KEYINPUT102), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n418_), .B1(new_n456_), .B2(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(G85gat), .B(G92gat), .Z(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT7), .ZN(new_n468_));
  INV_X1    g267(.A(G99gat), .ZN(new_n469_));
  INV_X1    g268(.A(G106gat), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n468_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G99gat), .A2(G106gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT6), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT6), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n477_), .A2(G99gat), .A3(G106gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  AOI211_X1 g278(.A(KEYINPUT8), .B(new_n467_), .C1(new_n474_), .C2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT8), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT66), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n479_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n476_), .A2(new_n478_), .A3(KEYINPUT66), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(new_n474_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n466_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n481_), .B1(new_n486_), .B2(KEYINPUT67), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n473_), .B1(new_n482_), .B2(new_n479_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n467_), .B1(new_n488_), .B2(new_n484_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT67), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n480_), .B1(new_n487_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT9), .ZN(new_n493_));
  INV_X1    g292(.A(G85gat), .ZN(new_n494_));
  INV_X1    g293(.A(G92gat), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n493_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n496_), .B1(new_n466_), .B2(new_n493_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT65), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT10), .B(G99gat), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n479_), .B1(new_n500_), .B2(G106gat), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n492_), .A2(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(G29gat), .B(G36gat), .Z(new_n504_));
  XOR2_X1   g303(.A(G43gat), .B(G50gat), .Z(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT15), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n503_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G232gat), .A2(G233gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT34), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n511_), .A2(KEYINPUT35), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n503_), .A2(new_n506_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n509_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(KEYINPUT35), .A3(new_n511_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n511_), .A2(KEYINPUT35), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n509_), .A2(new_n516_), .A3(new_n512_), .A4(new_n513_), .ZN(new_n517_));
  AND2_X1   g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G190gat), .B(G218gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G134gat), .B(G162gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n521_), .A2(KEYINPUT36), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n518_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n515_), .A2(new_n517_), .ZN(new_n524_));
  XOR2_X1   g323(.A(new_n521_), .B(KEYINPUT36), .Z(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n465_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT13), .ZN(new_n530_));
  INV_X1    g329(.A(new_n480_), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT8), .B1(new_n489_), .B2(new_n490_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n486_), .A2(KEYINPUT67), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n531_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n502_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G57gat), .B(G64gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G71gat), .B(G78gat), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n537_), .A2(new_n538_), .A3(KEYINPUT11), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n537_), .A2(KEYINPUT11), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n540_), .A2(new_n538_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n537_), .A2(KEYINPUT11), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n539_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n536_), .A2(new_n544_), .ZN(new_n545_));
  OAI211_X1 g344(.A(KEYINPUT12), .B(new_n544_), .C1(new_n492_), .C2(new_n502_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT68), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT68), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n536_), .A2(new_n548_), .A3(KEYINPUT12), .A4(new_n544_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n545_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT69), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n543_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n551_), .B1(new_n552_), .B2(KEYINPUT12), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT12), .ZN(new_n554_));
  OAI211_X1 g353(.A(KEYINPUT69), .B(new_n554_), .C1(new_n503_), .C2(new_n543_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G230gat), .A2(G233gat), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n557_), .B(KEYINPUT64), .Z(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n550_), .A2(new_n556_), .A3(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n558_), .B1(new_n545_), .B2(new_n552_), .ZN(new_n561_));
  XOR2_X1   g360(.A(G120gat), .B(G148gat), .Z(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT71), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G176gat), .B(G204gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT72), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n563_), .B(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n560_), .A2(new_n561_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n569_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n530_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n560_), .A2(new_n561_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(new_n568_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n575_), .A2(KEYINPUT13), .A3(new_n570_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G113gat), .B(G141gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G169gat), .B(G197gat), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n578_), .B(new_n579_), .Z(new_n580_));
  NOR2_X1   g379(.A1(new_n580_), .A2(KEYINPUT82), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT74), .B(G1gat), .ZN(new_n584_));
  INV_X1    g383(.A(G8gat), .ZN(new_n585_));
  OAI21_X1  g384(.A(KEYINPUT14), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G1gat), .B(G8gat), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G15gat), .B(G22gat), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n586_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n588_), .B1(new_n586_), .B2(new_n589_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n583_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n592_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(new_n582_), .A3(new_n590_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n596_), .A2(new_n508_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT81), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n506_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G229gat), .A2(G233gat), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n598_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT80), .ZN(new_n602_));
  INV_X1    g401(.A(new_n506_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n593_), .A2(new_n595_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n603_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n606_));
  OAI21_X1  g405(.A(KEYINPUT79), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT79), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n599_), .A2(new_n608_), .A3(new_n604_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n600_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n602_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  AOI211_X1 g411(.A(KEYINPUT80), .B(new_n600_), .C1(new_n607_), .C2(new_n609_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n601_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT83), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT83), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n601_), .B(new_n616_), .C1(new_n612_), .C2(new_n613_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n581_), .B1(new_n615_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n615_), .A2(new_n581_), .A3(new_n617_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n577_), .A2(KEYINPUT104), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT104), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n615_), .A2(new_n581_), .A3(new_n617_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(new_n618_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n573_), .A2(new_n576_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n623_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G231gat), .A2(G233gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT77), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n596_), .B(new_n629_), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n630_), .A2(new_n544_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n544_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(G127gat), .B(G155gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT16), .ZN(new_n635_));
  XOR2_X1   g434(.A(G183gat), .B(G211gat), .Z(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT17), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n638_), .A2(KEYINPUT17), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n633_), .A2(new_n640_), .A3(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT78), .ZN(new_n643_));
  INV_X1    g442(.A(new_n633_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n643_), .B1(new_n644_), .B2(new_n639_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n633_), .A2(KEYINPUT78), .A3(new_n640_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n642_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n622_), .A2(new_n627_), .A3(new_n647_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n529_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n310_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n527_), .A2(KEYINPUT37), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT37), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n525_), .B(KEYINPUT73), .Z(new_n654_));
  NAND2_X1  g453(.A1(new_n524_), .A2(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n653_), .B1(new_n523_), .B2(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n652_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n658_), .A2(new_n577_), .A3(new_n647_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n465_), .A2(new_n659_), .A3(new_n625_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n660_), .A2(new_n650_), .A3(new_n584_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT38), .ZN(new_n662_));
  AOI22_X1  g461(.A1(new_n651_), .A2(G1gat), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n661_), .A2(new_n662_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n664_), .A2(KEYINPUT103), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(KEYINPUT103), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n663_), .B1(new_n665_), .B2(new_n666_), .ZN(G1324gat));
  INV_X1    g466(.A(KEYINPUT40), .ZN(new_n668_));
  INV_X1    g467(.A(new_n418_), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n446_), .A2(new_n455_), .A3(new_n419_), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT102), .B1(new_n462_), .B2(new_n463_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n669_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n672_), .A2(new_n648_), .A3(new_n417_), .A4(new_n527_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT105), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n529_), .A2(new_n675_), .A3(new_n417_), .A4(new_n648_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n674_), .A2(new_n676_), .A3(G8gat), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n674_), .A2(new_n676_), .A3(KEYINPUT106), .A4(G8gat), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n679_), .A2(KEYINPUT39), .A3(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT39), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n677_), .A2(new_n678_), .A3(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n660_), .A2(new_n585_), .A3(new_n417_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n668_), .B1(new_n681_), .B2(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n679_), .A2(KEYINPUT39), .A3(new_n680_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n687_), .A2(KEYINPUT40), .A3(new_n684_), .A4(new_n683_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(G1325gat));
  NAND3_X1  g488(.A1(new_n660_), .A2(new_n243_), .A3(new_n258_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n649_), .A2(new_n258_), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n691_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(KEYINPUT41), .B1(new_n691_), .B2(G15gat), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n690_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT107), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n696_), .B(new_n690_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(G1326gat));
  INV_X1    g497(.A(G22gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n699_), .B1(new_n649_), .B2(new_n357_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT42), .Z(new_n701_));
  NAND3_X1  g500(.A1(new_n660_), .A2(new_n699_), .A3(new_n357_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1327gat));
  NOR3_X1   g502(.A1(new_n626_), .A2(new_n527_), .A3(new_n647_), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n672_), .A2(new_n621_), .A3(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(G29gat), .B1(new_n705_), .B2(new_n650_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n647_), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n622_), .A2(new_n627_), .A3(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n672_), .B2(new_n657_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n465_), .A2(KEYINPUT43), .A3(new_n658_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n708_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n713_), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n708_), .B(new_n715_), .C1(new_n710_), .C2(new_n711_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n714_), .A2(new_n716_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n650_), .A2(G29gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n706_), .B1(new_n717_), .B2(new_n718_), .ZN(G1328gat));
  INV_X1    g518(.A(KEYINPUT109), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT46), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n714_), .A2(new_n417_), .A3(new_n716_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(G36gat), .ZN(new_n725_));
  INV_X1    g524(.A(new_n417_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n726_), .A2(G36gat), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n672_), .A2(new_n621_), .A3(new_n704_), .A4(new_n727_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n728_), .A2(KEYINPUT45), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n728_), .A2(KEYINPUT45), .ZN(new_n730_));
  OAI22_X1  g529(.A1(new_n729_), .A2(new_n730_), .B1(KEYINPUT109), .B2(KEYINPUT46), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n723_), .B1(new_n725_), .B2(new_n732_), .ZN(new_n733_));
  AOI211_X1 g532(.A(new_n722_), .B(new_n731_), .C1(new_n724_), .C2(G36gat), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1329gat));
  NAND4_X1  g534(.A1(new_n714_), .A2(G43gat), .A3(new_n258_), .A4(new_n716_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n705_), .A2(new_n258_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n237_), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n736_), .A2(KEYINPUT47), .A3(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(KEYINPUT47), .B1(new_n736_), .B2(new_n738_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1330gat));
  AOI21_X1  g540(.A(G50gat), .B1(new_n705_), .B2(new_n357_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n357_), .A2(G50gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n717_), .B2(new_n743_), .ZN(G1331gat));
  NAND2_X1  g543(.A1(new_n626_), .A2(new_n647_), .ZN(new_n745_));
  NOR4_X1   g544(.A1(new_n465_), .A2(new_n621_), .A3(new_n528_), .A4(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n746_), .A2(G57gat), .A3(new_n650_), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n747_), .B(KEYINPUT112), .Z(new_n748_));
  NOR2_X1   g547(.A1(new_n657_), .A2(new_n745_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT110), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n465_), .A2(new_n621_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(new_n650_), .ZN(new_n753_));
  INV_X1    g552(.A(G57gat), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n753_), .A2(KEYINPUT111), .A3(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT111), .B1(new_n753_), .B2(new_n754_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n748_), .A2(new_n755_), .A3(new_n756_), .ZN(G1332gat));
  INV_X1    g556(.A(G64gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n746_), .B2(new_n417_), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT48), .Z(new_n760_));
  NAND3_X1  g559(.A1(new_n752_), .A2(new_n758_), .A3(new_n417_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(G1333gat));
  INV_X1    g561(.A(G71gat), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n752_), .A2(new_n763_), .A3(new_n258_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT49), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n746_), .A2(new_n258_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(G71gat), .ZN(new_n767_));
  AOI211_X1 g566(.A(KEYINPUT49), .B(new_n763_), .C1(new_n746_), .C2(new_n258_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT113), .Z(G1334gat));
  INV_X1    g569(.A(G78gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n771_), .B1(new_n746_), .B2(new_n357_), .ZN(new_n772_));
  XOR2_X1   g571(.A(new_n772_), .B(KEYINPUT50), .Z(new_n773_));
  NAND3_X1  g572(.A1(new_n752_), .A2(new_n771_), .A3(new_n357_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(G1335gat));
  AND4_X1   g574(.A1(new_n626_), .A2(new_n751_), .A3(new_n528_), .A4(new_n707_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n776_), .A2(new_n494_), .A3(new_n650_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n577_), .A2(new_n621_), .A3(new_n647_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n672_), .A2(new_n709_), .A3(new_n657_), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT43), .B1(new_n465_), .B2(new_n658_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n779_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n782_), .A2(KEYINPUT114), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n782_), .A2(KEYINPUT114), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n783_), .A2(new_n784_), .A3(new_n310_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n777_), .B1(new_n785_), .B2(new_n494_), .ZN(G1336gat));
  NAND3_X1  g585(.A1(new_n776_), .A2(new_n495_), .A3(new_n417_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n783_), .A2(new_n784_), .A3(new_n726_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n788_), .B2(new_n495_), .ZN(G1337gat));
  INV_X1    g588(.A(new_n500_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n776_), .A2(new_n258_), .A3(new_n790_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n782_), .A2(new_n258_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(new_n469_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g593(.A1(new_n776_), .A2(new_n470_), .A3(new_n357_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n782_), .A2(new_n357_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(G106gat), .ZN(new_n798_));
  AOI211_X1 g597(.A(KEYINPUT52), .B(new_n470_), .C1(new_n782_), .C2(new_n357_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n795_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT53), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n802_), .B(new_n795_), .C1(new_n798_), .C2(new_n799_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n803_), .ZN(G1339gat));
  OR4_X1    g603(.A1(new_n357_), .A2(new_n310_), .A3(new_n417_), .A4(new_n454_), .ZN(new_n805_));
  XOR2_X1   g604(.A(new_n805_), .B(KEYINPUT119), .Z(new_n806_));
  INV_X1    g605(.A(KEYINPUT58), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n559_), .B1(new_n550_), .B2(new_n556_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n560_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n550_), .A2(new_n556_), .A3(KEYINPUT55), .A4(new_n559_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n812_), .A2(KEYINPUT56), .A3(new_n568_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n569_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n815_), .A2(KEYINPUT56), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n814_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n611_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n819_));
  OR3_X1    g618(.A1(new_n819_), .A2(KEYINPUT117), .A3(new_n580_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n598_), .A2(new_n599_), .A3(new_n611_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT117), .B1(new_n819_), .B2(new_n580_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n820_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n601_), .B(new_n580_), .C1(new_n612_), .C2(new_n613_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n818_), .B1(new_n825_), .B2(new_n571_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n823_), .A2(new_n570_), .A3(KEYINPUT118), .A4(new_n824_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n807_), .B1(new_n817_), .B2(new_n828_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n826_), .A2(new_n827_), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n830_), .B(KEYINPUT58), .C1(new_n816_), .C2(new_n814_), .ZN(new_n831_));
  AND3_X1   g630(.A1(new_n829_), .A2(new_n657_), .A3(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n621_), .A2(new_n570_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n812_), .A2(new_n568_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT56), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n834_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT115), .B1(new_n815_), .B2(KEYINPUT56), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n815_), .A2(KEYINPUT116), .A3(KEYINPUT56), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT116), .B1(new_n815_), .B2(KEYINPUT56), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n833_), .B1(new_n839_), .B2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n825_), .B1(new_n575_), .B2(new_n570_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n527_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n832_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  OAI211_X1 g647(.A(KEYINPUT57), .B(new_n527_), .C1(new_n844_), .C2(new_n845_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n647_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n658_), .A2(new_n625_), .A3(new_n577_), .A4(new_n647_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n851_), .B(new_n852_), .ZN(new_n853_));
  OAI211_X1 g652(.A(KEYINPUT59), .B(new_n806_), .C1(new_n850_), .C2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n813_), .A2(new_n856_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n837_), .A2(new_n857_), .A3(new_n838_), .A4(new_n840_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n625_), .A2(new_n571_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n845_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n847_), .B1(new_n860_), .B2(new_n528_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n829_), .A2(new_n657_), .A3(new_n831_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n849_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n853_), .B1(new_n863_), .B2(new_n707_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n806_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n855_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n625_), .B1(new_n854_), .B2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(G113gat), .ZN(new_n868_));
  INV_X1    g667(.A(new_n864_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n806_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n621_), .A2(new_n868_), .ZN(new_n871_));
  OAI22_X1  g670(.A1(new_n867_), .A2(new_n868_), .B1(new_n870_), .B2(new_n871_), .ZN(G1340gat));
  AOI21_X1  g671(.A(new_n577_), .B1(new_n854_), .B2(new_n866_), .ZN(new_n873_));
  INV_X1    g672(.A(G120gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n874_), .B1(new_n577_), .B2(KEYINPUT60), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n875_), .B1(KEYINPUT60), .B2(new_n874_), .ZN(new_n876_));
  OAI22_X1  g675(.A1(new_n873_), .A2(new_n874_), .B1(new_n870_), .B2(new_n876_), .ZN(G1341gat));
  AOI21_X1  g676(.A(new_n707_), .B1(new_n854_), .B2(new_n866_), .ZN(new_n878_));
  INV_X1    g677(.A(G127gat), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n647_), .A2(new_n879_), .ZN(new_n880_));
  OAI22_X1  g679(.A1(new_n878_), .A2(new_n879_), .B1(new_n870_), .B2(new_n880_), .ZN(G1342gat));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n864_), .A2(new_n527_), .A3(new_n865_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(G134gat), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n528_), .B(new_n806_), .C1(new_n850_), .C2(new_n853_), .ZN(new_n885_));
  INV_X1    g684(.A(G134gat), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n885_), .A2(KEYINPUT120), .A3(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n854_), .A2(new_n866_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n657_), .A2(G134gat), .ZN(new_n889_));
  XOR2_X1   g688(.A(new_n889_), .B(KEYINPUT121), .Z(new_n890_));
  AOI22_X1  g689(.A1(new_n884_), .A2(new_n887_), .B1(new_n888_), .B2(new_n890_), .ZN(G1343gat));
  NAND2_X1  g690(.A1(new_n454_), .A2(new_n357_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n892_), .A2(new_n310_), .A3(new_n417_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n864_), .A2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n621_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n626_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(KEYINPUT122), .B(G148gat), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(G1345gat));
  NAND2_X1  g699(.A1(new_n895_), .A2(new_n647_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT61), .B(G155gat), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1346gat));
  NOR3_X1   g702(.A1(new_n864_), .A2(new_n527_), .A3(new_n894_), .ZN(new_n904_));
  OAI21_X1  g703(.A(KEYINPUT123), .B1(new_n904_), .B2(G162gat), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n528_), .B(new_n893_), .C1(new_n850_), .C2(new_n853_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n906_), .A2(new_n907_), .A3(new_n264_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n658_), .A2(new_n264_), .ZN(new_n909_));
  AOI22_X1  g708(.A1(new_n905_), .A2(new_n908_), .B1(new_n895_), .B2(new_n909_), .ZN(G1347gat));
  NOR3_X1   g709(.A1(new_n311_), .A2(new_n357_), .A3(new_n726_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n869_), .A2(new_n621_), .A3(new_n911_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n912_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n914_));
  INV_X1    g713(.A(new_n911_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n864_), .A2(new_n625_), .A3(new_n915_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n914_), .B1(new_n916_), .B2(new_n205_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n232_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n913_), .A2(new_n917_), .A3(new_n918_), .ZN(G1348gat));
  OR2_X1    g718(.A1(new_n206_), .A2(KEYINPUT124), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n206_), .A2(KEYINPUT124), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n864_), .A2(new_n915_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  OAI211_X1 g722(.A(new_n920_), .B(new_n921_), .C1(new_n923_), .C2(new_n577_), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n922_), .A2(KEYINPUT124), .A3(new_n206_), .A4(new_n626_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(G1349gat));
  AOI21_X1  g725(.A(new_n229_), .B1(new_n922_), .B2(new_n647_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n923_), .A2(new_n707_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n372_), .A2(new_n221_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n927_), .B1(new_n928_), .B2(new_n929_), .ZN(G1350gat));
  NAND2_X1  g729(.A1(new_n528_), .A2(new_n214_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(KEYINPUT125), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n864_), .A2(new_n658_), .A3(new_n915_), .ZN(new_n933_));
  INV_X1    g732(.A(G190gat), .ZN(new_n934_));
  OAI22_X1  g733(.A1(new_n923_), .A2(new_n932_), .B1(new_n933_), .B2(new_n934_), .ZN(G1351gat));
  NOR3_X1   g734(.A1(new_n892_), .A2(new_n650_), .A3(new_n726_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n864_), .A2(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(new_n621_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(G197gat), .ZN(G1352gat));
  AOI21_X1  g739(.A(new_n577_), .B1(KEYINPUT126), .B2(G204gat), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n938_), .A2(new_n941_), .ZN(new_n942_));
  OR2_X1    g741(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n942_), .B(new_n943_), .ZN(G1353gat));
  AOI21_X1  g743(.A(new_n707_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n938_), .A2(new_n945_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n947_));
  XOR2_X1   g746(.A(new_n947_), .B(KEYINPUT127), .Z(new_n948_));
  XNOR2_X1  g747(.A(new_n946_), .B(new_n948_), .ZN(G1354gat));
  INV_X1    g748(.A(G218gat), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n938_), .A2(new_n950_), .A3(new_n528_), .ZN(new_n951_));
  NOR3_X1   g750(.A1(new_n864_), .A2(new_n658_), .A3(new_n937_), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n951_), .B1(new_n950_), .B2(new_n952_), .ZN(G1355gat));
endmodule


