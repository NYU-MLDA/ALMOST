//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 0 0 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n772_, new_n773_, new_n774_, new_n775_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n784_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n933_, new_n934_, new_n935_, new_n937_,
    new_n938_, new_n940_, new_n941_, new_n942_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT34), .Z(new_n203_));
  INV_X1    g002(.A(KEYINPUT35), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G85gat), .A2(G92gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G85gat), .A2(G92gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT66), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(G85gat), .A2(G92gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT66), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n211_), .A2(new_n212_), .A3(new_n207_), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(KEYINPUT68), .A2(KEYINPUT6), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(KEYINPUT68), .A2(KEYINPUT6), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n216_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT68), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT6), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(new_n215_), .A3(new_n217_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT7), .ZN(new_n225_));
  INV_X1    g024(.A(G99gat), .ZN(new_n226_));
  INV_X1    g025(.A(G106gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n220_), .A2(new_n224_), .A3(new_n228_), .A4(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n214_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT8), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT8), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n210_), .A2(new_n213_), .A3(new_n233_), .ZN(new_n234_));
  AND2_X1   g033(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n235_));
  NOR2_X1   g034(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n216_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  OR2_X1    g036(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n238_));
  NAND2_X1  g037(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(new_n215_), .A3(new_n239_), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n237_), .A2(new_n240_), .A3(new_n228_), .A4(new_n229_), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n234_), .A2(new_n241_), .A3(KEYINPUT67), .ZN(new_n242_));
  AOI21_X1  g041(.A(KEYINPUT67), .B1(new_n234_), .B2(new_n241_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n232_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G29gat), .B(G36gat), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT72), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n245_), .A2(new_n246_), .ZN(new_n248_));
  XOR2_X1   g047(.A(G43gat), .B(G50gat), .Z(new_n249_));
  OR3_X1    g048(.A1(new_n247_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n249_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n211_), .A2(new_n207_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT9), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  AND3_X1   g056(.A1(new_n255_), .A2(KEYINPUT64), .A3(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(KEYINPUT64), .B1(new_n255_), .B2(new_n257_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT10), .B(G99gat), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n237_), .B(new_n240_), .C1(G106gat), .C2(new_n260_), .ZN(new_n261_));
  NOR3_X1   g060(.A1(new_n258_), .A2(new_n259_), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n244_), .A2(new_n253_), .A3(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT74), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n244_), .A2(new_n253_), .A3(new_n263_), .A4(KEYINPUT74), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(KEYINPUT73), .B(KEYINPUT15), .Z(new_n269_));
  NOR2_X1   g068(.A1(new_n252_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n269_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n271_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n233_), .B1(new_n214_), .B2(new_n230_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n276_));
  AND4_X1   g075(.A1(new_n228_), .A2(new_n237_), .A3(new_n240_), .A4(new_n229_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n210_), .A2(new_n213_), .A3(new_n233_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n276_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n234_), .A2(new_n241_), .A3(KEYINPUT67), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n275_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n274_), .B1(new_n281_), .B2(new_n262_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n244_), .A2(new_n263_), .A3(KEYINPUT71), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n273_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n203_), .A2(new_n204_), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n285_), .B(KEYINPUT75), .Z(new_n286_));
  INV_X1    g085(.A(KEYINPUT77), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  AND4_X1   g087(.A1(new_n206_), .A2(new_n268_), .A3(new_n284_), .A4(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n288_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n290_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n206_), .B1(new_n291_), .B2(new_n284_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G190gat), .B(G218gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT76), .ZN(new_n294_));
  XOR2_X1   g093(.A(G134gat), .B(G162gat), .Z(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT36), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NOR3_X1   g097(.A1(new_n289_), .A2(new_n292_), .A3(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n296_), .B(new_n297_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n268_), .A2(new_n284_), .A3(new_n288_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n205_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n291_), .A2(new_n206_), .A3(new_n284_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n300_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n299_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G1gat), .B(G29gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT0), .ZN(new_n307_));
  INV_X1    g106(.A(G57gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(G85gat), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT4), .ZN(new_n311_));
  INV_X1    g110(.A(G155gat), .ZN(new_n312_));
  INV_X1    g111(.A(G162gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n312_), .A2(new_n313_), .A3(KEYINPUT88), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT88), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n315_), .B1(G155gat), .B2(G162gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G155gat), .A2(G162gat), .ZN(new_n317_));
  AND3_X1   g116(.A1(new_n314_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT90), .ZN(new_n319_));
  INV_X1    g118(.A(G141gat), .ZN(new_n320_));
  INV_X1    g119(.A(G148gat), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT3), .ZN(new_n323_));
  NOR2_X1   g122(.A1(G141gat), .A2(G148gat), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT3), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(new_n319_), .A3(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n323_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  AND3_X1   g127(.A1(KEYINPUT87), .A2(G141gat), .A3(G148gat), .ZN(new_n329_));
  AOI21_X1  g128(.A(KEYINPUT87), .B1(G141gat), .B2(G148gat), .ZN(new_n330_));
  NOR3_X1   g129(.A1(new_n329_), .A2(new_n330_), .A3(KEYINPUT2), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n318_), .B1(new_n328_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT97), .ZN(new_n333_));
  AND3_X1   g132(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n334_));
  AOI21_X1  g133(.A(KEYINPUT1), .B1(G155gat), .B2(G162gat), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n314_), .B(new_n316_), .C1(new_n334_), .C2(new_n335_), .ZN(new_n336_));
  NOR3_X1   g135(.A1(new_n329_), .A2(new_n330_), .A3(new_n324_), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n336_), .A2(new_n337_), .A3(KEYINPUT89), .ZN(new_n338_));
  AOI21_X1  g137(.A(KEYINPUT89), .B1(new_n336_), .B2(new_n337_), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n332_), .B(new_n333_), .C1(new_n338_), .C2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G127gat), .B(G134gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G113gat), .B(G120gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n336_), .A2(new_n337_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT89), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n336_), .A2(new_n337_), .A3(KEYINPUT89), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n343_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n349_), .A2(new_n333_), .A3(new_n350_), .A4(new_n332_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n311_), .B1(new_n344_), .B2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n332_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n353_), .A2(new_n311_), .A3(new_n350_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n352_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n355_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n344_), .A2(new_n351_), .ZN(new_n359_));
  AOI211_X1 g158(.A(new_n310_), .B(new_n357_), .C1(new_n358_), .C2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n355_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT98), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n359_), .A2(KEYINPUT4), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n354_), .A2(new_n358_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n362_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  NOR3_X1   g165(.A1(new_n352_), .A2(KEYINPUT98), .A3(new_n364_), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n361_), .B(new_n310_), .C1(new_n366_), .C2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT33), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n363_), .A2(new_n362_), .A3(new_n365_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT98), .B1(new_n352_), .B2(new_n364_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT33), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n372_), .A2(new_n373_), .A3(new_n361_), .A4(new_n310_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n360_), .B1(new_n369_), .B2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G226gat), .A2(G233gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT19), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT22), .B(G169gat), .ZN(new_n378_));
  INV_X1    g177(.A(G176gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G183gat), .A2(G190gat), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT23), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n383_), .B(new_n384_), .C1(G183gat), .C2(G190gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G169gat), .A2(G176gat), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n380_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT25), .B(G183gat), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT26), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(G190gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT83), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n388_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(G190gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT26), .ZN(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT83), .B1(new_n390_), .B2(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n392_), .A2(new_n395_), .ZN(new_n396_));
  OR2_X1    g195(.A1(G169gat), .A2(G176gat), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n397_), .A2(KEYINPUT24), .A3(new_n386_), .ZN(new_n398_));
  NOR3_X1   g197(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n398_), .A2(new_n400_), .A3(new_n383_), .A4(new_n384_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n387_), .B1(new_n396_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT84), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT84), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n387_), .B(new_n404_), .C1(new_n396_), .C2(new_n401_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(G211gat), .B(G218gat), .Z(new_n407_));
  INV_X1    g206(.A(G197gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n408_), .A2(KEYINPUT92), .A3(G204gat), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT92), .ZN(new_n410_));
  INV_X1    g209(.A(G204gat), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n410_), .B1(new_n411_), .B2(G197gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT91), .B(G197gat), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n409_), .B(new_n412_), .C1(new_n413_), .C2(G204gat), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n407_), .B1(new_n414_), .B2(KEYINPUT21), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n408_), .A2(KEYINPUT91), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT91), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(G197gat), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n416_), .A2(new_n418_), .A3(G204gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT93), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT21), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT93), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n416_), .A2(new_n418_), .A3(new_n422_), .A4(G204gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n411_), .A2(G197gat), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n420_), .A2(new_n421_), .A3(new_n423_), .A4(new_n424_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n415_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n407_), .A2(KEYINPUT21), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT94), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n423_), .A2(new_n424_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n422_), .B1(new_n413_), .B2(G204gat), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n428_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n420_), .A2(KEYINPUT94), .A3(new_n423_), .A4(new_n424_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n427_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NOR3_X1   g232(.A1(new_n406_), .A2(new_n426_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n431_), .A2(new_n432_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n427_), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n435_), .A2(new_n436_), .B1(new_n425_), .B2(new_n415_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n383_), .A2(new_n384_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n438_), .A2(new_n399_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n388_), .A2(new_n390_), .A3(new_n394_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n440_), .A3(new_n398_), .ZN(new_n441_));
  AND2_X1   g240(.A1(new_n441_), .A2(new_n387_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT20), .B1(new_n437_), .B2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n377_), .B1(new_n434_), .B2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G8gat), .B(G36gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(KEYINPUT18), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT95), .ZN(new_n447_));
  XOR2_X1   g246(.A(G64gat), .B(G92gat), .Z(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n406_), .B1(new_n426_), .B2(new_n433_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n437_), .A2(new_n442_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n377_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n451_), .A2(new_n452_), .A3(KEYINPUT20), .A4(new_n453_), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n444_), .A2(new_n450_), .A3(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n450_), .B1(new_n444_), .B2(new_n454_), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT96), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n444_), .A2(new_n454_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n449_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT96), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n444_), .A2(new_n450_), .A3(new_n454_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n457_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n372_), .A2(new_n361_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n310_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n368_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n451_), .A2(KEYINPUT20), .A3(new_n452_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(new_n377_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT99), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n450_), .A2(KEYINPUT32), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT99), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n468_), .A2(new_n473_), .A3(new_n377_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n434_), .A2(new_n443_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(new_n453_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n470_), .A2(new_n472_), .A3(new_n474_), .A4(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n458_), .A2(new_n471_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  AOI22_X1  g278(.A1(new_n375_), .A2(new_n463_), .B1(new_n467_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n405_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n439_), .B(new_n398_), .C1(new_n392_), .C2(new_n395_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n404_), .B1(new_n482_), .B2(new_n387_), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT30), .B1(new_n481_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G227gat), .A2(G233gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(G15gat), .ZN(new_n486_));
  XOR2_X1   g285(.A(G71gat), .B(G99gat), .Z(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(KEYINPUT85), .B(G43gat), .Z(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT30), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n403_), .A2(new_n491_), .A3(new_n405_), .ZN(new_n492_));
  AND3_X1   g291(.A1(new_n484_), .A2(new_n490_), .A3(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n490_), .B1(new_n484_), .B2(new_n492_), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT86), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n484_), .A2(new_n492_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n490_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT86), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n484_), .A2(new_n490_), .A3(new_n492_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n498_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n343_), .B(KEYINPUT31), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n495_), .A2(new_n501_), .A3(new_n503_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n498_), .A2(new_n499_), .A3(new_n500_), .A4(new_n502_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  XOR2_X1   g305(.A(G22gat), .B(G50gat), .Z(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G228gat), .A2(G233gat), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT29), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n511_), .B1(new_n349_), .B2(new_n332_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n510_), .B1(new_n437_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n353_), .A2(KEYINPUT29), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n514_), .B(new_n509_), .C1(new_n426_), .C2(new_n433_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G78gat), .B(G106gat), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n513_), .A2(new_n515_), .A3(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n517_), .B1(new_n513_), .B2(new_n515_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n508_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n513_), .A2(new_n515_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(new_n516_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n513_), .A2(new_n515_), .A3(new_n517_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(new_n523_), .A3(new_n507_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n349_), .A2(new_n511_), .A3(new_n332_), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n525_), .B(KEYINPUT28), .Z(new_n526_));
  AND3_X1   g325(.A1(new_n520_), .A2(new_n524_), .A3(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n526_), .B1(new_n520_), .B2(new_n524_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n506_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n480_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n476_), .A2(new_n474_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n473_), .B1(new_n468_), .B2(new_n377_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n449_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT27), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT100), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n534_), .B1(new_n461_), .B2(new_n535_), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n533_), .B(new_n536_), .C1(new_n535_), .C2(new_n461_), .ZN(new_n537_));
  XOR2_X1   g336(.A(KEYINPUT101), .B(KEYINPUT27), .Z(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n539_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n537_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n467_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n504_), .A2(new_n505_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n543_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n526_), .ZN(new_n545_));
  NOR3_X1   g344(.A1(new_n518_), .A2(new_n519_), .A3(new_n508_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n507_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n545_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n520_), .A2(new_n524_), .A3(new_n526_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n548_), .A2(new_n506_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n544_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n541_), .A2(new_n542_), .A3(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n305_), .B1(new_n530_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n244_), .A2(new_n263_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G57gat), .B(G64gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G71gat), .B(G78gat), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n555_), .A2(new_n556_), .A3(KEYINPUT11), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(KEYINPUT11), .ZN(new_n558_));
  INV_X1    g357(.A(new_n556_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n555_), .A2(KEYINPUT11), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n557_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT69), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT69), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n564_), .B(new_n557_), .C1(new_n560_), .C2(new_n561_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(KEYINPUT70), .B1(new_n554_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n279_), .A2(new_n280_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n262_), .B1(new_n568_), .B2(new_n232_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT70), .ZN(new_n570_));
  INV_X1    g369(.A(new_n566_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n569_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n567_), .B(new_n572_), .C1(new_n569_), .C2(new_n571_), .ZN(new_n573_));
  AND2_X1   g372(.A1(G230gat), .A2(G233gat), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT12), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n562_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n282_), .A2(new_n283_), .A3(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n576_), .B1(new_n569_), .B2(new_n571_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n574_), .B1(new_n569_), .B2(new_n571_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G120gat), .B(G148gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT5), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G176gat), .B(G204gat), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n584_), .B(new_n585_), .Z(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n575_), .A2(new_n582_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n587_), .B1(new_n575_), .B2(new_n582_), .ZN(new_n590_));
  OR3_X1    g389(.A1(new_n589_), .A2(KEYINPUT13), .A3(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(KEYINPUT13), .B1(new_n589_), .B2(new_n590_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G15gat), .B(G22gat), .ZN(new_n594_));
  INV_X1    g393(.A(G1gat), .ZN(new_n595_));
  INV_X1    g394(.A(G8gat), .ZN(new_n596_));
  OAI21_X1  g395(.A(KEYINPUT14), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n594_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G1gat), .B(G8gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n273_), .A2(new_n600_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n252_), .A2(new_n600_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G229gat), .A2(G233gat), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n252_), .B(new_n600_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(new_n604_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(G113gat), .B(G141gat), .Z(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT81), .ZN(new_n610_));
  XOR2_X1   g409(.A(G169gat), .B(G197gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n605_), .A2(new_n608_), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n612_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n604_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n615_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n614_), .B1(new_n616_), .B2(new_n607_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n613_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT82), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT82), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n613_), .A2(new_n620_), .A3(new_n617_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n593_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n600_), .B(KEYINPUT78), .ZN(new_n625_));
  NAND2_X1  g424(.A1(G231gat), .A2(G233gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n627_), .A2(new_n562_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT17), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G127gat), .B(G155gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G183gat), .B(G211gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n628_), .A2(new_n629_), .A3(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n627_), .A2(new_n562_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n634_), .B(new_n629_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n638_), .B1(new_n627_), .B2(new_n566_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n639_), .B1(new_n566_), .B2(new_n627_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n637_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n553_), .A2(new_n624_), .A3(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G1gat), .B1(new_n643_), .B2(new_n542_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT37), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n645_), .B1(new_n299_), .B2(new_n304_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n300_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n647_), .B1(new_n289_), .B2(new_n292_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n298_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n302_), .A2(new_n649_), .A3(new_n303_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n648_), .A2(new_n650_), .A3(KEYINPUT37), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n646_), .A2(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n652_), .A2(new_n641_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT80), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n623_), .B1(new_n552_), .B2(new_n530_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n467_), .B(KEYINPUT102), .Z(new_n657_));
  NOR2_X1   g456(.A1(new_n657_), .A2(G1gat), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT103), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n656_), .A2(KEYINPUT103), .A3(new_n658_), .ZN(new_n662_));
  XOR2_X1   g461(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n663_));
  AND3_X1   g462(.A1(new_n661_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n644_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT105), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n668_), .B(new_n644_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(G1324gat));
  OAI21_X1  g469(.A(G8gat), .B1(new_n643_), .B2(new_n541_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT39), .ZN(new_n672_));
  INV_X1    g471(.A(new_n541_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n656_), .A2(new_n596_), .A3(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n675_), .B(new_n676_), .ZN(G1325gat));
  OAI21_X1  g476(.A(G15gat), .B1(new_n643_), .B2(new_n506_), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n678_), .A2(KEYINPUT41), .ZN(new_n679_));
  INV_X1    g478(.A(G15gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n656_), .A2(new_n680_), .A3(new_n543_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n678_), .A2(KEYINPUT41), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n679_), .A2(new_n681_), .A3(new_n682_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT107), .Z(G1326gat));
  NOR2_X1   g483(.A1(new_n527_), .A2(new_n528_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(G22gat), .B1(new_n643_), .B2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT42), .ZN(new_n688_));
  INV_X1    g487(.A(G22gat), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n656_), .A2(new_n689_), .A3(new_n685_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(G1327gat));
  NAND2_X1  g490(.A1(new_n305_), .A2(new_n641_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT110), .Z(new_n693_));
  NAND2_X1  g492(.A1(new_n655_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT111), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n655_), .A2(KEYINPUT111), .A3(new_n693_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G29gat), .B1(new_n698_), .B2(new_n467_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n544_), .A2(new_n550_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n537_), .A2(new_n542_), .A3(new_n540_), .ZN(new_n701_));
  OAI22_X1  g500(.A1(new_n700_), .A2(new_n701_), .B1(new_n480_), .B2(new_n529_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n702_), .A2(new_n703_), .A3(new_n652_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n648_), .A2(KEYINPUT37), .A3(new_n650_), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT37), .B1(new_n648_), .B2(new_n650_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n705_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n646_), .A2(KEYINPUT108), .A3(new_n651_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n703_), .B1(new_n702_), .B2(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n704_), .B1(new_n711_), .B2(KEYINPUT109), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT109), .ZN(new_n713_));
  AOI211_X1 g512(.A(new_n713_), .B(new_n703_), .C1(new_n702_), .C2(new_n710_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n712_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n623_), .A2(new_n642_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n715_), .A2(new_n716_), .A3(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(G29gat), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n719_), .A2(new_n720_), .A3(new_n657_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n716_), .B1(new_n715_), .B2(new_n718_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n699_), .B1(new_n721_), .B2(new_n722_), .ZN(G1328gat));
  AOI22_X1  g522(.A1(new_n530_), .A2(new_n552_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n713_), .B1(new_n724_), .B2(new_n703_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n711_), .A2(KEYINPUT109), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n725_), .A2(new_n726_), .A3(new_n704_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n727_), .A2(KEYINPUT44), .A3(new_n717_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n673_), .ZN(new_n729_));
  AOI21_X1  g528(.A(KEYINPUT44), .B1(new_n727_), .B2(new_n717_), .ZN(new_n730_));
  OAI21_X1  g529(.A(G36gat), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n541_), .A2(G36gat), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n696_), .A2(new_n697_), .A3(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT45), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n731_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT46), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n731_), .A2(KEYINPUT46), .A3(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1329gat));
  AND2_X1   g538(.A1(new_n698_), .A2(new_n543_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n722_), .A2(new_n728_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n543_), .A2(G43gat), .ZN(new_n742_));
  OAI22_X1  g541(.A1(G43gat), .A2(new_n740_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g543(.A(G50gat), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n685_), .A2(new_n745_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT112), .Z(new_n747_));
  NAND2_X1  g546(.A1(new_n698_), .A2(new_n747_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n719_), .A2(new_n730_), .A3(new_n686_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n749_), .B2(new_n745_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT113), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  OAI211_X1 g551(.A(KEYINPUT113), .B(new_n748_), .C1(new_n749_), .C2(new_n745_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(G1331gat));
  NOR2_X1   g553(.A1(new_n593_), .A2(new_n622_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n553_), .A2(new_n642_), .A3(new_n755_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n756_), .A2(new_n308_), .A3(new_n542_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n654_), .A2(new_n702_), .A3(new_n755_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n657_), .B1(new_n758_), .B2(KEYINPUT114), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n759_), .B1(KEYINPUT114), .B2(new_n758_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n757_), .B1(new_n760_), .B2(new_n308_), .ZN(G1332gat));
  OAI21_X1  g560(.A(G64gat), .B1(new_n756_), .B2(new_n541_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT48), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n541_), .A2(G64gat), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT115), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n763_), .B1(new_n758_), .B2(new_n765_), .ZN(G1333gat));
  OAI21_X1  g565(.A(G71gat), .B1(new_n756_), .B2(new_n506_), .ZN(new_n767_));
  XOR2_X1   g566(.A(KEYINPUT116), .B(KEYINPUT49), .Z(new_n768_));
  XNOR2_X1  g567(.A(new_n767_), .B(new_n768_), .ZN(new_n769_));
  OR2_X1    g568(.A1(new_n506_), .A2(G71gat), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(new_n758_), .B2(new_n770_), .ZN(G1334gat));
  OAI21_X1  g570(.A(G78gat), .B1(new_n756_), .B2(new_n686_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT50), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n686_), .A2(G78gat), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT117), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n773_), .B1(new_n758_), .B2(new_n775_), .ZN(G1335gat));
  INV_X1    g575(.A(G85gat), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n593_), .A2(new_n622_), .A3(new_n642_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n727_), .A2(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n777_), .B1(new_n779_), .B2(new_n467_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n693_), .A2(new_n702_), .A3(new_n755_), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n781_), .A2(G85gat), .A3(new_n657_), .ZN(new_n782_));
  OR2_X1    g581(.A1(new_n780_), .A2(new_n782_), .ZN(G1336gat));
  NOR3_X1   g582(.A1(new_n781_), .A2(G92gat), .A3(new_n541_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n779_), .A2(new_n673_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n785_), .B2(G92gat), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT118), .ZN(G1337gat));
  NAND2_X1  g586(.A1(KEYINPUT119), .A2(KEYINPUT51), .ZN(new_n788_));
  OR2_X1    g587(.A1(new_n506_), .A2(new_n260_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n788_), .B1(new_n781_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n779_), .A2(new_n543_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(G99gat), .ZN(new_n792_));
  NOR2_X1   g591(.A1(KEYINPUT119), .A2(KEYINPUT51), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n792_), .B(new_n793_), .ZN(G1338gat));
  OR3_X1    g593(.A1(new_n781_), .A2(G106gat), .A3(new_n686_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n685_), .B(new_n778_), .C1(new_n712_), .C2(new_n714_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n797_), .A3(G106gat), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n797_), .B1(new_n796_), .B2(G106gat), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(KEYINPUT120), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT120), .ZN(new_n801_));
  AOI211_X1 g600(.A(new_n801_), .B(new_n797_), .C1(new_n796_), .C2(G106gat), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n795_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT53), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n805_), .B(new_n795_), .C1(new_n800_), .C2(new_n802_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(G1339gat));
  NOR3_X1   g606(.A1(new_n673_), .A2(new_n657_), .A3(new_n544_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n614_), .B1(new_n606_), .B2(new_n604_), .ZN(new_n809_));
  XOR2_X1   g608(.A(new_n603_), .B(KEYINPUT122), .Z(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(new_n604_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n617_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n812_), .A2(new_n589_), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n579_), .A2(new_n567_), .A3(new_n580_), .A4(new_n572_), .ZN(new_n815_));
  AOI22_X1  g614(.A1(new_n814_), .A2(KEYINPUT55), .B1(new_n815_), .B2(new_n574_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT121), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n817_), .B1(new_n582_), .B2(new_n818_), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n582_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n816_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n821_), .A2(KEYINPUT56), .A3(new_n586_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT56), .B1(new_n821_), .B2(new_n586_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n823_), .B2(KEYINPUT123), .ZN(new_n824_));
  OAI21_X1  g623(.A(KEYINPUT121), .B1(new_n814_), .B2(KEYINPUT55), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n582_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n587_), .B1(new_n827_), .B2(new_n816_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT123), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n828_), .A2(new_n829_), .A3(KEYINPUT56), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n813_), .B1(new_n824_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n833_), .A2(KEYINPUT124), .A3(new_n652_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT124), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n829_), .B1(new_n828_), .B2(KEYINPUT56), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n821_), .A2(new_n586_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT56), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(KEYINPUT123), .A3(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n836_), .A2(new_n839_), .A3(new_n822_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT58), .B1(new_n840_), .B2(new_n813_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n652_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n835_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n831_), .A2(new_n832_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n834_), .A2(new_n843_), .A3(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n305_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n622_), .A2(new_n588_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n823_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(new_n822_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n589_), .A2(new_n590_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n812_), .A2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n847_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n822_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n622_), .B(new_n588_), .C1(new_n856_), .C2(new_n823_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n852_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n859_), .A2(KEYINPUT57), .A3(new_n847_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n855_), .A2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n642_), .B1(new_n846_), .B2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n622_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n653_), .A2(new_n863_), .A3(new_n593_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(KEYINPUT54), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n808_), .B1(new_n862_), .B2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT125), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n855_), .A2(new_n860_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n842_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n844_), .B1(new_n870_), .B2(KEYINPUT124), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n869_), .B1(new_n871_), .B2(new_n843_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n865_), .B1(new_n872_), .B2(new_n642_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT125), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n873_), .A2(new_n874_), .A3(new_n808_), .ZN(new_n875_));
  INV_X1    g674(.A(G113gat), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n868_), .A2(new_n875_), .A3(new_n876_), .A4(new_n622_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n867_), .A2(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n873_), .A2(KEYINPUT59), .A3(new_n808_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n863_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n877_), .B1(new_n881_), .B2(new_n876_), .ZN(G1340gat));
  INV_X1    g681(.A(new_n593_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT60), .ZN(new_n884_));
  INV_X1    g683(.A(G120gat), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n883_), .A2(new_n884_), .A3(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n886_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n868_), .A2(new_n875_), .A3(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n593_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(new_n885_), .ZN(G1341gat));
  INV_X1    g689(.A(G127gat), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n868_), .A2(new_n875_), .A3(new_n891_), .A4(new_n642_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n641_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n891_), .ZN(G1342gat));
  INV_X1    g693(.A(G134gat), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n868_), .A2(new_n875_), .A3(new_n895_), .A4(new_n305_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n842_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n897_), .B2(new_n895_), .ZN(G1343gat));
  INV_X1    g697(.A(new_n550_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n673_), .A2(new_n657_), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n873_), .A2(new_n899_), .A3(new_n622_), .A4(new_n900_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT126), .B(G141gat), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1344gat));
  NAND3_X1  g702(.A1(new_n873_), .A2(new_n899_), .A3(new_n900_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n905_), .A2(new_n321_), .A3(new_n883_), .ZN(new_n906_));
  OAI21_X1  g705(.A(G148gat), .B1(new_n904_), .B2(new_n593_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(G1345gat));
  NAND4_X1  g707(.A1(new_n873_), .A2(new_n899_), .A3(new_n642_), .A4(new_n900_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(KEYINPUT61), .B(G155gat), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n909_), .B(new_n910_), .ZN(G1346gat));
  AOI21_X1  g710(.A(new_n313_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n873_), .A2(new_n305_), .A3(new_n899_), .A4(new_n900_), .ZN(new_n913_));
  AOI22_X1  g712(.A1(new_n905_), .A2(new_n912_), .B1(new_n913_), .B2(new_n313_), .ZN(G1347gat));
  NAND3_X1  g713(.A1(new_n657_), .A2(new_n543_), .A3(new_n686_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(new_n541_), .ZN(new_n916_));
  OAI211_X1 g715(.A(new_n622_), .B(new_n916_), .C1(new_n862_), .C2(new_n866_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(G169gat), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n917_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n921_));
  INV_X1    g720(.A(new_n378_), .ZN(new_n922_));
  OAI211_X1 g721(.A(new_n920_), .B(new_n921_), .C1(new_n922_), .C2(new_n917_), .ZN(G1348gat));
  NAND3_X1  g722(.A1(new_n873_), .A2(new_n883_), .A3(new_n916_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(G176gat), .ZN(G1349gat));
  NOR2_X1   g724(.A1(new_n862_), .A2(new_n866_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n916_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n642_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(G183gat), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n928_), .A2(new_n388_), .A3(new_n642_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1350gat));
  NAND2_X1  g731(.A1(new_n928_), .A2(new_n652_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(G190gat), .ZN(new_n934_));
  NAND4_X1  g733(.A1(new_n928_), .A2(new_n305_), .A3(new_n390_), .A4(new_n394_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(G1351gat));
  NOR2_X1   g735(.A1(new_n541_), .A2(new_n467_), .ZN(new_n937_));
  NAND4_X1  g736(.A1(new_n873_), .A2(new_n899_), .A3(new_n622_), .A4(new_n937_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n593_), .B1(new_n940_), .B2(G204gat), .ZN(new_n941_));
  NAND4_X1  g740(.A1(new_n873_), .A2(new_n899_), .A3(new_n937_), .A4(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n411_), .A2(KEYINPUT127), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n942_), .B(new_n943_), .ZN(G1353gat));
  NAND3_X1  g743(.A1(new_n873_), .A2(new_n899_), .A3(new_n937_), .ZN(new_n945_));
  XOR2_X1   g744(.A(KEYINPUT63), .B(G211gat), .Z(new_n946_));
  OR3_X1    g745(.A1(new_n945_), .A2(new_n641_), .A3(new_n946_), .ZN(new_n947_));
  OAI22_X1  g746(.A1(new_n945_), .A2(new_n641_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(new_n948_), .ZN(G1354gat));
  OAI21_X1  g748(.A(G218gat), .B1(new_n945_), .B2(new_n842_), .ZN(new_n950_));
  OR2_X1    g749(.A1(new_n847_), .A2(G218gat), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n950_), .B1(new_n945_), .B2(new_n951_), .ZN(G1355gat));
endmodule


