//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 0 1 0 1 0 0 1 1 0 1 1 0 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n923_,
    new_n924_, new_n925_, new_n927_, new_n928_, new_n930_, new_n931_,
    new_n932_, new_n934_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_;
  INV_X1    g000(.A(KEYINPUT107), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G226gat), .A2(G233gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT25), .B(G183gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT26), .B(G190gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G169gat), .ZN(new_n215_));
  INV_X1    g014(.A(G176gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(KEYINPUT24), .A3(new_n218_), .ZN(new_n219_));
  OR3_X1    g018(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n209_), .A2(new_n214_), .A3(new_n219_), .A4(new_n220_), .ZN(new_n221_));
  OR2_X1    g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n212_), .A2(new_n222_), .A3(new_n213_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT22), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n224_), .B1(KEYINPUT83), .B2(G169gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(KEYINPUT83), .A3(G169gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(new_n216_), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n223_), .B(new_n218_), .C1(new_n225_), .C2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n221_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G197gat), .B(G204gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G211gat), .B(G218gat), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT89), .ZN(new_n232_));
  OAI211_X1 g031(.A(KEYINPUT21), .B(new_n230_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT21), .ZN(new_n234_));
  XOR2_X1   g033(.A(G211gat), .B(G218gat), .Z(new_n235_));
  AOI21_X1  g034(.A(new_n234_), .B1(new_n235_), .B2(KEYINPUT89), .ZN(new_n236_));
  XOR2_X1   g035(.A(G197gat), .B(G204gat), .Z(new_n237_));
  OAI21_X1  g036(.A(new_n237_), .B1(KEYINPUT21), .B2(new_n231_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n233_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT20), .B1(new_n229_), .B2(new_n239_), .ZN(new_n240_));
  AND4_X1   g039(.A1(new_n219_), .A2(new_n220_), .A3(new_n212_), .A4(new_n213_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n207_), .A2(KEYINPUT94), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT94), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT25), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n244_), .A2(G183gat), .ZN(new_n245_));
  INV_X1    g044(.A(G183gat), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n246_), .A2(KEYINPUT25), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n243_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n242_), .A2(new_n248_), .A3(new_n208_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n241_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT95), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n223_), .A2(new_n251_), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n212_), .A2(new_n222_), .A3(KEYINPUT95), .A4(new_n213_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT22), .B(G169gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(new_n216_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n252_), .A2(new_n218_), .A3(new_n253_), .A4(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n235_), .A2(new_n234_), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT21), .B1(new_n231_), .B2(new_n232_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(new_n258_), .A3(new_n237_), .ZN(new_n259_));
  AOI22_X1  g058(.A1(new_n250_), .A2(new_n256_), .B1(new_n259_), .B2(new_n233_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n206_), .B1(new_n240_), .B2(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(G8gat), .B(G36gat), .Z(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT18), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G64gat), .B(G92gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT20), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n266_), .B1(new_n229_), .B2(new_n239_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n250_), .A2(new_n256_), .A3(new_n259_), .A4(new_n233_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(new_n205_), .A3(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n261_), .A2(new_n265_), .A3(new_n269_), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n270_), .A2(KEYINPUT103), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(KEYINPUT103), .ZN(new_n272_));
  INV_X1    g071(.A(new_n265_), .ZN(new_n273_));
  NOR3_X1   g072(.A1(new_n240_), .A2(new_n260_), .A3(new_n206_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n205_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n273_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n271_), .A2(KEYINPUT27), .A3(new_n272_), .A4(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n261_), .A2(new_n269_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n273_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n280_), .A2(KEYINPUT96), .A3(new_n270_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT27), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT96), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n261_), .A2(new_n283_), .A3(new_n269_), .A4(new_n265_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n281_), .A2(new_n282_), .A3(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT104), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT104), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n281_), .A2(new_n287_), .A3(new_n282_), .A4(new_n284_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n278_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n239_), .A2(KEYINPUT90), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G228gat), .A2(G233gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  XOR2_X1   g092(.A(G141gat), .B(G148gat), .Z(new_n294_));
  INV_X1    g093(.A(G155gat), .ZN(new_n295_));
  INV_X1    g094(.A(G162gat), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n295_), .A2(new_n296_), .A3(KEYINPUT86), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT86), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n298_), .B1(G155gat), .B2(G162gat), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT1), .B1(new_n295_), .B2(new_n296_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT1), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n302_), .A2(G155gat), .A3(G162gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n294_), .B1(new_n300_), .B2(new_n304_), .ZN(new_n305_));
  AOI22_X1  g104(.A1(new_n297_), .A2(new_n299_), .B1(G155gat), .B2(G162gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G141gat), .A2(G148gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT87), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT2), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT3), .ZN(new_n311_));
  INV_X1    g110(.A(G141gat), .ZN(new_n312_));
  INV_X1    g111(.A(G148gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n311_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n310_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n309_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n306_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n305_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT29), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(new_n239_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n293_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G78gat), .B(G106gat), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n290_), .A2(new_n320_), .A3(new_n239_), .A4(new_n292_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n322_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n323_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT88), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n305_), .A2(new_n318_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT29), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n329_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NOR3_X1   g131(.A1(new_n319_), .A2(KEYINPUT88), .A3(KEYINPUT29), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT28), .B(G22gat), .ZN(new_n334_));
  INV_X1    g133(.A(G50gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NOR3_X1   g136(.A1(new_n332_), .A2(new_n333_), .A3(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n330_), .A2(new_n329_), .A3(new_n331_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT88), .B1(new_n319_), .B2(KEYINPUT29), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n336_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT91), .B1(new_n338_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT92), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n337_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT91), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n339_), .A2(new_n336_), .A3(new_n340_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n344_), .A2(new_n346_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT92), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(KEYINPUT91), .A3(new_n349_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n328_), .A2(new_n343_), .A3(new_n347_), .A4(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n322_), .A2(new_n324_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n323_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n354_), .A2(new_n347_), .A3(new_n325_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n349_), .B1(new_n348_), .B2(KEYINPUT91), .ZN(new_n356_));
  AOI211_X1 g155(.A(new_n345_), .B(KEYINPUT92), .C1(new_n344_), .C2(new_n346_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n355_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n351_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G227gat), .A2(G233gat), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n360_), .B(G71gat), .Z(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G15gat), .B(G43gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT84), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT30), .ZN(new_n365_));
  OR2_X1    g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n364_), .A2(new_n365_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(new_n229_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n229_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n362_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(G134gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(G127gat), .ZN(new_n375_));
  INV_X1    g174(.A(G127gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(G134gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(G120gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(G113gat), .ZN(new_n380_));
  INV_X1    g179(.A(G113gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(G120gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(KEYINPUT85), .B1(new_n378_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n378_), .A2(new_n383_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n375_), .A2(new_n377_), .A3(new_n380_), .A4(new_n382_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n384_), .B1(new_n387_), .B2(KEYINPUT85), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT31), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(G99gat), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n369_), .A2(new_n371_), .A3(new_n362_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n388_), .B(KEYINPUT31), .ZN(new_n393_));
  INV_X1    g192(.A(G99gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n373_), .A2(new_n391_), .A3(new_n392_), .A4(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n391_), .A2(new_n395_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n392_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n397_), .B1(new_n398_), .B2(new_n372_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n396_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G1gat), .B(G29gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(G85gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT0), .B(G57gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G225gat), .A2(G233gat), .ZN(new_n405_));
  XOR2_X1   g204(.A(new_n405_), .B(KEYINPUT99), .Z(new_n406_));
  NAND2_X1  g205(.A1(new_n388_), .A2(new_n319_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n406_), .B1(new_n407_), .B2(KEYINPUT4), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT97), .ZN(new_n409_));
  AND4_X1   g208(.A1(new_n375_), .A2(new_n377_), .A3(new_n380_), .A4(new_n382_), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n375_), .A2(new_n377_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n409_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n385_), .A2(KEYINPUT97), .A3(new_n386_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n412_), .A2(new_n318_), .A3(new_n305_), .A4(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n407_), .A2(KEYINPUT4), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT98), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT98), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n407_), .A2(new_n417_), .A3(new_n414_), .A4(KEYINPUT4), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n408_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n406_), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n407_), .A2(new_n420_), .A3(new_n414_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n404_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n416_), .A2(new_n418_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n408_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n421_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n404_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n400_), .A2(new_n422_), .A3(new_n427_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n359_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT106), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n289_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n430_), .B1(new_n289_), .B2(new_n429_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT33), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n434_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n435_));
  NOR4_X1   g234(.A1(new_n419_), .A2(KEYINPUT33), .A3(new_n421_), .A4(new_n404_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n407_), .A2(new_n406_), .A3(new_n414_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n404_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT100), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n407_), .A2(KEYINPUT4), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n423_), .A2(new_n420_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n261_), .A2(new_n265_), .A3(new_n269_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n265_), .B1(new_n261_), .B2(new_n269_), .ZN(new_n445_));
  NOR3_X1   g244(.A1(new_n444_), .A2(new_n445_), .A3(new_n283_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n284_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n443_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT101), .B1(new_n437_), .B2(new_n448_), .ZN(new_n449_));
  AOI22_X1  g248(.A1(new_n281_), .A2(new_n284_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT101), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n450_), .B(new_n451_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n427_), .A2(new_n422_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n279_), .B1(KEYINPUT32), .B2(new_n265_), .ZN(new_n454_));
  OAI211_X1 g253(.A(KEYINPUT32), .B(new_n265_), .C1(new_n274_), .C2(new_n275_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n454_), .B1(KEYINPUT102), .B2(new_n455_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n453_), .B(new_n456_), .C1(KEYINPUT102), .C2(new_n455_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n449_), .A2(new_n452_), .A3(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n359_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n453_), .B1(new_n351_), .B2(new_n358_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n289_), .A2(KEYINPUT105), .A3(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n286_), .A2(new_n288_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(new_n461_), .A3(new_n277_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT105), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n460_), .A2(new_n462_), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n400_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n433_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(G29gat), .B(G36gat), .Z(new_n470_));
  XOR2_X1   g269(.A(G43gat), .B(G50gat), .Z(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(KEYINPUT75), .B(KEYINPUT15), .Z(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G1gat), .B(G8gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT78), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G15gat), .B(G22gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G1gat), .A2(G8gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT14), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n476_), .A2(new_n480_), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n475_), .A2(KEYINPUT78), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n475_), .A2(KEYINPUT78), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n482_), .A2(new_n479_), .A3(new_n477_), .A4(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n481_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n474_), .A2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n481_), .A2(new_n472_), .A3(new_n484_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G229gat), .A2(G233gat), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT80), .ZN(new_n490_));
  INV_X1    g289(.A(new_n472_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n485_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(new_n487_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n488_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n490_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  AOI211_X1 g294(.A(KEYINPUT80), .B(new_n488_), .C1(new_n492_), .C2(new_n487_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n489_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G113gat), .B(G141gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT81), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G169gat), .B(G197gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n497_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n501_), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n489_), .B(new_n503_), .C1(new_n495_), .C2(new_n496_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT82), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n202_), .B1(new_n469_), .B2(new_n508_), .ZN(new_n509_));
  AOI22_X1  g308(.A1(new_n458_), .A2(new_n459_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n400_), .B1(new_n510_), .B2(new_n462_), .ZN(new_n511_));
  OAI211_X1 g310(.A(KEYINPUT107), .B(new_n507_), .C1(new_n511_), .C2(new_n433_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n509_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT74), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT71), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT67), .B(G71gat), .ZN(new_n516_));
  INV_X1    g315(.A(G78gat), .ZN(new_n517_));
  OR2_X1    g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(G57gat), .B(G64gat), .Z(new_n519_));
  INV_X1    g318(.A(KEYINPUT11), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n516_), .A2(new_n517_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n518_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT68), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT68), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n518_), .A2(new_n521_), .A3(new_n525_), .A4(new_n522_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n519_), .A2(new_n520_), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n524_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n527_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n515_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n524_), .A2(new_n526_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n527_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n524_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(KEYINPUT71), .A3(new_n534_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n530_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT72), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT69), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT8), .ZN(new_n539_));
  XOR2_X1   g338(.A(G85gat), .B(G92gat), .Z(new_n540_));
  NOR2_X1   g339(.A1(G99gat), .A2(G106gat), .ZN(new_n541_));
  NOR2_X1   g340(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G99gat), .A2(G106gat), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT6), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n539_), .B(new_n540_), .C1(new_n543_), .C2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n540_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT66), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n544_), .B(KEYINPUT6), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n543_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n546_), .A2(KEYINPUT66), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n548_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n538_), .B(new_n547_), .C1(new_n553_), .C2(new_n539_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n550_), .A2(new_n549_), .ZN(new_n555_));
  INV_X1    g354(.A(G106gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n394_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(new_n542_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n552_), .A2(new_n555_), .A3(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n539_), .B1(new_n559_), .B2(new_n540_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n547_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT69), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(KEYINPUT10), .B(G99gat), .Z(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(new_n556_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n540_), .A2(KEYINPUT9), .ZN(new_n565_));
  INV_X1    g364(.A(G85gat), .ZN(new_n566_));
  INV_X1    g365(.A(G92gat), .ZN(new_n567_));
  OR3_X1    g366(.A1(new_n566_), .A2(new_n567_), .A3(KEYINPUT9), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n564_), .A2(new_n565_), .A3(new_n550_), .A4(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT70), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n554_), .A2(new_n562_), .A3(new_n570_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n536_), .A2(new_n537_), .A3(KEYINPUT12), .A4(new_n571_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n571_), .A2(new_n530_), .A3(new_n535_), .A4(KEYINPUT12), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT72), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G230gat), .A2(G233gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT64), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n547_), .B1(new_n553_), .B2(new_n539_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(new_n569_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n533_), .A2(new_n534_), .ZN(new_n579_));
  OAI21_X1  g378(.A(KEYINPUT12), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n579_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n572_), .A2(new_n574_), .A3(new_n576_), .A4(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n576_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n581_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n578_), .A2(new_n579_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n584_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(G120gat), .B(G148gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G176gat), .B(G204gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n583_), .A2(new_n587_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n593_), .B1(new_n583_), .B2(new_n587_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n514_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n596_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n598_), .A2(KEYINPUT74), .A3(new_n594_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT13), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(KEYINPUT13), .B1(new_n597_), .B2(new_n599_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G231gat), .A2(G233gat), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n485_), .B(new_n605_), .Z(new_n606_));
  AND2_X1   g405(.A1(new_n536_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT17), .ZN(new_n608_));
  XOR2_X1   g407(.A(G127gat), .B(G155gat), .Z(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT16), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G183gat), .B(G211gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n607_), .A2(new_n608_), .A3(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n613_), .B1(new_n536_), .B2(new_n606_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n606_), .B(KEYINPUT79), .ZN(new_n615_));
  INV_X1    g414(.A(new_n579_), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n616_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n612_), .B(KEYINPUT17), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n617_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n614_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n578_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT35), .ZN(new_n623_));
  NAND2_X1  g422(.A1(G232gat), .A2(G233gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT34), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  AOI22_X1  g425(.A1(new_n622_), .A2(new_n472_), .B1(new_n623_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT76), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n571_), .A2(new_n628_), .A3(new_n474_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n628_), .B1(new_n571_), .B2(new_n474_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n627_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n626_), .A2(new_n623_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  XOR2_X1   g432(.A(G190gat), .B(G218gat), .Z(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT77), .ZN(new_n635_));
  XOR2_X1   g434(.A(G134gat), .B(G162gat), .Z(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n638_), .A2(KEYINPUT36), .ZN(new_n639_));
  OAI221_X1 g438(.A(new_n627_), .B1(new_n623_), .B2(new_n626_), .C1(new_n629_), .C2(new_n630_), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n633_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n637_), .B(KEYINPUT36), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n643_), .B1(new_n633_), .B2(new_n640_), .ZN(new_n644_));
  OAI21_X1  g443(.A(KEYINPUT37), .B1(new_n641_), .B2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n633_), .A2(new_n640_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(new_n642_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT37), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n633_), .A2(new_n640_), .A3(new_n639_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n647_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n645_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n604_), .A2(new_n621_), .A3(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n513_), .A2(new_n653_), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n654_), .A2(KEYINPUT108), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(KEYINPUT108), .ZN(new_n656_));
  INV_X1    g455(.A(new_n453_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n657_), .A2(G1gat), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n655_), .A2(new_n656_), .A3(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT38), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n641_), .A2(new_n644_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n469_), .A2(new_n621_), .A3(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n604_), .A2(new_n508_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G1gat), .B1(new_n665_), .B2(new_n657_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n659_), .A2(new_n660_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n661_), .A2(new_n666_), .A3(new_n667_), .ZN(G1324gat));
  OAI21_X1  g467(.A(G8gat), .B1(new_n665_), .B2(new_n289_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT39), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n289_), .A2(G8gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n655_), .A2(new_n656_), .A3(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT40), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n670_), .A2(KEYINPUT40), .A3(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1325gat));
  OAI21_X1  g476(.A(G15gat), .B1(new_n665_), .B2(new_n468_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT41), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n654_), .A2(G15gat), .A3(new_n468_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1326gat));
  OAI21_X1  g480(.A(G22gat), .B1(new_n665_), .B2(new_n459_), .ZN(new_n682_));
  XOR2_X1   g481(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n683_));
  XNOR2_X1  g482(.A(new_n682_), .B(new_n683_), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n459_), .A2(G22gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n684_), .B1(new_n654_), .B2(new_n685_), .ZN(G1327gat));
  INV_X1    g485(.A(new_n662_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n621_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n689_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT111), .B1(new_n513_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT111), .ZN(new_n693_));
  AOI211_X1 g492(.A(new_n693_), .B(new_n690_), .C1(new_n509_), .C2(new_n512_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n692_), .A2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G29gat), .B1(new_n695_), .B2(new_n453_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n467_), .A2(new_n468_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n433_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT110), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n651_), .B(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n651_), .A2(KEYINPUT43), .ZN(new_n704_));
  AOI22_X1  g503(.A1(new_n703_), .A2(KEYINPUT43), .B1(new_n700_), .B2(new_n704_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n604_), .A2(new_n508_), .A3(new_n688_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n697_), .B1(new_n705_), .B2(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n651_), .B(KEYINPUT110), .ZN(new_n709_));
  OAI21_X1  g508(.A(KEYINPUT43), .B1(new_n709_), .B2(new_n469_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n700_), .A2(new_n704_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n712_), .A2(KEYINPUT44), .A3(new_n706_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n708_), .A2(new_n713_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n453_), .A2(G29gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n696_), .B1(new_n714_), .B2(new_n715_), .ZN(G1328gat));
  INV_X1    g515(.A(new_n289_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n708_), .A2(new_n717_), .A3(new_n713_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(G36gat), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT45), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n289_), .A2(G36gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n695_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n721_), .ZN(new_n723_));
  NOR4_X1   g522(.A1(new_n692_), .A2(new_n694_), .A3(KEYINPUT45), .A4(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n719_), .B1(new_n722_), .B2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(KEYINPUT112), .B(KEYINPUT46), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n719_), .B(new_n726_), .C1(new_n722_), .C2(new_n724_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1329gat));
  XNOR2_X1  g529(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n731_));
  INV_X1    g530(.A(G43gat), .ZN(new_n732_));
  INV_X1    g531(.A(new_n695_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(new_n468_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n708_), .A2(G43gat), .A3(new_n400_), .A4(new_n713_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n731_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n692_), .A2(new_n694_), .A3(new_n468_), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n735_), .B(new_n731_), .C1(new_n737_), .C2(G43gat), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n736_), .A2(new_n739_), .ZN(G1330gat));
  NAND3_X1  g539(.A1(new_n695_), .A2(new_n335_), .A3(new_n359_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT114), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n714_), .A2(new_n742_), .A3(new_n359_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(G50gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n742_), .B1(new_n714_), .B2(new_n359_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n741_), .B1(new_n744_), .B2(new_n745_), .ZN(G1331gat));
  INV_X1    g545(.A(G57gat), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n602_), .A2(new_n603_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n748_), .A2(new_n507_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(new_n663_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT115), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n747_), .B1(new_n751_), .B2(new_n453_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n748_), .A2(new_n507_), .A3(new_n469_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n621_), .B1(new_n645_), .B2(new_n650_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n755_), .A2(new_n747_), .A3(new_n453_), .ZN(new_n756_));
  OR2_X1    g555(.A1(new_n752_), .A2(new_n756_), .ZN(G1332gat));
  INV_X1    g556(.A(G64gat), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n755_), .A2(new_n758_), .A3(new_n717_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT48), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n751_), .A2(new_n717_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(G64gat), .ZN(new_n762_));
  AOI211_X1 g561(.A(KEYINPUT48), .B(new_n758_), .C1(new_n751_), .C2(new_n717_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n759_), .B1(new_n762_), .B2(new_n763_), .ZN(G1333gat));
  NOR2_X1   g563(.A1(new_n468_), .A2(G71gat), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT116), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n755_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n751_), .A2(new_n400_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT49), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n768_), .A2(new_n769_), .A3(G71gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n768_), .B2(G71gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n770_), .B2(new_n771_), .ZN(G1334gat));
  NAND3_X1  g571(.A1(new_n755_), .A2(new_n517_), .A3(new_n359_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n751_), .A2(new_n359_), .ZN(new_n774_));
  XOR2_X1   g573(.A(KEYINPUT117), .B(KEYINPUT50), .Z(new_n775_));
  AND3_X1   g574(.A1(new_n774_), .A2(G78gat), .A3(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n774_), .B2(G78gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(G1335gat));
  NAND3_X1  g577(.A1(new_n712_), .A2(new_n621_), .A3(new_n749_), .ZN(new_n779_));
  OAI21_X1  g578(.A(G85gat), .B1(new_n779_), .B2(new_n657_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n753_), .A2(new_n689_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n782_), .A2(new_n566_), .A3(new_n453_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n780_), .A2(new_n783_), .ZN(G1336gat));
  OAI21_X1  g583(.A(G92gat), .B1(new_n779_), .B2(new_n289_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n782_), .A2(new_n567_), .A3(new_n717_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(G1337gat));
  OAI21_X1  g586(.A(G99gat), .B1(new_n779_), .B2(new_n468_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n400_), .A2(new_n563_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n788_), .B1(new_n781_), .B2(new_n789_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g590(.A1(new_n782_), .A2(new_n556_), .A3(new_n359_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n712_), .A2(new_n359_), .A3(new_n621_), .A4(new_n749_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n793_), .A2(new_n794_), .A3(G106gat), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n793_), .B2(G106gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n792_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g597(.A(KEYINPUT59), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n507_), .A2(new_n594_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n583_), .A2(new_n801_), .ZN(new_n802_));
  AOI22_X1  g601(.A1(new_n573_), .A2(KEYINPUT72), .B1(new_n580_), .B2(new_n581_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n572_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n584_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n803_), .A2(new_n572_), .A3(KEYINPUT55), .A4(new_n576_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n802_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n592_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT56), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n807_), .A2(KEYINPUT56), .A3(new_n592_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n800_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT119), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n486_), .A2(new_n487_), .A3(new_n494_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n494_), .B1(new_n492_), .B2(new_n487_), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT118), .B1(new_n815_), .B2(new_n503_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n815_), .A2(KEYINPUT118), .A3(new_n503_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n813_), .B(new_n814_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n504_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n818_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n816_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n813_), .B1(new_n822_), .B2(new_n814_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n820_), .A2(new_n823_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n597_), .A2(new_n599_), .A3(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n687_), .B1(new_n812_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n824_), .A2(new_n594_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT120), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT120), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n824_), .A2(new_n831_), .A3(new_n594_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n811_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT56), .B1(new_n807_), .B2(new_n592_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n833_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT58), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT121), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n836_), .A2(new_n839_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n833_), .B(new_n838_), .C1(new_n834_), .C2(new_n835_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n841_), .A3(new_n652_), .ZN(new_n842_));
  OAI211_X1 g641(.A(KEYINPUT57), .B(new_n687_), .C1(new_n812_), .C2(new_n825_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n828_), .A2(new_n842_), .A3(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n748_), .A2(new_n845_), .A3(new_n508_), .A4(new_n754_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n508_), .B(new_n754_), .C1(new_n602_), .C2(new_n603_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT54), .ZN(new_n848_));
  AOI22_X1  g647(.A1(new_n844_), .A2(new_n621_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n849_));
  NOR4_X1   g648(.A1(new_n717_), .A2(new_n468_), .A3(new_n657_), .A4(new_n359_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n799_), .B1(new_n849_), .B2(new_n851_), .ZN(new_n852_));
  AOI22_X1  g651(.A1(new_n810_), .A2(new_n811_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n651_), .B1(new_n853_), .B2(new_n838_), .ZN(new_n854_));
  AOI22_X1  g653(.A1(new_n840_), .A2(new_n854_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n688_), .B1(new_n855_), .B2(new_n843_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n846_), .A2(new_n848_), .ZN(new_n857_));
  OAI211_X1 g656(.A(KEYINPUT59), .B(new_n850_), .C1(new_n856_), .C2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n852_), .A2(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n508_), .A2(new_n381_), .ZN(new_n860_));
  XOR2_X1   g659(.A(new_n860_), .B(KEYINPUT122), .Z(new_n861_));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n844_), .A2(new_n621_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n846_), .A2(new_n848_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n850_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n381_), .B1(new_n866_), .B2(new_n508_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n862_), .A2(KEYINPUT123), .A3(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT123), .ZN(new_n869_));
  INV_X1    g668(.A(new_n861_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(new_n852_), .B2(new_n858_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n849_), .A2(new_n851_), .ZN(new_n872_));
  AOI21_X1  g671(.A(G113gat), .B1(new_n872_), .B2(new_n507_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n869_), .B1(new_n871_), .B2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n868_), .A2(new_n874_), .ZN(G1340gat));
  OAI21_X1  g674(.A(new_n379_), .B1(new_n748_), .B2(KEYINPUT60), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n872_), .B(new_n876_), .C1(KEYINPUT60), .C2(new_n379_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n748_), .B1(new_n852_), .B2(new_n858_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n878_), .B2(new_n379_), .ZN(G1341gat));
  OAI21_X1  g678(.A(new_n376_), .B1(new_n866_), .B2(new_n621_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  OAI211_X1 g681(.A(KEYINPUT124), .B(new_n376_), .C1(new_n866_), .C2(new_n621_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n688_), .A2(G127gat), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n882_), .A2(new_n883_), .B1(new_n859_), .B2(new_n885_), .ZN(G1342gat));
  NAND3_X1  g685(.A1(new_n872_), .A2(new_n374_), .A3(new_n662_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n651_), .B1(new_n852_), .B2(new_n858_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n888_), .B2(new_n374_), .ZN(G1343gat));
  NOR4_X1   g688(.A1(new_n717_), .A2(new_n400_), .A3(new_n657_), .A4(new_n459_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n849_), .A2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n507_), .ZN(new_n893_));
  XOR2_X1   g692(.A(KEYINPUT125), .B(G141gat), .Z(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1344gat));
  NAND2_X1  g694(.A1(new_n892_), .A2(new_n604_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g696(.A1(new_n865_), .A2(new_n688_), .A3(new_n890_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(KEYINPUT126), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT126), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n892_), .A2(new_n900_), .A3(new_n688_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT61), .B(G155gat), .ZN(new_n902_));
  AND3_X1   g701(.A1(new_n899_), .A2(new_n901_), .A3(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n902_), .B1(new_n899_), .B2(new_n901_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1346gat));
  AOI21_X1  g704(.A(G162gat), .B1(new_n892_), .B2(new_n662_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n709_), .A2(new_n296_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n892_), .B2(new_n907_), .ZN(G1347gat));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n289_), .A2(new_n359_), .A3(new_n428_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n865_), .A2(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(new_n508_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n909_), .B1(new_n912_), .B2(new_n215_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n254_), .ZN(new_n914_));
  OAI211_X1 g713(.A(KEYINPUT62), .B(G169gat), .C1(new_n911_), .C2(new_n508_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n913_), .A2(new_n914_), .A3(new_n915_), .ZN(G1348gat));
  NOR2_X1   g715(.A1(KEYINPUT127), .A2(G176gat), .ZN(new_n917_));
  NOR3_X1   g716(.A1(new_n911_), .A2(new_n748_), .A3(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n911_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(new_n604_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(KEYINPUT127), .B(G176gat), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n918_), .B1(new_n920_), .B2(new_n921_), .ZN(G1349gat));
  AND2_X1   g721(.A1(new_n242_), .A2(new_n248_), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n911_), .A2(new_n923_), .A3(new_n621_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n919_), .A2(new_n688_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n924_), .B1(new_n246_), .B2(new_n925_), .ZN(G1350gat));
  OAI21_X1  g725(.A(G190gat), .B1(new_n911_), .B2(new_n651_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n662_), .A2(new_n208_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n927_), .B1(new_n911_), .B2(new_n928_), .ZN(G1351gat));
  NAND3_X1  g728(.A1(new_n717_), .A2(new_n468_), .A3(new_n461_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n849_), .A2(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(new_n507_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g732(.A1(new_n931_), .A2(new_n604_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g734(.A(KEYINPUT63), .B(G211gat), .C1(new_n931_), .C2(new_n688_), .ZN(new_n936_));
  NOR3_X1   g735(.A1(new_n849_), .A2(new_n621_), .A3(new_n930_), .ZN(new_n937_));
  XOR2_X1   g736(.A(KEYINPUT63), .B(G211gat), .Z(new_n938_));
  AOI21_X1  g737(.A(new_n936_), .B1(new_n937_), .B2(new_n938_), .ZN(G1354gat));
  INV_X1    g738(.A(G218gat), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n931_), .A2(new_n940_), .A3(new_n662_), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n849_), .A2(new_n651_), .A3(new_n930_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n941_), .B1(new_n942_), .B2(new_n940_), .ZN(G1355gat));
endmodule


