//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1 0 1 0 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n786_, new_n787_, new_n788_, new_n790_, new_n791_,
    new_n792_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n881_,
    new_n883_, new_n885_, new_n886_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n916_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G169gat), .ZN(new_n202_));
  INV_X1    g001(.A(G176gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  AOI21_X1  g003(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND3_X1  g005(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n207_));
  INV_X1    g006(.A(G183gat), .ZN(new_n208_));
  INV_X1    g007(.A(G190gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n206_), .A2(new_n207_), .A3(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n204_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT78), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(KEYINPUT24), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n218_), .A2(KEYINPUT78), .A3(KEYINPUT24), .A4(new_n212_), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n208_), .A2(KEYINPUT25), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT25), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(G183gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n209_), .A2(KEYINPUT26), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT26), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(G190gat), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n221_), .A2(new_n223_), .A3(new_n224_), .A4(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n207_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n228_), .A2(new_n205_), .ZN(new_n229_));
  NOR3_X1   g028(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n227_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n213_), .B1(new_n220_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT79), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n217_), .A2(new_n219_), .ZN(new_n235_));
  NOR3_X1   g034(.A1(new_n228_), .A2(new_n230_), .A3(new_n205_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n236_), .A3(new_n227_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT79), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(new_n238_), .A3(new_n213_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n234_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G71gat), .B(G99gat), .ZN(new_n241_));
  INV_X1    g040(.A(G43gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n240_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G127gat), .B(G134gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT80), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G113gat), .B(G120gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n244_), .B(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G227gat), .A2(G233gat), .ZN(new_n250_));
  INV_X1    g049(.A(G15gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT30), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT31), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n249_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n249_), .A2(new_n255_), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(G155gat), .ZN(new_n260_));
  INV_X1    g059(.A(G162gat), .ZN(new_n261_));
  OR3_X1    g060(.A1(new_n260_), .A2(new_n261_), .A3(KEYINPUT1), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT1), .B1(new_n260_), .B2(new_n261_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n262_), .B(new_n263_), .C1(G155gat), .C2(G162gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G141gat), .A2(G148gat), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT81), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(G141gat), .ZN(new_n269_));
  INV_X1    g068(.A(G148gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT82), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n269_), .A2(new_n270_), .A3(KEYINPUT82), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n264_), .A2(new_n268_), .A3(new_n273_), .A4(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(G155gat), .B(G162gat), .Z(new_n276_));
  NOR2_X1   g075(.A1(new_n267_), .A2(KEYINPUT2), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n271_), .A2(KEYINPUT3), .ZN(new_n278_));
  OR3_X1    g077(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT2), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n278_), .B(new_n279_), .C1(new_n280_), .C2(new_n265_), .ZN(new_n281_));
  OAI211_X1 g080(.A(KEYINPUT83), .B(new_n276_), .C1(new_n277_), .C2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n265_), .A2(new_n280_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n284_), .B1(KEYINPUT3), .B2(new_n271_), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n285_), .B(new_n279_), .C1(new_n267_), .C2(KEYINPUT2), .ZN(new_n286_));
  AOI21_X1  g085(.A(KEYINPUT83), .B1(new_n286_), .B2(new_n276_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n275_), .B1(new_n283_), .B2(new_n287_), .ZN(new_n288_));
  OR3_X1    g087(.A1(new_n288_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT28), .B1(new_n288_), .B2(KEYINPUT29), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G22gat), .B(G50gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n288_), .A2(KEYINPUT29), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT85), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT87), .ZN(new_n296_));
  INV_X1    g095(.A(G204gat), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT86), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n298_), .A2(G197gat), .ZN(new_n299_));
  INV_X1    g098(.A(G197gat), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n300_), .A2(KEYINPUT86), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n296_), .B(new_n297_), .C1(new_n299_), .C2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT21), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n300_), .A2(KEYINPUT86), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n298_), .A2(G197gat), .ZN(new_n305_));
  AOI21_X1  g104(.A(G204gat), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n296_), .B1(new_n300_), .B2(G204gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT88), .B1(new_n303_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT21), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n311_), .B1(new_n306_), .B2(new_n296_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT88), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT86), .B(G197gat), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n307_), .B1(new_n314_), .B2(G204gat), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n312_), .A2(new_n313_), .A3(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(G197gat), .A2(G204gat), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n318_), .B1(new_n314_), .B2(new_n297_), .ZN(new_n319_));
  INV_X1    g118(.A(G211gat), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n320_), .A2(G218gat), .ZN(new_n321_));
  INV_X1    g120(.A(G218gat), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n322_), .A2(G211gat), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT89), .B1(new_n321_), .B2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(G211gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n320_), .A2(G218gat), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT89), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n325_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  AOI22_X1  g127(.A1(new_n319_), .A2(new_n311_), .B1(new_n324_), .B2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n310_), .A2(new_n316_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT90), .ZN(new_n331_));
  INV_X1    g130(.A(new_n328_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n327_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n331_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n324_), .A2(KEYINPUT90), .A3(new_n328_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n297_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n336_));
  NOR3_X1   g135(.A1(new_n336_), .A2(new_n311_), .A3(new_n317_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n334_), .A2(new_n335_), .A3(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n330_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n294_), .A2(new_n295_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(G233gat), .ZN(new_n341_));
  NOR2_X1   g140(.A1(KEYINPUT84), .A2(G228gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(KEYINPUT84), .A2(G228gat), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n341_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n340_), .A2(new_n345_), .ZN(new_n346_));
  AND3_X1   g145(.A1(new_n334_), .A2(new_n335_), .A3(new_n337_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n313_), .B1(new_n312_), .B2(new_n315_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n324_), .A2(new_n328_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n336_), .A2(new_n317_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n349_), .B1(new_n350_), .B2(KEYINPUT21), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n348_), .A2(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n347_), .B1(new_n352_), .B2(new_n316_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n353_), .A2(KEYINPUT85), .ZN(new_n354_));
  INV_X1    g153(.A(new_n345_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(new_n355_), .A3(new_n294_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G78gat), .B(G106gat), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n346_), .A2(new_n356_), .A3(new_n358_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n293_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT93), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n346_), .A2(new_n356_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n358_), .B1(new_n362_), .B2(KEYINPUT92), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT92), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n346_), .A2(new_n364_), .A3(new_n356_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n361_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n356_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n355_), .B1(new_n354_), .B2(new_n294_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT92), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  AND4_X1   g168(.A1(new_n361_), .A2(new_n369_), .A3(new_n357_), .A4(new_n365_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n360_), .B1(new_n366_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT91), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n359_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n362_), .A2(new_n357_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n346_), .A2(KEYINPUT91), .A3(new_n356_), .A4(new_n358_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n373_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n293_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n371_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G225gat), .A2(G233gat), .ZN(new_n380_));
  INV_X1    g179(.A(new_n248_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n288_), .A2(new_n381_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n248_), .B(new_n275_), .C1(new_n287_), .C2(new_n283_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(KEYINPUT4), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT4), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n288_), .A2(new_n385_), .A3(new_n381_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n380_), .B1(new_n384_), .B2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G1gat), .B(G29gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(G85gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT0), .B(G57gat), .ZN(new_n390_));
  XOR2_X1   g189(.A(new_n389_), .B(new_n390_), .Z(new_n391_));
  INV_X1    g190(.A(new_n380_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n392_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n393_));
  OR3_X1    g192(.A1(new_n387_), .A2(new_n391_), .A3(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n391_), .B1(new_n387_), .B2(new_n393_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT27), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n212_), .A2(KEYINPUT97), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n212_), .A2(KEYINPUT97), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n204_), .A2(new_n211_), .A3(new_n399_), .A4(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT94), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n215_), .A2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n212_), .A2(KEYINPUT94), .A3(KEYINPUT24), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n404_), .A2(new_n218_), .A3(new_n405_), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n406_), .A2(KEYINPUT95), .A3(new_n227_), .ZN(new_n407_));
  AOI21_X1  g206(.A(KEYINPUT95), .B1(new_n406_), .B2(new_n227_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n236_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n402_), .B1(new_n409_), .B2(KEYINPUT96), .ZN(new_n410_));
  INV_X1    g209(.A(new_n236_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT95), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n212_), .A2(KEYINPUT94), .A3(KEYINPUT24), .ZN(new_n413_));
  AOI21_X1  g212(.A(KEYINPUT94), .B1(new_n212_), .B2(KEYINPUT24), .ZN(new_n414_));
  NOR3_X1   g213(.A1(new_n413_), .A2(new_n414_), .A3(new_n216_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n227_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n412_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n406_), .A2(KEYINPUT95), .A3(new_n227_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n411_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT96), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n410_), .A2(new_n353_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT99), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT99), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n410_), .A2(new_n353_), .A3(new_n424_), .A4(new_n421_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT20), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n427_), .B1(new_n339_), .B2(new_n240_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G226gat), .A2(G233gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT19), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n426_), .A2(new_n433_), .ZN(new_n434_));
  XOR2_X1   g233(.A(G8gat), .B(G36gat), .Z(new_n435_));
  XNOR2_X1  g234(.A(G64gat), .B(G92gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n401_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n409_), .A2(KEYINPUT96), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n339_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n237_), .A2(new_n238_), .A3(new_n213_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n238_), .B1(new_n237_), .B2(new_n213_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n427_), .B1(new_n353_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n443_), .A2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT98), .B1(new_n448_), .B2(new_n430_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT98), .ZN(new_n450_));
  AOI211_X1 g249(.A(new_n450_), .B(new_n431_), .C1(new_n443_), .C2(new_n447_), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n434_), .B(new_n440_), .C1(new_n449_), .C2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n410_), .A2(new_n421_), .B1(new_n330_), .B2(new_n338_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT20), .B1(new_n339_), .B2(new_n240_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n430_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n450_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n448_), .A2(KEYINPUT98), .A3(new_n430_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n440_), .B1(new_n459_), .B2(new_n434_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n398_), .B1(new_n453_), .B2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n432_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n462_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n398_), .B1(new_n463_), .B2(new_n440_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n443_), .A2(new_n447_), .A3(new_n431_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT102), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n443_), .A2(new_n447_), .A3(KEYINPUT102), .A4(new_n431_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n330_), .A2(new_n409_), .A3(new_n338_), .A4(new_n401_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n431_), .B1(new_n428_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n467_), .A2(new_n468_), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(new_n439_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT103), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n472_), .A2(KEYINPUT103), .A3(new_n439_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n464_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n379_), .A2(new_n397_), .A3(new_n461_), .A4(new_n477_), .ZN(new_n478_));
  AND2_X1   g277(.A1(new_n440_), .A2(KEYINPUT32), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n472_), .A2(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n434_), .B1(new_n449_), .B2(new_n451_), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n479_), .B(KEYINPUT101), .Z(new_n482_));
  OAI211_X1 g281(.A(new_n396_), .B(new_n480_), .C1(new_n481_), .C2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n439_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n452_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT33), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n395_), .A2(new_n486_), .ZN(new_n487_));
  OAI211_X1 g286(.A(KEYINPUT33), .B(new_n391_), .C1(new_n387_), .C2(new_n393_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n384_), .A2(new_n380_), .A3(new_n386_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n391_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n382_), .A2(new_n392_), .A3(new_n383_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n487_), .A2(new_n488_), .A3(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n483_), .B1(new_n485_), .B2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n369_), .A2(new_n357_), .A3(new_n365_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT93), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n363_), .A2(new_n361_), .A3(new_n365_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  AOI22_X1  g297(.A1(new_n498_), .A2(new_n360_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n494_), .A2(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n259_), .B1(new_n478_), .B2(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n258_), .A2(new_n396_), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n477_), .A2(new_n461_), .A3(KEYINPUT104), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT104), .B1(new_n477_), .B2(new_n461_), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n499_), .B(new_n502_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT105), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT104), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n452_), .A2(KEYINPUT27), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n470_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n509_));
  AOI211_X1 g308(.A(new_n474_), .B(new_n440_), .C1(new_n509_), .C2(new_n468_), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT103), .B1(new_n472_), .B2(new_n439_), .ZN(new_n511_));
  NOR3_X1   g310(.A1(new_n508_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(KEYINPUT27), .B1(new_n484_), .B2(new_n452_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n507_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n477_), .A2(new_n461_), .A3(KEYINPUT104), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT105), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n516_), .A2(new_n517_), .A3(new_n499_), .A4(new_n502_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n501_), .B1(new_n506_), .B2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G15gat), .B(G22gat), .ZN(new_n520_));
  INV_X1    g319(.A(G1gat), .ZN(new_n521_));
  INV_X1    g320(.A(G8gat), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT14), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G1gat), .B(G8gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G29gat), .B(G36gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G43gat), .B(G50gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  XOR2_X1   g328(.A(new_n526_), .B(new_n529_), .Z(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT76), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n531_), .A2(G229gat), .A3(G233gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n529_), .B(KEYINPUT15), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(new_n526_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G229gat), .A2(G233gat), .ZN(new_n535_));
  INV_X1    g334(.A(new_n526_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(new_n529_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n534_), .A2(new_n535_), .A3(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n532_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G113gat), .B(G141gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT77), .ZN(new_n541_));
  XOR2_X1   g340(.A(G169gat), .B(G197gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n539_), .B(new_n543_), .Z(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  XOR2_X1   g344(.A(G57gat), .B(G64gat), .Z(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT67), .B(G71gat), .ZN(new_n547_));
  INV_X1    g346(.A(G78gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT11), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n546_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n547_), .B(G78gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT11), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n552_), .A2(KEYINPUT11), .A3(new_n546_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G231gat), .A2(G233gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT74), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(new_n526_), .ZN(new_n560_));
  XOR2_X1   g359(.A(G127gat), .B(G155gat), .Z(new_n561_));
  XNOR2_X1  g360(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G183gat), .B(G211gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(KEYINPUT17), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n560_), .A2(new_n566_), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n565_), .A2(KEYINPUT17), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n560_), .A2(new_n566_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G99gat), .A2(G106gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT6), .ZN(new_n573_));
  XOR2_X1   g372(.A(KEYINPUT10), .B(G99gat), .Z(new_n574_));
  INV_X1    g373(.A(G106gat), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G85gat), .A2(G92gat), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n580_), .A2(KEYINPUT65), .ZN(new_n581_));
  INV_X1    g380(.A(G85gat), .ZN(new_n582_));
  INV_X1    g381(.A(G92gat), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n579_), .A2(KEYINPUT9), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n584_), .B(new_n585_), .C1(new_n580_), .C2(KEYINPUT65), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n573_), .B(new_n576_), .C1(new_n581_), .C2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n584_), .A2(new_n578_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT66), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT8), .ZN(new_n591_));
  OAI21_X1  g390(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n592_));
  OR3_X1    g391(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n573_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n590_), .A2(new_n591_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n591_), .B1(new_n590_), .B2(new_n594_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n587_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n556_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT12), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n556_), .A2(new_n598_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n599_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G230gat), .A2(G233gat), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n598_), .A2(KEYINPUT69), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n554_), .A2(new_n555_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n605_), .A2(new_n600_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT69), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n607_), .B(new_n587_), .C1(new_n596_), .C2(new_n597_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n604_), .A2(new_n606_), .A3(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n602_), .A2(new_n603_), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n598_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(new_n605_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n612_), .A2(KEYINPUT68), .A3(new_n601_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n603_), .ZN(new_n614_));
  OR3_X1    g413(.A1(new_n556_), .A2(new_n598_), .A3(KEYINPUT68), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n613_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n610_), .A2(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G120gat), .B(G148gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT5), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G176gat), .B(G204gat), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n619_), .B(new_n620_), .Z(new_n621_));
  NAND2_X1  g420(.A1(new_n617_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n621_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n610_), .A2(new_n616_), .A3(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT13), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n622_), .A2(KEYINPUT13), .A3(new_n624_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT72), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT35), .ZN(new_n632_));
  NAND2_X1  g431(.A1(G232gat), .A2(G233gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT71), .ZN(new_n634_));
  XOR2_X1   g433(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  AOI22_X1  g435(.A1(new_n611_), .A2(new_n529_), .B1(new_n632_), .B2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n604_), .A2(new_n533_), .A3(new_n608_), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n636_), .A2(new_n632_), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n637_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n639_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(G190gat), .B(G218gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(G134gat), .B(G162gat), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(KEYINPUT36), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n631_), .B1(new_n642_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n646_), .ZN(new_n648_));
  NOR4_X1   g447(.A1(new_n640_), .A2(new_n641_), .A3(KEYINPUT72), .A4(new_n648_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n645_), .A2(KEYINPUT36), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n648_), .B(new_n651_), .C1(new_n640_), .C2(new_n641_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n650_), .A2(KEYINPUT73), .A3(KEYINPUT37), .A4(new_n652_), .ZN(new_n653_));
  OAI211_X1 g452(.A(new_n652_), .B(KEYINPUT73), .C1(new_n647_), .C2(new_n649_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT37), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n571_), .A2(new_n630_), .A3(new_n653_), .A4(new_n656_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n519_), .A2(new_n545_), .A3(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n658_), .A2(new_n521_), .A3(new_n396_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT38), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n650_), .A2(new_n652_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n519_), .A2(new_n663_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n629_), .A2(new_n545_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n664_), .A2(new_n571_), .A3(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(G1gat), .B1(new_n666_), .B2(new_n397_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n659_), .A2(new_n660_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n661_), .A2(new_n667_), .A3(new_n668_), .ZN(G1324gat));
  NOR2_X1   g468(.A1(new_n503_), .A2(new_n504_), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n658_), .A2(new_n522_), .A3(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(G8gat), .B1(new_n666_), .B2(new_n516_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT39), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT39), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n674_), .B(G8gat), .C1(new_n666_), .C2(new_n516_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n671_), .B1(new_n673_), .B2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n676_), .B(new_n678_), .ZN(G1325gat));
  INV_X1    g478(.A(new_n666_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n251_), .B1(new_n680_), .B2(new_n259_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n682_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n658_), .A2(new_n251_), .A3(new_n259_), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n685_), .B(KEYINPUT107), .Z(new_n686_));
  NAND3_X1  g485(.A1(new_n683_), .A2(new_n684_), .A3(new_n686_), .ZN(G1326gat));
  INV_X1    g486(.A(G22gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n658_), .A2(new_n688_), .A3(new_n379_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G22gat), .B1(new_n666_), .B2(new_n499_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n690_), .A2(KEYINPUT42), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(KEYINPUT42), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n689_), .B1(new_n691_), .B2(new_n692_), .ZN(G1327gat));
  NOR2_X1   g492(.A1(new_n519_), .A2(new_n545_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n570_), .A2(new_n663_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n695_), .A2(new_n629_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G29gat), .B1(new_n698_), .B2(new_n396_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n570_), .A2(new_n665_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n702_));
  INV_X1    g501(.A(new_n501_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n505_), .A2(KEYINPUT105), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n379_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n517_), .B1(new_n705_), .B2(new_n502_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n703_), .B1(new_n704_), .B2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n653_), .A2(new_n656_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n702_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n708_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n519_), .A2(KEYINPUT43), .A3(new_n710_), .ZN(new_n711_));
  OAI211_X1 g510(.A(KEYINPUT44), .B(new_n701_), .C1(new_n709_), .C2(new_n711_), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n712_), .A2(G29gat), .A3(new_n396_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n701_), .B1(new_n709_), .B2(new_n711_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n699_), .B1(new_n713_), .B2(new_n716_), .ZN(G1328gat));
  INV_X1    g516(.A(G36gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n707_), .A2(new_n702_), .A3(new_n708_), .ZN(new_n719_));
  OAI21_X1  g518(.A(KEYINPUT43), .B1(new_n519_), .B2(new_n710_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n700_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n516_), .B1(new_n721_), .B2(KEYINPUT44), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n718_), .B1(new_n722_), .B2(new_n716_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n516_), .A2(G36gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n694_), .A2(new_n696_), .A3(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT45), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n694_), .A2(new_n727_), .A3(new_n696_), .A4(new_n724_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n723_), .A2(new_n730_), .A3(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n712_), .A2(new_n670_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n721_), .A2(KEYINPUT44), .ZN(new_n735_));
  OAI21_X1  g534(.A(G36gat), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n731_), .B1(new_n736_), .B2(new_n729_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n733_), .A2(new_n737_), .ZN(G1329gat));
  OAI21_X1  g537(.A(new_n242_), .B1(new_n697_), .B2(new_n258_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n712_), .A2(G43gat), .A3(new_n259_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n740_), .B2(new_n735_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g541(.A(G50gat), .B1(new_n698_), .B2(new_n379_), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n712_), .A2(G50gat), .A3(new_n379_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n744_), .B2(new_n716_), .ZN(G1331gat));
  NOR2_X1   g544(.A1(new_n519_), .A2(new_n544_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n708_), .A2(new_n570_), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n746_), .A2(new_n629_), .A3(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(G57gat), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n748_), .A2(new_n749_), .A3(new_n396_), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n664_), .A2(new_n545_), .A3(new_n629_), .A4(new_n571_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n751_), .A2(KEYINPUT109), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(KEYINPUT109), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n752_), .A2(new_n396_), .A3(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n750_), .B1(new_n754_), .B2(new_n749_), .ZN(G1332gat));
  INV_X1    g554(.A(G64gat), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n748_), .A2(new_n756_), .A3(new_n670_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n752_), .A2(new_n670_), .A3(new_n753_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT48), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n758_), .A2(new_n759_), .A3(G64gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n758_), .B2(G64gat), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n757_), .B1(new_n760_), .B2(new_n761_), .ZN(G1333gat));
  NOR2_X1   g561(.A1(new_n258_), .A2(G71gat), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT111), .Z(new_n764_));
  NAND2_X1  g563(.A1(new_n748_), .A2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n752_), .A2(new_n259_), .A3(new_n753_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n766_), .A2(G71gat), .A3(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n766_), .B2(G71gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n765_), .B1(new_n768_), .B2(new_n769_), .ZN(G1334gat));
  NAND3_X1  g569(.A1(new_n748_), .A2(new_n548_), .A3(new_n379_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n752_), .A2(new_n379_), .A3(new_n753_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT50), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n772_), .A2(new_n773_), .A3(G78gat), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n773_), .B1(new_n772_), .B2(G78gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n771_), .B1(new_n774_), .B2(new_n775_), .ZN(G1335gat));
  NAND3_X1  g575(.A1(new_n570_), .A2(new_n545_), .A3(new_n629_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n777_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(G85gat), .B1(new_n779_), .B2(new_n397_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n695_), .A2(new_n630_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n746_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(new_n582_), .A3(new_n396_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n780_), .A2(new_n784_), .ZN(G1336gat));
  OAI21_X1  g584(.A(new_n583_), .B1(new_n782_), .B2(new_n516_), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n786_), .B(KEYINPUT112), .Z(new_n787_));
  NOR3_X1   g586(.A1(new_n779_), .A2(new_n583_), .A3(new_n516_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(G1337gat));
  NAND2_X1  g588(.A1(new_n778_), .A2(new_n259_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n259_), .A2(new_n574_), .ZN(new_n791_));
  AOI22_X1  g590(.A1(new_n790_), .A2(G99gat), .B1(new_n783_), .B2(new_n791_), .ZN(new_n792_));
  XOR2_X1   g591(.A(new_n792_), .B(KEYINPUT51), .Z(G1338gat));
  XNOR2_X1  g592(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797_));
  OAI21_X1  g596(.A(G106gat), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n798_), .B1(new_n778_), .B2(new_n379_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n796_), .A2(new_n797_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n783_), .A2(new_n575_), .A3(new_n379_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n803_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n795_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n799_), .A2(new_n800_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n806_), .A2(new_n801_), .A3(new_n803_), .A4(new_n794_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(G1339gat));
  NAND2_X1  g607(.A1(new_n601_), .A2(new_n600_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n612_), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n604_), .A2(new_n606_), .A3(new_n608_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n810_), .A2(new_n811_), .A3(new_n614_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n614_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n813_), .B2(KEYINPUT55), .ZN(new_n814_));
  AND4_X1   g613(.A1(KEYINPUT55), .A2(new_n602_), .A3(new_n603_), .A4(new_n609_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n621_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT56), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT56), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n818_), .B(new_n621_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n817_), .A2(new_n624_), .A3(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n539_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n531_), .A2(new_n535_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n535_), .B1(new_n536_), .B2(new_n529_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n543_), .B1(new_n534_), .B2(new_n823_), .ZN(new_n824_));
  AOI22_X1  g623(.A1(new_n821_), .A2(new_n543_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT58), .B1(new_n820_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n624_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n827_), .B1(new_n816_), .B2(KEYINPUT56), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n828_), .A2(KEYINPUT58), .A3(new_n825_), .A4(new_n819_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n708_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n817_), .A2(new_n544_), .A3(new_n624_), .A4(new_n819_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n825_), .A2(new_n625_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n663_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  OAI22_X1  g632(.A1(new_n826_), .A2(new_n830_), .B1(new_n833_), .B2(KEYINPUT57), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n833_), .A2(KEYINPUT57), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n570_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(KEYINPUT54), .B1(new_n657_), .B2(new_n544_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n747_), .A2(new_n838_), .A3(new_n545_), .A4(new_n630_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT115), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n705_), .A2(new_n396_), .A3(new_n259_), .ZN(new_n842_));
  AOI22_X1  g641(.A1(new_n836_), .A2(new_n840_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  OR2_X1    g642(.A1(new_n842_), .A2(new_n841_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(KEYINPUT59), .A3(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT59), .B1(new_n843_), .B2(new_n844_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(G113gat), .B1(new_n848_), .B2(new_n545_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n836_), .A2(new_n840_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n842_), .A2(new_n841_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n850_), .A2(new_n844_), .A3(new_n851_), .ZN(new_n852_));
  OR3_X1    g651(.A1(new_n852_), .A2(G113gat), .A3(new_n545_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n849_), .A2(new_n853_), .ZN(G1340gat));
  OAI21_X1  g653(.A(G120gat), .B1(new_n848_), .B2(new_n630_), .ZN(new_n855_));
  INV_X1    g654(.A(G120gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n856_), .B1(new_n630_), .B2(KEYINPUT60), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(KEYINPUT60), .B2(new_n856_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n855_), .B1(new_n852_), .B2(new_n858_), .ZN(G1341gat));
  OAI21_X1  g658(.A(G127gat), .B1(new_n848_), .B2(new_n570_), .ZN(new_n860_));
  OR3_X1    g659(.A1(new_n852_), .A2(G127gat), .A3(new_n570_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1342gat));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n850_), .A2(new_n663_), .A3(new_n844_), .A4(new_n851_), .ZN(new_n864_));
  INV_X1    g663(.A(G134gat), .ZN(new_n865_));
  AND3_X1   g664(.A1(new_n864_), .A2(KEYINPUT116), .A3(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(KEYINPUT116), .B1(new_n864_), .B2(new_n865_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(KEYINPUT117), .B(G134gat), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n710_), .A2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n852_), .A2(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n871_), .B1(new_n873_), .B2(new_n845_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n863_), .B1(new_n868_), .B2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n870_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n876_), .B(KEYINPUT118), .C1(new_n867_), .C2(new_n866_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(G1343gat));
  NOR3_X1   g677(.A1(new_n499_), .A2(new_n397_), .A3(new_n259_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n850_), .A2(new_n516_), .A3(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n880_), .A2(new_n545_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(new_n269_), .ZN(G1344gat));
  NOR2_X1   g681(.A1(new_n880_), .A2(new_n630_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(new_n270_), .ZN(G1345gat));
  NOR2_X1   g683(.A1(new_n880_), .A2(new_n570_), .ZN(new_n885_));
  XOR2_X1   g684(.A(KEYINPUT61), .B(G155gat), .Z(new_n886_));
  XNOR2_X1  g685(.A(new_n885_), .B(new_n886_), .ZN(G1346gat));
  OAI21_X1  g686(.A(G162gat), .B1(new_n880_), .B2(new_n710_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n663_), .A2(new_n261_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n880_), .B2(new_n889_), .ZN(G1347gat));
  NAND2_X1  g689(.A1(new_n850_), .A2(new_n499_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n670_), .A2(new_n502_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n893_), .A2(new_n202_), .A3(new_n544_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT62), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n892_), .A2(new_n545_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(KEYINPUT119), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n850_), .A2(new_n499_), .A3(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n895_), .B1(new_n898_), .B2(G169gat), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n898_), .A2(new_n895_), .A3(G169gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n894_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(KEYINPUT120), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n894_), .B(new_n903_), .C1(new_n899_), .C2(new_n900_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n904_), .ZN(G1348gat));
  AOI21_X1  g704(.A(G176gat), .B1(new_n893_), .B2(new_n629_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n891_), .B(KEYINPUT121), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n892_), .A2(new_n203_), .A3(new_n630_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n906_), .B1(new_n907_), .B2(new_n908_), .ZN(G1349gat));
  NAND2_X1  g708(.A1(new_n221_), .A2(new_n223_), .ZN(new_n910_));
  AND3_X1   g709(.A1(new_n893_), .A2(new_n910_), .A3(new_n571_), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n907_), .A2(new_n670_), .A3(new_n502_), .A4(new_n571_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n911_), .B1(new_n912_), .B2(new_n208_), .ZN(G1350gat));
  INV_X1    g712(.A(new_n893_), .ZN(new_n914_));
  OAI21_X1  g713(.A(G190gat), .B1(new_n914_), .B2(new_n710_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n663_), .A2(new_n224_), .A3(new_n226_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n914_), .B2(new_n916_), .ZN(G1351gat));
  NOR4_X1   g716(.A1(new_n516_), .A2(new_n499_), .A3(new_n396_), .A4(new_n259_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n850_), .A2(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n919_), .A2(new_n545_), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n920_), .A2(KEYINPUT122), .A3(G197gat), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n300_), .B1(new_n919_), .B2(new_n545_), .ZN(new_n922_));
  AND2_X1   g721(.A1(new_n922_), .A2(KEYINPUT122), .ZN(new_n923_));
  AOI211_X1 g722(.A(new_n921_), .B(new_n923_), .C1(G197gat), .C2(new_n920_), .ZN(G1352gat));
  INV_X1    g723(.A(new_n919_), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT124), .ZN(new_n926_));
  OAI211_X1 g725(.A(new_n925_), .B(new_n629_), .C1(new_n926_), .C2(new_n297_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n297_), .B2(KEYINPUT123), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n927_), .B(new_n928_), .ZN(G1353gat));
  AOI21_X1  g728(.A(new_n570_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n925_), .A2(new_n930_), .ZN(new_n931_));
  AND2_X1   g730(.A1(new_n931_), .A2(KEYINPUT125), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n931_), .A2(KEYINPUT125), .ZN(new_n933_));
  OAI22_X1  g732(.A1(new_n932_), .A2(new_n933_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n934_));
  OR2_X1    g733(.A1(new_n931_), .A2(KEYINPUT125), .ZN(new_n935_));
  NOR2_X1   g734(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n931_), .A2(KEYINPUT125), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n935_), .A2(new_n936_), .A3(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n934_), .A2(new_n938_), .ZN(G1354gat));
  XOR2_X1   g738(.A(KEYINPUT126), .B(G218gat), .Z(new_n940_));
  NOR3_X1   g739(.A1(new_n919_), .A2(new_n710_), .A3(new_n940_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n925_), .A2(new_n663_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n941_), .B1(new_n942_), .B2(new_n940_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n943_), .B(new_n944_), .ZN(G1355gat));
endmodule


