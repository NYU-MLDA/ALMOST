//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 1 1 1 1 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n818_, new_n819_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n829_, new_n830_, new_n831_, new_n832_, new_n834_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n866_, new_n867_, new_n868_, new_n870_, new_n871_,
    new_n872_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_;
  INV_X1    g000(.A(KEYINPUT78), .ZN(new_n202_));
  XOR2_X1   g001(.A(G15gat), .B(G22gat), .Z(new_n203_));
  NAND2_X1  g002(.A1(G1gat), .A2(G8gat), .ZN(new_n204_));
  AOI21_X1  g003(.A(new_n203_), .B1(KEYINPUT14), .B2(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT73), .ZN(new_n206_));
  XOR2_X1   g005(.A(G1gat), .B(G8gat), .Z(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT73), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n205_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n207_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n208_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G29gat), .B(G36gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G43gat), .B(G50gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT15), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n213_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n208_), .A2(new_n212_), .A3(new_n216_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G229gat), .A2(G233gat), .ZN(new_n220_));
  XOR2_X1   g019(.A(new_n220_), .B(KEYINPUT77), .Z(new_n221_));
  NAND3_X1  g020(.A1(new_n218_), .A2(new_n219_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n216_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n213_), .A2(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n220_), .B1(new_n225_), .B2(new_n219_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G113gat), .B(G141gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G169gat), .B(G197gat), .ZN(new_n228_));
  XOR2_X1   g027(.A(new_n227_), .B(new_n228_), .Z(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NOR3_X1   g029(.A1(new_n223_), .A2(new_n226_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n225_), .A2(new_n219_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n220_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n229_), .B1(new_n234_), .B2(new_n222_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n202_), .B1(new_n231_), .B2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n230_), .B1(new_n223_), .B2(new_n226_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n234_), .A2(new_n222_), .A3(new_n229_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(new_n238_), .A3(KEYINPUT78), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n236_), .A2(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n240_), .B(KEYINPUT79), .Z(new_n241_));
  INV_X1    g040(.A(G197gat), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n242_), .A2(G204gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT88), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT89), .B(G204gat), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n245_), .A2(G197gat), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT21), .B1(new_n244_), .B2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G211gat), .B(G218gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT91), .ZN(new_n249_));
  MUX2_X1   g048(.A(G204gat), .B(new_n245_), .S(G197gat), .Z(new_n250_));
  XOR2_X1   g049(.A(KEYINPUT90), .B(KEYINPUT21), .Z(new_n251_));
  OAI211_X1 g050(.A(new_n247_), .B(new_n249_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(KEYINPUT92), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n248_), .B(KEYINPUT91), .Z(new_n254_));
  INV_X1    g053(.A(KEYINPUT92), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n245_), .A2(new_n242_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(G197gat), .A2(G204gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n255_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n253_), .A2(new_n254_), .A3(KEYINPUT21), .A4(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n252_), .A2(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(G141gat), .A2(G148gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT3), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G141gat), .A2(G148gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT2), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G155gat), .B(G162gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT85), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n261_), .B(new_n267_), .ZN(new_n268_));
  AND2_X1   g067(.A1(G155gat), .A2(G162gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT1), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n268_), .A2(new_n263_), .A3(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n266_), .A2(KEYINPUT1), .ZN(new_n272_));
  OAI22_X1  g071(.A1(new_n265_), .A2(new_n266_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT29), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n260_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(G233gat), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT87), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n277_), .A2(G228gat), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(G228gat), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n276_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n275_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G78gat), .B(G106gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT93), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n273_), .A2(KEYINPUT29), .ZN(new_n286_));
  XOR2_X1   g085(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n287_));
  XNOR2_X1  g086(.A(G22gat), .B(G50gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n286_), .B(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n285_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n282_), .B(new_n283_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G227gat), .A2(G233gat), .ZN(new_n294_));
  XOR2_X1   g093(.A(new_n294_), .B(KEYINPUT83), .Z(new_n295_));
  OR2_X1    g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n296_), .A2(KEYINPUT24), .A3(new_n297_), .ZN(new_n298_));
  XOR2_X1   g097(.A(KEYINPUT25), .B(G183gat), .Z(new_n299_));
  XOR2_X1   g098(.A(KEYINPUT26), .B(G190gat), .Z(new_n300_));
  OAI221_X1 g099(.A(new_n298_), .B1(KEYINPUT24), .B2(new_n296_), .C1(new_n299_), .C2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT23), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n302_), .A2(G183gat), .A3(G190gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT80), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n302_), .B1(G183gat), .B2(G190gat), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n301_), .A2(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(KEYINPUT82), .B(G176gat), .Z(new_n309_));
  INV_X1    g108(.A(KEYINPUT81), .ZN(new_n310_));
  INV_X1    g109(.A(G169gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT22), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n311_), .A2(KEYINPUT22), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n309_), .B(new_n312_), .C1(new_n310_), .C2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(G183gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n315_), .A2(KEYINPUT23), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n306_), .B1(G190gat), .B2(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(G183gat), .A2(G190gat), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n314_), .B(new_n297_), .C1(new_n317_), .C2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n308_), .A2(KEYINPUT30), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(G15gat), .B(G43gat), .Z(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT30), .B1(new_n308_), .B2(new_n319_), .ZN(new_n323_));
  NOR3_X1   g122(.A1(new_n321_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n322_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n308_), .A2(new_n319_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT30), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n325_), .B1(new_n328_), .B2(new_n320_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n295_), .B1(new_n324_), .B2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G71gat), .B(G99gat), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n322_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n295_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n328_), .A2(new_n325_), .A3(new_n320_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n332_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n330_), .A2(new_n331_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT84), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n331_), .B1(new_n330_), .B2(new_n335_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT31), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(G127gat), .B(G134gat), .Z(new_n341_));
  XOR2_X1   g140(.A(G113gat), .B(G120gat), .Z(new_n342_));
  XOR2_X1   g141(.A(new_n341_), .B(new_n342_), .Z(new_n343_));
  NAND2_X1  g142(.A1(new_n330_), .A2(new_n335_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n331_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT31), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n346_), .A2(new_n337_), .A3(new_n347_), .A4(new_n336_), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n340_), .A2(new_n343_), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n343_), .B1(new_n340_), .B2(new_n348_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n293_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n340_), .A2(new_n348_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n343_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n291_), .B(new_n292_), .Z(new_n355_));
  NAND3_X1  g154(.A1(new_n340_), .A2(new_n343_), .A3(new_n348_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n351_), .A2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n307_), .A2(new_n318_), .ZN(new_n359_));
  XOR2_X1   g158(.A(KEYINPUT22), .B(G169gat), .Z(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n309_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(new_n297_), .ZN(new_n363_));
  OAI22_X1  g162(.A1(new_n359_), .A2(new_n363_), .B1(new_n301_), .B2(new_n317_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n260_), .A2(new_n364_), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n365_), .B(KEYINPUT20), .C1(new_n260_), .C2(new_n326_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT94), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G226gat), .A2(G233gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT19), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n366_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT20), .B1(new_n260_), .B2(new_n364_), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n260_), .A2(new_n326_), .ZN(new_n373_));
  OR3_X1    g172(.A1(new_n372_), .A2(new_n373_), .A3(new_n369_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n367_), .B1(new_n366_), .B2(new_n369_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n371_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G8gat), .B(G36gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT18), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G64gat), .B(G92gat), .ZN(new_n379_));
  XOR2_X1   g178(.A(new_n378_), .B(new_n379_), .Z(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT27), .B1(new_n376_), .B2(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n369_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n383_));
  OR2_X1    g182(.A1(new_n383_), .A2(KEYINPUT97), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n366_), .A2(new_n369_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(KEYINPUT97), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n384_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n387_), .A2(new_n381_), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT98), .B1(new_n382_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n375_), .A2(new_n374_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n381_), .B1(new_n390_), .B2(new_n370_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n387_), .A2(new_n381_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT98), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n392_), .A2(new_n393_), .A3(new_n394_), .A4(KEYINPUT27), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n353_), .B(new_n273_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT4), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT4), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n273_), .A2(new_n398_), .A3(new_n343_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G225gat), .A2(G233gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT95), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n397_), .A2(new_n399_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n396_), .A2(new_n400_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G1gat), .B(G29gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(G85gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT0), .B(G57gat), .ZN(new_n406_));
  XOR2_X1   g205(.A(new_n405_), .B(new_n406_), .Z(new_n407_));
  NAND3_X1  g206(.A1(new_n402_), .A2(new_n403_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n407_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT27), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n390_), .A2(new_n370_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n413_), .A2(new_n380_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n412_), .B1(new_n414_), .B2(new_n391_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n389_), .A2(new_n395_), .A3(new_n411_), .A4(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n358_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n380_), .A2(KEYINPUT32), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n411_), .B1(new_n387_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT96), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n413_), .A2(new_n422_), .A3(new_n419_), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT96), .B1(new_n376_), .B2(new_n420_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n421_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n376_), .A2(new_n381_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n396_), .A2(new_n401_), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n427_), .A2(new_n407_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n397_), .A2(new_n400_), .A3(new_n399_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT33), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n408_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n409_), .A2(KEYINPUT33), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n392_), .A2(new_n426_), .A3(new_n431_), .A4(new_n432_), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n425_), .A2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n355_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n435_));
  OR2_X1    g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n241_), .B1(new_n418_), .B2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G57gat), .B(G64gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT11), .ZN(new_n439_));
  XOR2_X1   g238(.A(G71gat), .B(G78gat), .Z(new_n440_));
  OR2_X1    g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n438_), .A2(KEYINPUT11), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(new_n440_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n441_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT68), .ZN(new_n445_));
  AND2_X1   g244(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n446_));
  NOR2_X1   g245(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n447_));
  OAI22_X1  g246(.A1(new_n446_), .A2(new_n447_), .B1(G99gat), .B2(G106gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G99gat), .A2(G106gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT6), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n451_), .A2(G99gat), .A3(G106gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(G99gat), .A2(G106gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n448_), .A2(new_n453_), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(G85gat), .ZN(new_n458_));
  INV_X1    g257(.A(G92gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G85gat), .A2(G92gat), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n457_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT8), .ZN(new_n464_));
  OR2_X1    g263(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n465_));
  INV_X1    g264(.A(G106gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT64), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT64), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n465_), .A2(new_n470_), .A3(new_n466_), .A4(new_n467_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n460_), .A2(KEYINPUT9), .A3(new_n461_), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n461_), .A2(KEYINPUT9), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n453_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  AOI22_X1  g274(.A1(new_n463_), .A2(new_n464_), .B1(new_n472_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT66), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT65), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT7), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n454_), .B1(new_n480_), .B2(new_n455_), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n454_), .A2(new_n455_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n477_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n448_), .A2(KEYINPUT66), .A3(new_n456_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(new_n484_), .A3(new_n453_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n462_), .A2(KEYINPUT8), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n476_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n445_), .A2(KEYINPUT12), .A3(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n476_), .A2(new_n488_), .A3(new_n444_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G230gat), .A2(G233gat), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n444_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n463_), .A2(new_n464_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n472_), .A2(new_n475_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n448_), .A2(new_n456_), .ZN(new_n498_));
  AOI22_X1  g297(.A1(new_n498_), .A2(new_n477_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n486_), .B1(new_n499_), .B2(new_n484_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n494_), .B1(new_n497_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT12), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT69), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n444_), .B1(new_n476_), .B2(new_n488_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT69), .ZN(new_n505_));
  NOR3_X1   g304(.A1(new_n504_), .A2(new_n505_), .A3(KEYINPUT12), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n490_), .B(new_n493_), .C1(new_n503_), .C2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT67), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n491_), .B(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n492_), .B1(new_n510_), .B2(new_n501_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n508_), .A2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G120gat), .B(G148gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT5), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G176gat), .B(G204gat), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n514_), .B(new_n515_), .Z(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(KEYINPUT70), .B1(new_n512_), .B2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n518_), .B1(new_n512_), .B2(new_n517_), .ZN(new_n519_));
  OAI211_X1 g318(.A(KEYINPUT70), .B(new_n516_), .C1(new_n508_), .C2(new_n511_), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n519_), .A2(KEYINPUT13), .A3(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(KEYINPUT13), .B1(new_n519_), .B2(new_n520_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n213_), .A2(KEYINPUT74), .ZN(new_n525_));
  INV_X1    g324(.A(G231gat), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n526_), .A2(new_n276_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT74), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n208_), .A2(new_n212_), .A3(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n525_), .A2(new_n527_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n527_), .B1(new_n525_), .B2(new_n529_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n445_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n532_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n445_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(new_n530_), .ZN(new_n536_));
  XOR2_X1   g335(.A(G127gat), .B(G155gat), .Z(new_n537_));
  XNOR2_X1  g336(.A(G183gat), .B(G211gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT17), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n533_), .A2(new_n536_), .A3(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT76), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n533_), .A2(new_n536_), .A3(KEYINPUT76), .A4(new_n543_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n531_), .A2(new_n532_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(new_n494_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n444_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n541_), .B(KEYINPUT17), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n550_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n548_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n489_), .A2(new_n217_), .ZN(new_n555_));
  XOR2_X1   g354(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n556_));
  NAND2_X1  g355(.A1(G232gat), .A2(G233gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  OAI221_X1 g357(.A(new_n555_), .B1(KEYINPUT35), .B2(new_n558_), .C1(new_n224_), .C2(new_n489_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(KEYINPUT35), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G190gat), .B(G218gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G134gat), .B(G162gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n564_), .A2(KEYINPUT36), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n561_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(KEYINPUT72), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT72), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n561_), .A2(new_n568_), .A3(new_n565_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n564_), .B(KEYINPUT36), .Z(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n561_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(KEYINPUT37), .B1(new_n570_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT37), .ZN(new_n576_));
  AOI211_X1 g375(.A(new_n576_), .B(new_n573_), .C1(new_n567_), .C2(new_n569_), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n554_), .A2(new_n575_), .A3(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n437_), .A2(new_n524_), .A3(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n411_), .B(KEYINPUT99), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NOR3_X1   g380(.A1(new_n579_), .A2(G1gat), .A3(new_n581_), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n582_), .A2(KEYINPUT38), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(KEYINPUT38), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n418_), .A2(new_n436_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT100), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n586_), .B1(new_n523_), .B2(new_n240_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n240_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n588_), .B(KEYINPUT100), .C1(new_n521_), .C2(new_n522_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n570_), .A2(new_n574_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT101), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n591_), .A2(new_n554_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n585_), .A2(new_n587_), .A3(new_n589_), .A4(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(G1gat), .B1(new_n593_), .B2(new_n411_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n583_), .A2(new_n584_), .A3(new_n594_), .ZN(G1324gat));
  NAND3_X1  g394(.A1(new_n389_), .A2(new_n415_), .A3(new_n395_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NOR3_X1   g396(.A1(new_n579_), .A2(G8gat), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT102), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT39), .ZN(new_n600_));
  OAI211_X1 g399(.A(G8gat), .B(new_n600_), .C1(new_n593_), .C2(new_n597_), .ZN(new_n601_));
  OR3_X1    g400(.A1(new_n601_), .A2(new_n599_), .A3(KEYINPUT39), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n601_), .B1(new_n599_), .B2(KEYINPUT39), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n598_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n604_), .B(new_n605_), .Z(G1325gat));
  NOR2_X1   g405(.A1(new_n349_), .A2(new_n350_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  OR3_X1    g407(.A1(new_n579_), .A2(G15gat), .A3(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n593_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(new_n607_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n611_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n612_));
  AOI21_X1  g411(.A(KEYINPUT41), .B1(new_n611_), .B2(G15gat), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n609_), .B1(new_n612_), .B2(new_n613_), .ZN(G1326gat));
  OR3_X1    g413(.A1(new_n579_), .A2(G22gat), .A3(new_n355_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n610_), .A2(new_n293_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n616_), .A2(G22gat), .A3(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n617_), .B1(new_n616_), .B2(G22gat), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n615_), .B1(new_n618_), .B2(new_n619_), .ZN(G1327gat));
  OR2_X1    g419(.A1(new_n575_), .A2(new_n577_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n416_), .B1(new_n351_), .B2(new_n357_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n434_), .A2(new_n435_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n621_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT43), .ZN(new_n628_));
  OAI221_X1 g427(.A(new_n621_), .B1(KEYINPUT105), .B2(new_n628_), .C1(new_n622_), .C2(new_n623_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n587_), .A2(new_n554_), .A3(new_n589_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(KEYINPUT44), .B1(new_n630_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT44), .ZN(new_n634_));
  AOI211_X1 g433(.A(new_n634_), .B(new_n631_), .C1(new_n627_), .C2(new_n629_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(new_n580_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(G29gat), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n591_), .A2(new_n554_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n639_), .A2(new_n523_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n437_), .A2(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n411_), .A2(G29gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT106), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n638_), .B1(new_n641_), .B2(new_n643_), .ZN(G1328gat));
  OR2_X1    g443(.A1(new_n596_), .A2(KEYINPUT108), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n596_), .A2(KEYINPUT108), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n641_), .A2(G36gat), .A3(new_n648_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT45), .Z(new_n650_));
  AND2_X1   g449(.A1(new_n627_), .A2(new_n629_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n634_), .B1(new_n651_), .B2(new_n631_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n630_), .A2(KEYINPUT44), .A3(new_n632_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n652_), .A2(KEYINPUT107), .A3(new_n596_), .A4(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(G36gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT107), .B1(new_n636_), .B2(new_n596_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n650_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n650_), .B(new_n658_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1329gat));
  NAND3_X1  g461(.A1(new_n636_), .A2(G43gat), .A3(new_n607_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n641_), .A2(new_n608_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n663_), .B1(G43gat), .B2(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g465(.A(new_n641_), .ZN(new_n667_));
  AOI21_X1  g466(.A(G50gat), .B1(new_n667_), .B2(new_n293_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n293_), .A2(G50gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n636_), .B2(new_n669_), .ZN(G1331gat));
  NAND4_X1  g469(.A1(new_n585_), .A2(new_n241_), .A3(new_n523_), .A4(new_n592_), .ZN(new_n671_));
  INV_X1    g470(.A(G57gat), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n671_), .A2(new_n672_), .A3(new_n411_), .ZN(new_n673_));
  AOI211_X1 g472(.A(new_n588_), .B(new_n524_), .C1(new_n418_), .C2(new_n436_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(new_n578_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n581_), .B1(new_n675_), .B2(KEYINPUT110), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n676_), .B1(KEYINPUT110), .B2(new_n675_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n673_), .B1(new_n677_), .B2(new_n672_), .ZN(G1332gat));
  OAI21_X1  g477(.A(G64gat), .B1(new_n671_), .B2(new_n648_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT48), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n648_), .A2(G64gat), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n680_), .B1(new_n675_), .B2(new_n681_), .ZN(G1333gat));
  OR3_X1    g481(.A1(new_n675_), .A2(G71gat), .A3(new_n608_), .ZN(new_n683_));
  OAI21_X1  g482(.A(G71gat), .B1(new_n671_), .B2(new_n608_), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n684_), .A2(KEYINPUT49), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n684_), .A2(KEYINPUT49), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n683_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT111), .Z(G1334gat));
  OAI21_X1  g488(.A(G78gat), .B1(new_n671_), .B2(new_n355_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT50), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n355_), .A2(G78gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(new_n675_), .B2(new_n692_), .ZN(G1335gat));
  INV_X1    g492(.A(new_n554_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n694_), .A2(new_n588_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(new_n523_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n651_), .A2(KEYINPUT112), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT112), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n630_), .A2(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n696_), .B1(new_n697_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G85gat), .B1(new_n701_), .B2(new_n411_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n639_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n674_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n705_), .A2(new_n458_), .A3(new_n580_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n702_), .A2(new_n706_), .ZN(G1336gat));
  OAI21_X1  g506(.A(G92gat), .B1(new_n701_), .B2(new_n648_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n705_), .A2(new_n459_), .A3(new_n596_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1337gat));
  INV_X1    g509(.A(G99gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n711_), .B1(new_n700_), .B2(new_n607_), .ZN(new_n712_));
  AND4_X1   g511(.A1(new_n607_), .A2(new_n705_), .A3(new_n465_), .A4(new_n467_), .ZN(new_n713_));
  OR3_X1    g512(.A1(new_n712_), .A2(KEYINPUT51), .A3(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(KEYINPUT51), .B1(new_n712_), .B2(new_n713_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1338gat));
  NAND3_X1  g515(.A1(new_n705_), .A2(new_n466_), .A3(new_n293_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n695_), .A2(new_n293_), .A3(new_n523_), .ZN(new_n718_));
  OAI21_X1  g517(.A(G106gat), .B1(new_n651_), .B2(new_n718_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n719_), .A2(KEYINPUT52), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(KEYINPUT52), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g522(.A(KEYINPUT59), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n524_), .A2(new_n241_), .A3(new_n578_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT54), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n725_), .B(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n591_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n218_), .A2(new_n219_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT116), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n221_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n731_), .B1(new_n730_), .B2(new_n729_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n229_), .B1(new_n232_), .B2(new_n221_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n231_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n519_), .A2(new_n520_), .A3(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n512_), .A2(new_n517_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n236_), .A2(new_n736_), .A3(new_n239_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT114), .ZN(new_n738_));
  AND2_X1   g537(.A1(G230gat), .A2(G233gat), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n501_), .A2(KEYINPUT69), .A3(new_n502_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n505_), .B1(new_n504_), .B2(KEYINPUT12), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n742_), .A2(new_n510_), .A3(new_n490_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n744_));
  AOI22_X1  g543(.A1(new_n739_), .A2(new_n743_), .B1(new_n507_), .B2(new_n744_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n742_), .A2(KEYINPUT55), .A3(new_n490_), .A4(new_n493_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n738_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n743_), .A2(new_n739_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n507_), .A2(new_n744_), .ZN(new_n749_));
  AND4_X1   g548(.A1(new_n738_), .A2(new_n748_), .A3(new_n746_), .A4(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n516_), .B1(new_n747_), .B2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT56), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n748_), .A2(new_n749_), .A3(new_n746_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT114), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n745_), .A2(new_n738_), .A3(new_n746_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n757_), .A2(KEYINPUT56), .A3(new_n516_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n737_), .B1(new_n753_), .B2(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n735_), .B1(new_n759_), .B2(KEYINPUT115), .ZN(new_n760_));
  INV_X1    g559(.A(new_n737_), .ZN(new_n761_));
  AOI21_X1  g560(.A(KEYINPUT56), .B1(new_n757_), .B2(new_n516_), .ZN(new_n762_));
  AOI211_X1 g561(.A(new_n752_), .B(new_n517_), .C1(new_n755_), .C2(new_n756_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n761_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT115), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n728_), .B1(new_n760_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT57), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  OAI211_X1 g568(.A(KEYINPUT57), .B(new_n728_), .C1(new_n760_), .C2(new_n766_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n734_), .A2(new_n736_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n771_), .B1(new_n762_), .B2(KEYINPUT117), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n753_), .A2(new_n773_), .A3(new_n758_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT58), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n772_), .A2(new_n774_), .A3(KEYINPUT58), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n777_), .A2(new_n621_), .A3(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n769_), .A2(new_n770_), .A3(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n727_), .B1(new_n780_), .B2(new_n554_), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n357_), .A2(new_n596_), .A3(new_n581_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n724_), .B1(new_n781_), .B2(new_n783_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n778_), .A2(new_n621_), .ZN(new_n785_));
  AOI22_X1  g584(.A1(new_n767_), .A2(new_n768_), .B1(new_n785_), .B2(new_n777_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n694_), .B1(new_n786_), .B2(new_n770_), .ZN(new_n787_));
  OAI211_X1 g586(.A(KEYINPUT59), .B(new_n782_), .C1(new_n787_), .C2(new_n727_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n784_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(G113gat), .B1(new_n790_), .B2(new_n241_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n735_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n759_), .A2(KEYINPUT115), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n591_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n779_), .B1(new_n795_), .B2(KEYINPUT57), .ZN(new_n796_));
  INV_X1    g595(.A(new_n770_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n554_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n727_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n783_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  OR2_X1    g600(.A1(new_n240_), .A2(G113gat), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n791_), .B1(new_n801_), .B2(new_n802_), .ZN(G1340gat));
  INV_X1    g602(.A(G120gat), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n789_), .B2(new_n523_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n798_), .A2(new_n799_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT60), .ZN(new_n807_));
  AOI21_X1  g606(.A(G120gat), .B1(new_n523_), .B2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n808_), .B1(new_n807_), .B2(G120gat), .ZN(new_n809_));
  AND4_X1   g608(.A1(KEYINPUT118), .A2(new_n806_), .A3(new_n782_), .A4(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT118), .B1(new_n800_), .B2(new_n809_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(KEYINPUT119), .B1(new_n805_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n524_), .B1(new_n784_), .B2(new_n788_), .ZN(new_n815_));
  OAI221_X1 g614(.A(new_n814_), .B1(new_n810_), .B2(new_n811_), .C1(new_n815_), .C2(new_n804_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n813_), .A2(new_n816_), .ZN(G1341gat));
  OAI21_X1  g616(.A(G127gat), .B1(new_n790_), .B2(new_n554_), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n554_), .A2(G127gat), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n818_), .B1(new_n801_), .B2(new_n819_), .ZN(G1342gat));
  INV_X1    g619(.A(G134gat), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n821_), .B1(new_n801_), .B2(new_n728_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT120), .ZN(new_n823_));
  OR2_X1    g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n823_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n621_), .A2(G134gat), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(KEYINPUT121), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n824_), .A2(new_n825_), .B1(new_n789_), .B2(new_n827_), .ZN(G1343gat));
  NOR3_X1   g627(.A1(new_n647_), .A2(new_n351_), .A3(new_n581_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n806_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n588_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n523_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g634(.A1(new_n830_), .A2(new_n554_), .ZN(new_n836_));
  XOR2_X1   g635(.A(KEYINPUT61), .B(G155gat), .Z(new_n837_));
  XNOR2_X1  g636(.A(new_n836_), .B(new_n837_), .ZN(G1346gat));
  NOR2_X1   g637(.A1(new_n830_), .A2(new_n728_), .ZN(new_n839_));
  OR3_X1    g638(.A1(new_n839_), .A2(KEYINPUT122), .A3(G162gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT122), .B1(new_n839_), .B2(G162gat), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n621_), .A2(G162gat), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(KEYINPUT123), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n840_), .A2(new_n841_), .B1(new_n831_), .B2(new_n843_), .ZN(G1347gat));
  NOR2_X1   g643(.A1(new_n781_), .A2(new_n293_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n647_), .A2(new_n607_), .A3(new_n581_), .ZN(new_n846_));
  XOR2_X1   g645(.A(new_n846_), .B(KEYINPUT124), .Z(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(G169gat), .B1(new_n848_), .B2(new_n240_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT62), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n845_), .A2(new_n847_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n852_), .A2(new_n361_), .A3(new_n588_), .ZN(new_n853_));
  OAI211_X1 g652(.A(KEYINPUT62), .B(G169gat), .C1(new_n848_), .C2(new_n240_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n851_), .A2(new_n853_), .A3(new_n854_), .ZN(G1348gat));
  NAND2_X1  g654(.A1(new_n852_), .A2(new_n523_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n845_), .A2(KEYINPUT125), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT125), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n781_), .B2(new_n293_), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n847_), .A2(G176gat), .A3(new_n523_), .ZN(new_n861_));
  AOI22_X1  g660(.A1(new_n309_), .A2(new_n856_), .B1(new_n860_), .B2(new_n861_), .ZN(G1349gat));
  NAND4_X1  g661(.A1(new_n857_), .A2(new_n694_), .A3(new_n847_), .A4(new_n859_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n694_), .A2(new_n299_), .ZN(new_n864_));
  AOI22_X1  g663(.A1(new_n863_), .A2(new_n315_), .B1(new_n852_), .B2(new_n864_), .ZN(G1350gat));
  NAND2_X1  g664(.A1(new_n852_), .A2(new_n621_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(G190gat), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n728_), .A2(new_n300_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n848_), .B2(new_n868_), .ZN(G1351gat));
  INV_X1    g668(.A(new_n411_), .ZN(new_n870_));
  NOR4_X1   g669(.A1(new_n781_), .A2(new_n351_), .A3(new_n870_), .A4(new_n648_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n588_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n523_), .ZN(new_n874_));
  MUX2_X1   g673(.A(new_n245_), .B(G204gat), .S(new_n874_), .Z(G1353gat));
  AOI21_X1  g674(.A(new_n554_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n876_));
  XOR2_X1   g675(.A(new_n876_), .B(KEYINPUT126), .Z(new_n877_));
  NOR2_X1   g676(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(KEYINPUT127), .B2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n871_), .A2(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n878_), .A2(KEYINPUT127), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n880_), .B(new_n881_), .ZN(G1354gat));
  INV_X1    g681(.A(G218gat), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n871_), .A2(new_n883_), .A3(new_n591_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n871_), .A2(new_n621_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(new_n883_), .ZN(G1355gat));
endmodule


