//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 1 0 1 0 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n785_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n947_,
    new_n948_, new_n950_, new_n951_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n960_, new_n961_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n972_, new_n973_, new_n974_, new_n975_;
  INV_X1    g000(.A(KEYINPUT20), .ZN(new_n202_));
  NOR3_X1   g001(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206_));
  AOI21_X1  g005(.A(new_n203_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT23), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(G183gat), .A3(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT26), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT26), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(G190gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT25), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(G183gat), .ZN(new_n218_));
  INV_X1    g017(.A(G183gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT25), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n214_), .A2(new_n216_), .A3(new_n218_), .A4(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n207_), .A2(new_n212_), .A3(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT89), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n208_), .A2(new_n210_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n219_), .A2(new_n213_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT90), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT90), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n210_), .B1(G183gat), .B2(G190gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n208_), .A2(KEYINPUT23), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n229_), .B(new_n225_), .C1(new_n230_), .C2(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(G169gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n228_), .A2(new_n232_), .A3(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT89), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n207_), .A2(new_n236_), .A3(new_n212_), .A4(new_n221_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n223_), .A2(new_n235_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(G197gat), .ZN(new_n239_));
  INV_X1    g038(.A(G204gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G197gat), .A2(G204gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n241_), .A2(KEYINPUT21), .A3(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G211gat), .B(G218gat), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT21), .ZN(new_n246_));
  INV_X1    g045(.A(new_n242_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(G197gat), .A2(G204gat), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n246_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n245_), .A2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n202_), .B1(new_n238_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n251_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT83), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n212_), .A2(new_n254_), .A3(new_n225_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n227_), .A2(KEYINPUT83), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(new_n256_), .A3(new_n234_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT26), .B(G190gat), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT25), .B1(new_n219_), .B2(KEYINPUT82), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n258_), .B(new_n259_), .C1(KEYINPUT82), .C2(new_n218_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n260_), .A2(new_n212_), .A3(new_n207_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n253_), .A2(new_n257_), .A3(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n252_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G226gat), .A2(G233gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT19), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(G8gat), .B(G36gat), .Z(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT18), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G64gat), .B(G92gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n253_), .A2(new_n223_), .A3(new_n235_), .A4(new_n237_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n257_), .A2(new_n261_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n251_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n265_), .A2(new_n202_), .ZN(new_n274_));
  AND3_X1   g073(.A1(new_n271_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n266_), .A2(new_n270_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n270_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n265_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n279_), .B1(new_n252_), .B2(new_n262_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n278_), .B1(new_n280_), .B2(new_n275_), .ZN(new_n281_));
  AOI21_X1  g080(.A(KEYINPUT27), .B1(new_n277_), .B2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n222_), .A2(new_n250_), .A3(new_n245_), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n228_), .A2(new_n232_), .A3(new_n234_), .ZN(new_n284_));
  OAI211_X1 g083(.A(KEYINPUT95), .B(KEYINPUT20), .C1(new_n283_), .C2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n273_), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n235_), .A2(new_n250_), .A3(new_n245_), .A4(new_n222_), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT95), .B1(new_n287_), .B2(KEYINPUT20), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n265_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n252_), .A2(new_n279_), .A3(new_n262_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n270_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  OAI211_X1 g090(.A(KEYINPUT27), .B(new_n277_), .C1(new_n291_), .C2(KEYINPUT96), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(KEYINPUT96), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n282_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT97), .ZN(new_n296_));
  INV_X1    g095(.A(G228gat), .ZN(new_n297_));
  INV_X1    g096(.A(G233gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n251_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT86), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n300_), .B1(new_n301_), .B2(KEYINPUT1), .ZN(new_n302_));
  OR2_X1    g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT1), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n304_), .A2(KEYINPUT86), .A3(G155gat), .A4(G162gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n301_), .A2(KEYINPUT1), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n302_), .A2(new_n303_), .A3(new_n305_), .A4(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(G141gat), .ZN(new_n308_));
  INV_X1    g107(.A(G148gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n308_), .A2(new_n309_), .A3(KEYINPUT85), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT85), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n311_), .B1(G141gat), .B2(G148gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G141gat), .A2(G148gat), .ZN(new_n313_));
  AND3_X1   g112(.A1(new_n310_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT3), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n315_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT2), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n313_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n316_), .A2(new_n318_), .A3(new_n319_), .A4(new_n320_), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n303_), .A2(new_n301_), .ZN(new_n322_));
  AOI22_X1  g121(.A1(new_n307_), .A2(new_n314_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT29), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n299_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT87), .B(KEYINPUT29), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n251_), .B1(new_n323_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT88), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n297_), .A2(new_n298_), .ZN(new_n331_));
  AND3_X1   g130(.A1(new_n329_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n330_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n327_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(G78gat), .B(G106gat), .Z(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n329_), .A2(new_n331_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT88), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n329_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n335_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(new_n341_), .A3(new_n327_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n307_), .A2(new_n314_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n321_), .A2(new_n322_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT28), .B1(new_n345_), .B2(KEYINPUT29), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT28), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n323_), .A2(new_n347_), .A3(new_n324_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G22gat), .B(G50gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  AND3_X1   g149(.A1(new_n346_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n350_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n336_), .A2(new_n342_), .A3(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n353_), .B1(new_n336_), .B2(new_n342_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT84), .B(G43gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT31), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(KEYINPUT30), .B1(new_n257_), .B2(new_n261_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(G71gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G227gat), .A2(G233gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(G15gat), .ZN(new_n364_));
  INV_X1    g163(.A(G15gat), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(G227gat), .A3(G233gat), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n362_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n364_), .A2(new_n366_), .A3(new_n362_), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n368_), .A2(G99gat), .A3(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(G99gat), .B1(new_n368_), .B2(new_n369_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n257_), .A2(new_n261_), .A3(KEYINPUT30), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n361_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n370_), .A2(new_n371_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n257_), .A2(new_n261_), .A3(KEYINPUT30), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n375_), .B1(new_n376_), .B2(new_n360_), .ZN(new_n377_));
  INV_X1    g176(.A(G134gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(G127gat), .ZN(new_n379_));
  INV_X1    g178(.A(G127gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(G134gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(G120gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(G113gat), .ZN(new_n384_));
  INV_X1    g183(.A(G113gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(G120gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n382_), .A2(new_n387_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n379_), .A2(new_n381_), .A3(new_n384_), .A4(new_n386_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  AND3_X1   g189(.A1(new_n374_), .A2(new_n377_), .A3(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n390_), .B1(new_n374_), .B2(new_n377_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n359_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n374_), .A2(new_n377_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n388_), .A2(new_n389_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n374_), .A2(new_n377_), .A3(new_n390_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n396_), .A2(new_n358_), .A3(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G225gat), .A2(G233gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT91), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n323_), .A2(new_n390_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT4), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n401_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n345_), .A2(new_n395_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n323_), .A2(new_n390_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(KEYINPUT4), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n404_), .A2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n323_), .B(new_n395_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(new_n401_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G1gat), .B(G29gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G57gat), .B(G85gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(KEYINPUT92), .B(KEYINPUT0), .Z(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n408_), .A2(new_n410_), .A3(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n416_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n393_), .A2(new_n398_), .A3(new_n419_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n295_), .A2(new_n296_), .A3(new_n356_), .A4(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n289_), .A2(new_n290_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n278_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT96), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NOR3_X1   g224(.A1(new_n280_), .A2(new_n278_), .A3(new_n275_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT27), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n425_), .A2(new_n294_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n282_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n429_), .A2(new_n356_), .A3(new_n430_), .A4(new_n420_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT97), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n270_), .A2(KEYINPUT32), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n422_), .A2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n266_), .A2(new_n433_), .A3(new_n276_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n408_), .A2(new_n410_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(new_n415_), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n407_), .A2(new_n404_), .B1(new_n409_), .B2(new_n401_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n416_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n435_), .A2(new_n436_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT33), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n443_), .B1(new_n439_), .B2(new_n416_), .ZN(new_n444_));
  AND4_X1   g243(.A1(new_n443_), .A2(new_n408_), .A3(new_n410_), .A4(new_n416_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n277_), .B(new_n281_), .C1(new_n444_), .C2(new_n445_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n407_), .B(new_n401_), .C1(KEYINPUT4), .C2(new_n405_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n405_), .A2(new_n406_), .A3(new_n400_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT93), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n448_), .A2(new_n449_), .A3(new_n415_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n449_), .B1(new_n448_), .B2(new_n415_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n447_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT94), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT94), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n447_), .B(new_n454_), .C1(new_n450_), .C2(new_n451_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n442_), .B1(new_n446_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n356_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n353_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n341_), .B1(new_n340_), .B2(new_n327_), .ZN(new_n460_));
  AOI211_X1 g259(.A(new_n335_), .B(new_n326_), .C1(new_n338_), .C2(new_n339_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n459_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n336_), .A2(new_n342_), .A3(new_n353_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n441_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n429_), .A2(new_n464_), .A3(new_n430_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n458_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n393_), .A2(new_n398_), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n421_), .A2(new_n432_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(G85gat), .ZN(new_n469_));
  INV_X1    g268(.A(G92gat), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(new_n470_), .A3(KEYINPUT9), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n471_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n472_));
  XOR2_X1   g271(.A(KEYINPUT65), .B(KEYINPUT9), .Z(new_n473_));
  OR2_X1    g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G99gat), .A2(G106gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT6), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT6), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n477_), .A2(G99gat), .A3(G106gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n472_), .A2(new_n473_), .ZN(new_n480_));
  XOR2_X1   g279(.A(KEYINPUT10), .B(G99gat), .Z(new_n481_));
  INV_X1    g280(.A(G106gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n474_), .A2(new_n479_), .A3(new_n480_), .A4(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G43gat), .B(G50gat), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(G36gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(G29gat), .ZN(new_n488_));
  INV_X1    g287(.A(G29gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(G36gat), .ZN(new_n490_));
  AND3_X1   g289(.A1(new_n488_), .A2(new_n490_), .A3(KEYINPUT68), .ZN(new_n491_));
  AOI21_X1  g290(.A(KEYINPUT68), .B1(new_n488_), .B2(new_n490_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n486_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT68), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n489_), .A2(G36gat), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n487_), .A2(G29gat), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n494_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n488_), .A2(new_n490_), .A3(KEYINPUT68), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n497_), .A2(new_n498_), .A3(new_n485_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n493_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT66), .ZN(new_n501_));
  NOR2_X1   g300(.A1(G99gat), .A2(G106gat), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT7), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n501_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  OAI211_X1 g303(.A(KEYINPUT66), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  AOI22_X1  g305(.A1(new_n476_), .A2(new_n478_), .B1(new_n503_), .B2(new_n502_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT8), .ZN(new_n509_));
  XOR2_X1   g308(.A(G85gat), .B(G92gat), .Z(new_n510_));
  NAND3_X1  g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n509_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n484_), .B(new_n500_), .C1(new_n512_), .C2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT69), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n508_), .A2(new_n510_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT8), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(new_n511_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT69), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n518_), .A2(new_n519_), .A3(new_n500_), .A4(new_n484_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n484_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n493_), .A2(new_n499_), .A3(KEYINPUT15), .ZN(new_n522_));
  AOI21_X1  g321(.A(KEYINPUT15), .B1(new_n493_), .B2(new_n499_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n515_), .A2(new_n520_), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT35), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT70), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n515_), .A2(new_n525_), .A3(new_n520_), .A4(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G232gat), .A2(G233gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n528_), .A2(new_n530_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT71), .ZN(new_n535_));
  AOI22_X1  g334(.A1(new_n514_), .A2(KEYINPUT69), .B1(new_n521_), .B2(new_n524_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n533_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n536_), .A2(new_n529_), .A3(new_n520_), .A4(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G190gat), .B(G218gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G134gat), .B(G162gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n541_), .A2(KEYINPUT36), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n534_), .A2(new_n535_), .A3(new_n538_), .A4(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n530_), .A2(new_n533_), .ZN(new_n544_));
  AOI21_X1  g343(.A(KEYINPUT35), .B1(new_n536_), .B2(new_n520_), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n538_), .B(new_n542_), .C1(new_n544_), .C2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT71), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n541_), .B(KEYINPUT36), .Z(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n549_), .B1(new_n534_), .B2(new_n538_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n543_), .B1(new_n547_), .B2(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n468_), .A2(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(G127gat), .B(G155gat), .Z(new_n553_));
  XNOR2_X1  g352(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G183gat), .B(G211gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT17), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT11), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G71gat), .B(G78gat), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G57gat), .B(G64gat), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT67), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n564_), .ZN(new_n566_));
  AOI211_X1 g365(.A(new_n560_), .B(new_n562_), .C1(new_n565_), .C2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n565_), .A2(new_n560_), .A3(new_n566_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n563_), .B(new_n564_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n561_), .B1(new_n569_), .B2(KEYINPUT11), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n567_), .B1(new_n568_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(G231gat), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n572_), .A2(new_n298_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n569_), .A2(KEYINPUT11), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n575_), .A2(new_n562_), .A3(new_n568_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n569_), .A2(KEYINPUT11), .A3(new_n561_), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n576_), .A2(new_n577_), .A3(new_n573_), .ZN(new_n578_));
  OAI21_X1  g377(.A(KEYINPUT73), .B1(new_n574_), .B2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n577_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n580_), .B1(new_n572_), .B2(new_n298_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT73), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n571_), .A2(new_n573_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n581_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G15gat), .B(G22gat), .ZN(new_n585_));
  INV_X1    g384(.A(G1gat), .ZN(new_n586_));
  INV_X1    g385(.A(G8gat), .ZN(new_n587_));
  OAI21_X1  g386(.A(KEYINPUT14), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n585_), .A2(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(G1gat), .B(G8gat), .Z(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  AND3_X1   g390(.A1(new_n579_), .A2(new_n584_), .A3(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n591_), .B1(new_n579_), .B2(new_n584_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n559_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT75), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  OAI211_X1 g395(.A(KEYINPUT75), .B(new_n559_), .C1(new_n592_), .C2(new_n593_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n557_), .B(new_n558_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n592_), .A2(new_n593_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n598_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G230gat), .A2(G233gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT64), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n580_), .A2(new_n518_), .A3(new_n484_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n571_), .A2(new_n521_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n607_), .A2(new_n608_), .A3(KEYINPUT12), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT12), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n571_), .A2(new_n521_), .A3(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n606_), .B1(new_n609_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n607_), .A2(new_n608_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(new_n606_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G120gat), .B(G148gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT5), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G176gat), .B(G204gat), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n618_), .B(new_n619_), .Z(new_n620_));
  NAND2_X1  g419(.A1(new_n616_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n620_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n613_), .A2(new_n615_), .A3(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT13), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n591_), .A2(new_n500_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n627_), .A2(KEYINPUT77), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT77), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n629_), .B1(new_n591_), .B2(new_n500_), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(G229gat), .A2(G233gat), .ZN(new_n632_));
  OR3_X1    g431(.A1(new_n522_), .A2(new_n523_), .A3(new_n591_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n631_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT79), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n591_), .A2(new_n500_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n636_), .B1(new_n628_), .B2(new_n630_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(KEYINPUT78), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT78), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n636_), .B(new_n639_), .C1(new_n628_), .C2(new_n630_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n632_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n635_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  AOI211_X1 g442(.A(KEYINPUT79), .B(new_n632_), .C1(new_n638_), .C2(new_n640_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n634_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(G113gat), .B(G141gat), .Z(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT80), .ZN(new_n647_));
  XNOR2_X1  g446(.A(G169gat), .B(G197gat), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n647_), .B(new_n648_), .Z(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n645_), .A2(new_n650_), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n634_), .B(new_n649_), .C1(new_n643_), .C2(new_n644_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n626_), .A2(new_n654_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n552_), .A2(new_n603_), .A3(new_n655_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n656_), .A2(new_n441_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n657_), .A2(new_n586_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT38), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT76), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n660_), .B1(new_n598_), .B2(new_n601_), .ZN(new_n661_));
  AOI211_X1 g460(.A(KEYINPUT76), .B(new_n600_), .C1(new_n596_), .C2(new_n597_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n624_), .B(KEYINPUT13), .ZN(new_n664_));
  OAI21_X1  g463(.A(KEYINPUT37), .B1(new_n550_), .B2(KEYINPUT72), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n551_), .B(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n663_), .A2(new_n664_), .A3(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n653_), .B(KEYINPUT81), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n669_), .A2(new_n468_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n672_), .A2(new_n586_), .A3(new_n441_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n658_), .B1(new_n659_), .B2(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n674_), .B1(new_n659_), .B2(new_n673_), .ZN(G1324gat));
  INV_X1    g474(.A(new_n294_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n430_), .B1(new_n292_), .B2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n656_), .A2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(KEYINPUT98), .B1(new_n678_), .B2(G8gat), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT39), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n672_), .A2(new_n587_), .A3(new_n677_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n678_), .A2(KEYINPUT98), .A3(G8gat), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n679_), .A2(new_n680_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n683_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT40), .ZN(G1325gat));
  INV_X1    g486(.A(new_n467_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n365_), .B1(new_n656_), .B2(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT41), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n672_), .A2(new_n365_), .A3(new_n688_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1326gat));
  INV_X1    g491(.A(G22gat), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n462_), .A2(new_n463_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n656_), .B2(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(KEYINPUT99), .B(KEYINPUT42), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n695_), .B(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n356_), .A2(G22gat), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT100), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n697_), .B1(new_n671_), .B2(new_n699_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT101), .Z(G1327gat));
  OAI21_X1  g500(.A(KEYINPUT43), .B1(new_n468_), .B2(new_n666_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n703_));
  OAI211_X1 g502(.A(new_n665_), .B(new_n543_), .C1(new_n550_), .C2(new_n547_), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n550_), .A2(KEYINPUT72), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n551_), .A2(new_n705_), .A3(KEYINPUT37), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n431_), .B(new_n296_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n688_), .B1(new_n458_), .B2(new_n465_), .ZN(new_n709_));
  OAI211_X1 g508(.A(new_n703_), .B(new_n707_), .C1(new_n708_), .C2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n702_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n663_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(new_n712_), .A3(new_n655_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(KEYINPUT102), .A2(KEYINPUT44), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n711_), .A2(new_n712_), .A3(new_n655_), .A4(new_n714_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n489_), .B1(new_n718_), .B2(new_n441_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n551_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n663_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(new_n664_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n670_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n724_), .A2(G29gat), .A3(new_n419_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n719_), .A2(new_n725_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT103), .Z(G1328gat));
  NOR2_X1   g526(.A1(new_n295_), .A2(G36gat), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n670_), .A2(new_n721_), .A3(new_n664_), .A4(new_n728_), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n729_), .A2(KEYINPUT104), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(KEYINPUT104), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n730_), .A2(KEYINPUT45), .A3(new_n731_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n295_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n734_), .B(new_n735_), .C1(new_n487_), .C2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT46), .ZN(G1329gat));
  NOR3_X1   g539(.A1(new_n724_), .A2(G43gat), .A3(new_n467_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n718_), .A2(new_n688_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n742_), .B2(G43gat), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g543(.A(new_n724_), .ZN(new_n745_));
  AOI21_X1  g544(.A(G50gat), .B1(new_n745_), .B2(new_n694_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n694_), .A2(G50gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n718_), .B2(new_n747_), .ZN(G1331gat));
  NOR2_X1   g547(.A1(new_n712_), .A2(new_n707_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n626_), .A2(new_n654_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n750_), .A2(new_n468_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n419_), .B1(new_n752_), .B2(KEYINPUT106), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n753_), .B1(KEYINPUT106), .B2(new_n752_), .ZN(new_n754_));
  INV_X1    g553(.A(G57gat), .ZN(new_n755_));
  AND4_X1   g554(.A1(new_n669_), .A2(new_n552_), .A3(new_n626_), .A4(new_n663_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n419_), .A2(new_n755_), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n754_), .A2(new_n755_), .B1(new_n756_), .B2(new_n757_), .ZN(G1332gat));
  INV_X1    g557(.A(G64gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n756_), .B2(new_n677_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT48), .Z(new_n761_));
  INV_X1    g560(.A(new_n752_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n762_), .A2(new_n759_), .A3(new_n677_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1333gat));
  AOI21_X1  g563(.A(new_n362_), .B1(new_n756_), .B2(new_n688_), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT49), .Z(new_n766_));
  NAND3_X1  g565(.A1(new_n762_), .A2(new_n362_), .A3(new_n688_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(G1334gat));
  INV_X1    g567(.A(G78gat), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n769_), .B1(new_n756_), .B2(new_n694_), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n770_), .B(KEYINPUT50), .Z(new_n771_));
  NAND3_X1  g570(.A1(new_n762_), .A2(new_n769_), .A3(new_n694_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT107), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n773_), .B(new_n774_), .ZN(G1335gat));
  AND2_X1   g574(.A1(new_n751_), .A2(new_n721_), .ZN(new_n776_));
  AOI21_X1  g575(.A(G85gat), .B1(new_n776_), .B2(new_n441_), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n626_), .B(new_n654_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n778_), .B1(new_n702_), .B2(new_n710_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n441_), .A2(G85gat), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT108), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n777_), .B1(new_n779_), .B2(new_n781_), .ZN(G1336gat));
  INV_X1    g581(.A(new_n779_), .ZN(new_n783_));
  OAI21_X1  g582(.A(G92gat), .B1(new_n783_), .B2(new_n295_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n776_), .A2(new_n470_), .A3(new_n677_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(G1337gat));
  NAND3_X1  g585(.A1(new_n776_), .A2(new_n688_), .A3(new_n481_), .ZN(new_n787_));
  XOR2_X1   g586(.A(new_n787_), .B(KEYINPUT109), .Z(new_n788_));
  OAI21_X1  g587(.A(G99gat), .B1(new_n783_), .B2(new_n467_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT110), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n791_));
  AOI22_X1  g590(.A1(new_n788_), .A2(new_n789_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n790_), .A2(new_n791_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n792_), .B(new_n793_), .ZN(G1338gat));
  INV_X1    g593(.A(KEYINPUT113), .ZN(new_n795_));
  INV_X1    g594(.A(new_n778_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n421_), .A2(new_n432_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n466_), .A2(new_n467_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n703_), .B1(new_n799_), .B2(new_n707_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n468_), .A2(new_n666_), .A3(KEYINPUT43), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n694_), .B(new_n796_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT111), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n779_), .A2(new_n804_), .A3(new_n694_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n482_), .B1(new_n803_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n795_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  AND4_X1   g607(.A1(new_n804_), .A2(new_n711_), .A3(new_n694_), .A4(new_n796_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n804_), .B1(new_n779_), .B2(new_n694_), .ZN(new_n810_));
  OAI21_X1  g609(.A(G106gat), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n811_), .A2(KEYINPUT113), .A3(KEYINPUT52), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n482_), .A2(KEYINPUT52), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT112), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  OAI211_X1 g615(.A(KEYINPUT112), .B(new_n813_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n808_), .A2(new_n812_), .A3(new_n816_), .A4(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n776_), .A2(new_n482_), .A3(new_n694_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT53), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n818_), .A2(new_n822_), .A3(new_n819_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(G1339gat));
  NOR2_X1   g623(.A1(new_n677_), .A2(new_n694_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n467_), .A2(new_n419_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n609_), .A2(new_n606_), .A3(new_n611_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n612_), .B1(new_n828_), .B2(KEYINPUT55), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830_));
  AOI211_X1 g629(.A(new_n830_), .B(new_n606_), .C1(new_n609_), .C2(new_n611_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n620_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT56), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(KEYINPUT114), .A3(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n623_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n832_), .A2(new_n833_), .ZN(new_n837_));
  OAI211_X1 g636(.A(KEYINPUT56), .B(new_n620_), .C1(new_n829_), .C2(new_n831_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n834_), .B(new_n836_), .C1(new_n839_), .C2(KEYINPUT114), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n641_), .A2(new_n632_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n631_), .A2(new_n642_), .A3(new_n633_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n841_), .A2(new_n650_), .A3(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n624_), .A2(new_n652_), .A3(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n551_), .B1(new_n840_), .B2(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(KEYINPUT116), .A2(KEYINPUT58), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n652_), .A2(new_n848_), .A3(new_n623_), .A4(new_n843_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n839_), .A2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n652_), .A2(new_n623_), .A3(new_n843_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(KEYINPUT115), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n847_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n839_), .A2(new_n852_), .A3(new_n847_), .A4(new_n849_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n707_), .ZN(new_n855_));
  OAI22_X1  g654(.A1(new_n845_), .A2(KEYINPUT57), .B1(new_n853_), .B2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n837_), .A2(new_n857_), .A3(new_n838_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n836_), .A2(new_n834_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n844_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n720_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n602_), .B1(new_n856_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n668_), .A2(new_n865_), .A3(new_n669_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n669_), .ZN(new_n867_));
  OAI21_X1  g666(.A(KEYINPUT54), .B1(new_n667_), .B2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n827_), .B1(new_n864_), .B2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT59), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n854_), .A2(new_n707_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n839_), .A2(new_n849_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n852_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n846_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  AOI22_X1  g674(.A1(new_n861_), .A2(new_n862_), .B1(new_n872_), .B2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n845_), .A2(KEYINPUT57), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n663_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n866_), .A2(new_n868_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n827_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n871_), .ZN(new_n882_));
  OAI22_X1  g681(.A1(new_n870_), .A2(new_n871_), .B1(new_n880_), .B2(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(G113gat), .B1(new_n883_), .B2(new_n669_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n870_), .A2(new_n385_), .A3(new_n653_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1340gat));
  OAI21_X1  g685(.A(G120gat), .B1(new_n883_), .B2(new_n664_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n603_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n881_), .B1(new_n888_), .B2(new_n879_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n383_), .B1(new_n664_), .B2(KEYINPUT60), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n890_), .B1(KEYINPUT60), .B2(new_n383_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n887_), .B1(new_n889_), .B2(new_n891_), .ZN(G1341gat));
  OAI21_X1  g691(.A(new_n380_), .B1(new_n889_), .B2(new_n712_), .ZN(new_n893_));
  OR2_X1    g692(.A1(new_n893_), .A2(KEYINPUT117), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(KEYINPUT117), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n712_), .B1(new_n856_), .B2(new_n863_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n882_), .B1(new_n896_), .B2(new_n869_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n897_), .B1(new_n889_), .B2(KEYINPUT59), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n603_), .A2(G127gat), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(KEYINPUT118), .ZN(new_n900_));
  AOI22_X1  g699(.A1(new_n894_), .A2(new_n895_), .B1(new_n898_), .B2(new_n900_), .ZN(G1342gat));
  AOI21_X1  g700(.A(new_n378_), .B1(new_n898_), .B2(new_n707_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n889_), .A2(G134gat), .A3(new_n720_), .ZN(new_n903_));
  OAI21_X1  g702(.A(KEYINPUT119), .B1(new_n902_), .B2(new_n903_), .ZN(new_n904_));
  OAI21_X1  g703(.A(G134gat), .B1(new_n883_), .B2(new_n666_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n906_));
  INV_X1    g705(.A(new_n903_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n905_), .A2(new_n906_), .A3(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n904_), .A2(new_n908_), .ZN(G1343gat));
  NAND2_X1  g708(.A1(new_n864_), .A2(new_n869_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n694_), .A2(new_n441_), .A3(new_n467_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n677_), .A2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n910_), .A2(new_n912_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(new_n654_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(KEYINPUT120), .B(G141gat), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n914_), .B(new_n915_), .ZN(G1344gat));
  NOR2_X1   g715(.A1(new_n913_), .A2(new_n664_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(KEYINPUT121), .B(G148gat), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n917_), .B(new_n918_), .ZN(G1345gat));
  INV_X1    g718(.A(KEYINPUT122), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n920_), .B1(new_n913_), .B2(new_n712_), .ZN(new_n921_));
  NAND4_X1  g720(.A1(new_n910_), .A2(KEYINPUT122), .A3(new_n663_), .A4(new_n912_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(KEYINPUT61), .B(G155gat), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n923_), .B(new_n924_), .ZN(G1346gat));
  OAI21_X1  g724(.A(G162gat), .B1(new_n913_), .B2(new_n666_), .ZN(new_n926_));
  OR2_X1    g725(.A1(new_n720_), .A2(G162gat), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n913_), .B2(new_n927_), .ZN(G1347gat));
  INV_X1    g727(.A(G169gat), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n677_), .A2(new_n420_), .ZN(new_n930_));
  AOI211_X1 g729(.A(new_n694_), .B(new_n930_), .C1(new_n896_), .C2(new_n869_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n929_), .B1(new_n931_), .B2(new_n653_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT62), .ZN(new_n933_));
  AND2_X1   g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n932_), .A2(new_n933_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n931_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(KEYINPUT22), .B(G169gat), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n653_), .A2(new_n937_), .ZN(new_n938_));
  XOR2_X1   g737(.A(new_n938_), .B(KEYINPUT123), .Z(new_n939_));
  OAI22_X1  g738(.A1(new_n934_), .A2(new_n935_), .B1(new_n936_), .B2(new_n939_), .ZN(G1348gat));
  AOI21_X1  g739(.A(G176gat), .B1(new_n931_), .B2(new_n626_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n910_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n942_), .A2(new_n694_), .ZN(new_n943_));
  INV_X1    g742(.A(G176gat), .ZN(new_n944_));
  NOR3_X1   g743(.A1(new_n664_), .A2(new_n944_), .A3(new_n930_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n941_), .B1(new_n943_), .B2(new_n945_), .ZN(G1349gat));
  NAND4_X1  g745(.A1(new_n943_), .A2(new_n677_), .A3(new_n420_), .A4(new_n663_), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n602_), .B1(new_n218_), .B2(new_n220_), .ZN(new_n948_));
  AOI22_X1  g747(.A1(new_n947_), .A2(new_n219_), .B1(new_n931_), .B2(new_n948_), .ZN(G1350gat));
  OAI21_X1  g748(.A(G190gat), .B1(new_n936_), .B2(new_n666_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n931_), .A2(new_n258_), .A3(new_n551_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n950_), .A2(new_n951_), .ZN(G1351gat));
  NAND2_X1  g751(.A1(new_n464_), .A2(new_n467_), .ZN(new_n953_));
  OR2_X1    g752(.A1(new_n953_), .A2(KEYINPUT124), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n953_), .A2(KEYINPUT124), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n954_), .A2(new_n677_), .A3(new_n955_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n942_), .A2(new_n956_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n957_), .A2(new_n653_), .ZN(new_n958_));
  XNOR2_X1  g757(.A(new_n958_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g758(.A1(new_n957_), .A2(new_n626_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(KEYINPUT125), .B(G204gat), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n960_), .B(new_n961_), .ZN(G1353gat));
  NOR3_X1   g761(.A1(new_n942_), .A2(new_n602_), .A3(new_n956_), .ZN(new_n963_));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n964_));
  INV_X1    g763(.A(KEYINPUT63), .ZN(new_n965_));
  INV_X1    g764(.A(G211gat), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n965_), .A2(new_n966_), .ZN(new_n967_));
  OR3_X1    g766(.A1(new_n963_), .A2(new_n964_), .A3(new_n967_), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n964_), .B1(new_n963_), .B2(new_n967_), .ZN(new_n969_));
  XOR2_X1   g768(.A(KEYINPUT63), .B(G211gat), .Z(new_n970_));
  AOI22_X1  g769(.A1(new_n968_), .A2(new_n969_), .B1(new_n963_), .B2(new_n970_), .ZN(G1354gat));
  AND3_X1   g770(.A1(new_n957_), .A2(G218gat), .A3(new_n707_), .ZN(new_n972_));
  NOR3_X1   g771(.A1(new_n942_), .A2(new_n720_), .A3(new_n956_), .ZN(new_n973_));
  OR2_X1    g772(.A1(new_n973_), .A2(KEYINPUT127), .ZN(new_n974_));
  AOI21_X1  g773(.A(G218gat), .B1(new_n973_), .B2(KEYINPUT127), .ZN(new_n975_));
  AOI21_X1  g774(.A(new_n972_), .B1(new_n974_), .B2(new_n975_), .ZN(G1355gat));
endmodule


