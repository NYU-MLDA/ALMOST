//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 1 1 0 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0 0 0 0 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n874_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT21), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT85), .ZN(new_n205_));
  INV_X1    g004(.A(G204gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n205_), .B1(new_n206_), .B2(G197gat), .ZN(new_n207_));
  INV_X1    g006(.A(G197gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n208_), .A2(KEYINPUT85), .A3(G204gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n206_), .A2(G197gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n207_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n204_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G218gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(G211gat), .ZN(new_n214_));
  INV_X1    g013(.A(G211gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(G218gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n208_), .A2(G204gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(new_n210_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n217_), .B1(KEYINPUT21), .B2(new_n219_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n207_), .A2(new_n209_), .A3(new_n203_), .A4(new_n210_), .ZN(new_n221_));
  AOI21_X1  g020(.A(KEYINPUT86), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n206_), .A2(G197gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n208_), .A2(G204gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT21), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  AND4_X1   g024(.A1(KEYINPUT86), .A2(new_n221_), .A3(new_n225_), .A4(new_n202_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n212_), .B1(new_n222_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(G190gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT26), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT26), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(G190gat), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G183gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT25), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT25), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(G183gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n232_), .A2(new_n234_), .A3(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT23), .B1(new_n233_), .B2(new_n228_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT23), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n239_), .A2(G183gat), .A3(G190gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(G169gat), .ZN(new_n242_));
  INV_X1    g041(.A(G176gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n244_), .A2(KEYINPUT24), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G169gat), .A2(G176gat), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n244_), .A2(KEYINPUT24), .A3(new_n247_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n237_), .A2(new_n241_), .A3(new_n246_), .A4(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n247_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT22), .B(G169gat), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n250_), .B1(new_n251_), .B2(new_n243_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n239_), .B1(G183gat), .B2(G190gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT79), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n240_), .A2(new_n254_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n239_), .A2(KEYINPUT79), .A3(G183gat), .A4(G190gat), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n253_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(G183gat), .A2(G190gat), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n252_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n249_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n227_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT77), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n262_), .B1(new_n235_), .B2(G183gat), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n233_), .A2(KEYINPUT77), .A3(KEYINPUT25), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n229_), .A2(new_n231_), .A3(new_n236_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n248_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT78), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  OAI211_X1 g068(.A(KEYINPUT78), .B(new_n248_), .C1(new_n265_), .C2(new_n266_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n257_), .A2(new_n245_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT86), .ZN(new_n273_));
  INV_X1    g072(.A(new_n221_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G197gat), .B(G204gat), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n202_), .B1(new_n275_), .B2(new_n203_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n273_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n220_), .A2(KEYINPUT86), .A3(new_n221_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n252_), .A2(KEYINPUT80), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n242_), .A2(KEYINPUT22), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT22), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(G169gat), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n281_), .A2(new_n283_), .A3(new_n243_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(new_n247_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT80), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n241_), .B1(G183gat), .B2(G190gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n280_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n272_), .A2(new_n279_), .A3(new_n212_), .A4(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n261_), .A2(new_n290_), .A3(KEYINPUT20), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G226gat), .A2(G233gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT19), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT88), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT20), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n272_), .A2(new_n289_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n295_), .B1(new_n296_), .B2(new_n227_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n260_), .ZN(new_n298_));
  AOI22_X1  g097(.A1(new_n277_), .A2(new_n278_), .B1(new_n211_), .B2(new_n204_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n293_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  AOI22_X1  g099(.A1(new_n291_), .A2(new_n294_), .B1(new_n297_), .B2(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(G8gat), .B(G36gat), .Z(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G64gat), .B(G92gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n301_), .A2(new_n306_), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n307_), .A2(KEYINPUT27), .ZN(new_n308_));
  INV_X1    g107(.A(new_n294_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n261_), .A2(new_n290_), .A3(KEYINPUT20), .A4(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n260_), .A2(KEYINPUT95), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT95), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n249_), .A2(new_n259_), .A3(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n311_), .A2(new_n299_), .A3(new_n313_), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n297_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n293_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n310_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n306_), .ZN(new_n318_));
  AOI21_X1  g117(.A(KEYINPUT98), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n316_), .B1(new_n297_), .B2(new_n314_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n310_), .ZN(new_n321_));
  OAI211_X1 g120(.A(KEYINPUT98), .B(new_n318_), .C1(new_n320_), .C2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n308_), .B1(new_n319_), .B2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n291_), .A2(new_n294_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n297_), .A2(new_n300_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n318_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT90), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n328_), .A2(new_n329_), .A3(new_n307_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n329_), .B1(new_n301_), .B2(new_n306_), .ZN(new_n331_));
  AND3_X1   g130(.A1(new_n325_), .A2(new_n326_), .A3(new_n306_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  XOR2_X1   g132(.A(KEYINPUT99), .B(KEYINPUT27), .Z(new_n334_));
  NAND3_X1  g133(.A1(new_n330_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n324_), .A2(new_n335_), .ZN(new_n336_));
  XOR2_X1   g135(.A(G127gat), .B(G134gat), .Z(new_n337_));
  XOR2_X1   g136(.A(G113gat), .B(G120gat), .Z(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(G155gat), .A2(G162gat), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT81), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G155gat), .A2(G162gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT82), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(KEYINPUT82), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G141gat), .A2(G148gat), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT2), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(G141gat), .ZN(new_n354_));
  INV_X1    g153(.A(G148gat), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(new_n355_), .A3(KEYINPUT3), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT3), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n357_), .B1(G141gat), .B2(G148gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n350_), .A2(new_n353_), .A3(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT83), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n356_), .A2(new_n358_), .B1(new_n352_), .B2(new_n351_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(KEYINPUT83), .A3(new_n350_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n345_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(G141gat), .A2(G148gat), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(new_n351_), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n344_), .B(KEYINPUT1), .Z(new_n369_));
  AOI21_X1  g168(.A(new_n368_), .B1(new_n369_), .B2(new_n343_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n340_), .B1(new_n365_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n345_), .ZN(new_n372_));
  AND3_X1   g171(.A1(new_n363_), .A2(KEYINPUT83), .A3(new_n350_), .ZN(new_n373_));
  AOI21_X1  g172(.A(KEYINPUT83), .B1(new_n363_), .B2(new_n350_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n372_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n370_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(new_n339_), .A3(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G225gat), .A2(G233gat), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n371_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT91), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT91), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n371_), .A2(new_n377_), .A3(new_n381_), .A4(new_n378_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n339_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT4), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n378_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n371_), .A2(KEYINPUT4), .A3(new_n377_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n383_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G1gat), .B(G29gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(G85gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT0), .B(G57gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n389_), .A2(KEYINPUT97), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT97), .ZN(new_n395_));
  AOI22_X1  g194(.A1(new_n380_), .A2(new_n382_), .B1(new_n387_), .B2(new_n386_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n393_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n395_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n393_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n383_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n394_), .A2(new_n398_), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  XOR2_X1   g201(.A(G22gat), .B(G50gat), .Z(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT29), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n375_), .A2(new_n405_), .A3(new_n376_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT28), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT84), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT28), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n375_), .A2(new_n409_), .A3(new_n405_), .A4(new_n376_), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n407_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n408_), .B1(new_n407_), .B2(new_n410_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n404_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n407_), .A2(new_n410_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT84), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n407_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n415_), .A2(new_n403_), .A3(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n375_), .A2(new_n376_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n299_), .B1(new_n418_), .B2(KEYINPUT29), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G228gat), .A2(G233gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(G78gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(G106gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n419_), .B(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n413_), .A2(new_n417_), .A3(KEYINPUT87), .A4(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n413_), .A2(new_n417_), .A3(KEYINPUT87), .ZN(new_n425_));
  INV_X1    g224(.A(new_n423_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(KEYINPUT87), .B1(new_n413_), .B2(new_n417_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n424_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G71gat), .B(G99gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(G43gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n296_), .B(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(new_n340_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G227gat), .A2(G233gat), .ZN(new_n434_));
  XOR2_X1   g233(.A(new_n434_), .B(G15gat), .Z(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT30), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT31), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n433_), .A2(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n433_), .A2(new_n437_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n336_), .A2(new_n402_), .A3(new_n429_), .A4(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n306_), .A2(KEYINPUT32), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n327_), .A2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n443_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT96), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  OAI211_X1 g246(.A(KEYINPUT96), .B(new_n443_), .C1(new_n320_), .C2(new_n321_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n444_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n401_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT92), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT33), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n451_), .B1(new_n400_), .B2(new_n452_), .ZN(new_n453_));
  AOI211_X1 g252(.A(KEYINPUT92), .B(KEYINPUT33), .C1(new_n383_), .C2(new_n399_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n331_), .A2(new_n332_), .ZN(new_n455_));
  NOR3_X1   g254(.A1(new_n327_), .A2(new_n329_), .A3(new_n318_), .ZN(new_n456_));
  OAI22_X1  g255(.A1(new_n453_), .A2(new_n454_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n378_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n371_), .A2(new_n377_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(new_n393_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT93), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n459_), .A2(KEYINPUT93), .A3(new_n393_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n387_), .B(new_n378_), .C1(KEYINPUT4), .C2(new_n371_), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT94), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n459_), .A2(KEYINPUT93), .A3(new_n393_), .ZN(new_n467_));
  AOI21_X1  g266(.A(KEYINPUT93), .B1(new_n459_), .B2(new_n393_), .ZN(new_n468_));
  OAI211_X1 g267(.A(KEYINPUT94), .B(new_n465_), .C1(new_n467_), .C2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  OAI22_X1  g269(.A1(new_n466_), .A2(new_n470_), .B1(new_n452_), .B2(new_n400_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n450_), .B1(new_n457_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(new_n429_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n424_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n425_), .A2(new_n426_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n428_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n474_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n336_), .A2(new_n477_), .A3(new_n402_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n473_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n440_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n442_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G1gat), .B(G8gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT75), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G15gat), .B(G22gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G1gat), .A2(G8gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT14), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n483_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n483_), .A2(new_n487_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G29gat), .B(G36gat), .Z(new_n491_));
  XOR2_X1   g290(.A(G43gat), .B(G50gat), .Z(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n490_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT76), .ZN(new_n495_));
  OR2_X1    g294(.A1(new_n490_), .A2(new_n493_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G229gat), .A2(G233gat), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n490_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n493_), .B(KEYINPUT15), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n503_), .A2(new_n498_), .A3(new_n494_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n500_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G113gat), .B(G141gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G169gat), .B(G197gat), .ZN(new_n507_));
  XOR2_X1   g306(.A(new_n506_), .B(new_n507_), .Z(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n505_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n500_), .A2(new_n504_), .A3(new_n508_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n481_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(G85gat), .ZN(new_n515_));
  INV_X1    g314(.A(G92gat), .ZN(new_n516_));
  NOR3_X1   g315(.A1(new_n515_), .A2(new_n516_), .A3(KEYINPUT9), .ZN(new_n517_));
  XOR2_X1   g316(.A(G85gat), .B(G92gat), .Z(new_n518_));
  AOI21_X1  g317(.A(new_n517_), .B1(new_n518_), .B2(KEYINPUT9), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT10), .B(G99gat), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n520_), .A2(G106gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT64), .B(KEYINPUT6), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n522_), .A2(G99gat), .A3(G106gat), .ZN(new_n523_));
  XOR2_X1   g322(.A(KEYINPUT64), .B(KEYINPUT6), .Z(new_n524_));
  NAND2_X1  g323(.A1(G99gat), .A2(G106gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n519_), .A2(new_n521_), .A3(new_n523_), .A4(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(G99gat), .A2(G106gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT7), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n526_), .A2(new_n523_), .A3(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n530_), .A2(new_n518_), .A3(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n531_), .B1(new_n530_), .B2(new_n518_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n527_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT66), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT66), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n536_), .B(new_n527_), .C1(new_n532_), .C2(new_n533_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G57gat), .B(G64gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT11), .ZN(new_n539_));
  XOR2_X1   g338(.A(G71gat), .B(G78gat), .Z(new_n540_));
  OR2_X1    g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n538_), .A2(KEYINPUT11), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n539_), .A2(new_n540_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n541_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT67), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n535_), .A2(new_n537_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n544_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n534_), .A2(KEYINPUT12), .A3(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n545_), .B1(new_n535_), .B2(new_n537_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n546_), .B(new_n548_), .C1(new_n549_), .C2(KEYINPUT12), .ZN(new_n550_));
  INV_X1    g349(.A(G230gat), .ZN(new_n551_));
  INV_X1    g350(.A(G233gat), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n550_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n546_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n553_), .B1(new_n555_), .B2(new_n549_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G120gat), .B(G148gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT5), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G176gat), .B(G204gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n559_), .B(new_n560_), .Z(new_n561_));
  NAND2_X1  g360(.A1(new_n557_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n561_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n554_), .A2(new_n556_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT13), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n562_), .A2(KEYINPUT13), .A3(new_n564_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n490_), .B(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n573_), .A2(new_n547_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT17), .ZN(new_n575_));
  XOR2_X1   g374(.A(G127gat), .B(G155gat), .Z(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT16), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G183gat), .B(G211gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  NOR3_X1   g378(.A1(new_n574_), .A2(new_n575_), .A3(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n580_), .B1(new_n544_), .B2(new_n572_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n573_), .A2(new_n545_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n573_), .A2(new_n545_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n579_), .B(KEYINPUT17), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n582_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n581_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n535_), .A2(new_n493_), .A3(new_n537_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G232gat), .A2(G233gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT34), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(KEYINPUT68), .B(KEYINPUT35), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  AOI22_X1  g392(.A1(new_n534_), .A2(new_n502_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n587_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n593_), .B1(new_n587_), .B2(new_n594_), .ZN(new_n596_));
  XOR2_X1   g395(.A(KEYINPUT71), .B(KEYINPUT36), .Z(new_n597_));
  XOR2_X1   g396(.A(G190gat), .B(G218gat), .Z(new_n598_));
  XNOR2_X1  g397(.A(G134gat), .B(G162gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NOR4_X1   g402(.A1(new_n595_), .A2(new_n596_), .A3(new_n597_), .A4(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n602_), .B(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n606_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(KEYINPUT74), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT74), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n609_), .B(new_n606_), .C1(new_n595_), .C2(new_n596_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n604_), .B1(new_n608_), .B2(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n611_), .A2(KEYINPUT37), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT73), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n607_), .A2(new_n613_), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n607_), .A2(new_n613_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n604_), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n615_), .A2(new_n616_), .A3(KEYINPUT37), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n612_), .B1(new_n614_), .B2(new_n617_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n514_), .A2(new_n570_), .A3(new_n586_), .A4(new_n618_), .ZN(new_n619_));
  OR3_X1    g418(.A1(new_n619_), .A2(G1gat), .A3(new_n402_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT38), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT102), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n611_), .B(KEYINPUT100), .Z(new_n624_));
  INV_X1    g423(.A(KEYINPUT101), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n627_), .A2(new_n481_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n570_), .A2(new_n512_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n586_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G1gat), .B1(new_n632_), .B2(new_n402_), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n623_), .B(new_n633_), .C1(new_n621_), .C2(new_n620_), .ZN(G1324gat));
  OR3_X1    g433(.A1(new_n619_), .A2(G8gat), .A3(new_n336_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n336_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n628_), .A2(new_n636_), .A3(new_n631_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT39), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n637_), .A2(new_n638_), .A3(G8gat), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n637_), .B2(G8gat), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n635_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g441(.A1(new_n628_), .A2(new_n440_), .A3(new_n631_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n643_), .A2(G15gat), .ZN(new_n644_));
  XOR2_X1   g443(.A(KEYINPUT103), .B(KEYINPUT41), .Z(new_n645_));
  OR2_X1    g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  OR3_X1    g445(.A1(new_n619_), .A2(G15gat), .A3(new_n480_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n644_), .A2(new_n645_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n646_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT104), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT104), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n646_), .A2(new_n651_), .A3(new_n647_), .A4(new_n648_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(G1326gat));
  OR3_X1    g452(.A1(new_n619_), .A2(G22gat), .A3(new_n429_), .ZN(new_n654_));
  OAI21_X1  g453(.A(G22gat), .B1(new_n632_), .B2(new_n429_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n655_), .A2(new_n656_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n654_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT106), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  OAI211_X1 g460(.A(KEYINPUT106), .B(new_n654_), .C1(new_n657_), .C2(new_n658_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1327gat));
  INV_X1    g462(.A(G29gat), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT43), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n617_), .A2(new_n614_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n666_), .B1(new_n611_), .B2(KEYINPUT37), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n440_), .B1(new_n473_), .B2(new_n478_), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n665_), .B(new_n667_), .C1(new_n668_), .C2(new_n442_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT107), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n429_), .A2(new_n401_), .ZN(new_n671_));
  AOI22_X1  g470(.A1(new_n472_), .A2(new_n429_), .B1(new_n671_), .B2(new_n336_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n441_), .B1(new_n672_), .B2(new_n440_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT107), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n673_), .A2(new_n674_), .A3(new_n665_), .A4(new_n667_), .ZN(new_n675_));
  OAI21_X1  g474(.A(KEYINPUT43), .B1(new_n481_), .B2(new_n618_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n670_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n629_), .A2(new_n586_), .ZN(new_n678_));
  AOI21_X1  g477(.A(KEYINPUT44), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n677_), .A2(KEYINPUT44), .A3(new_n678_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT108), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT108), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n677_), .A2(new_n682_), .A3(KEYINPUT44), .A4(new_n678_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n679_), .B1(new_n681_), .B2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n664_), .B1(new_n684_), .B2(new_n401_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT109), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n624_), .A2(new_n586_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n514_), .A2(new_n570_), .A3(new_n688_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n689_), .A2(G29gat), .A3(new_n402_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n686_), .A2(new_n687_), .A3(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT109), .B1(new_n685_), .B2(new_n690_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1328gat));
  NAND2_X1  g493(.A1(new_n681_), .A2(new_n683_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n679_), .A2(new_n336_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(G36gat), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT46), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n689_), .A2(G36gat), .A3(new_n336_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT45), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n698_), .A2(KEYINPUT110), .A3(new_n699_), .A4(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n699_), .A2(KEYINPUT110), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n699_), .A2(KEYINPUT110), .ZN(new_n705_));
  INV_X1    g504(.A(G36gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n704_), .B(new_n705_), .C1(new_n707_), .C2(new_n701_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n703_), .A2(new_n708_), .ZN(G1329gat));
  INV_X1    g508(.A(G43gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n710_), .B1(new_n689_), .B2(new_n480_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n684_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n440_), .A2(G43gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n711_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT47), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT47), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n716_), .B(new_n711_), .C1(new_n712_), .C2(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(G1330gat));
  OR3_X1    g517(.A1(new_n689_), .A2(G50gat), .A3(new_n429_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT111), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n684_), .A2(new_n720_), .A3(new_n477_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(G50gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n720_), .B1(new_n684_), .B2(new_n477_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n719_), .B1(new_n722_), .B2(new_n723_), .ZN(G1331gat));
  NAND2_X1  g523(.A1(new_n513_), .A2(new_n586_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n570_), .A2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n626_), .A2(new_n673_), .A3(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT113), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n728_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(G57gat), .B1(new_n731_), .B2(new_n402_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n618_), .A2(new_n569_), .A3(new_n586_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT112), .Z(new_n734_));
  NOR2_X1   g533(.A1(new_n481_), .A2(new_n512_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n402_), .A2(G57gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n732_), .B1(new_n736_), .B2(new_n737_), .ZN(G1332gat));
  INV_X1    g537(.A(KEYINPUT48), .ZN(new_n739_));
  INV_X1    g538(.A(new_n731_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(new_n636_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n739_), .B1(new_n741_), .B2(G64gat), .ZN(new_n742_));
  INV_X1    g541(.A(G64gat), .ZN(new_n743_));
  AOI211_X1 g542(.A(KEYINPUT48), .B(new_n743_), .C1(new_n740_), .C2(new_n636_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n636_), .A2(new_n743_), .ZN(new_n745_));
  OAI22_X1  g544(.A1(new_n742_), .A2(new_n744_), .B1(new_n736_), .B2(new_n745_), .ZN(G1333gat));
  OR3_X1    g545(.A1(new_n736_), .A2(G71gat), .A3(new_n480_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n729_), .A2(new_n440_), .A3(new_n730_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT49), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n748_), .A2(new_n749_), .A3(G71gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n748_), .B2(G71gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n747_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT114), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n747_), .B(KEYINPUT114), .C1(new_n750_), .C2(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1334gat));
  OR3_X1    g555(.A1(new_n736_), .A2(G78gat), .A3(new_n429_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n740_), .A2(new_n477_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT50), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n758_), .A2(new_n759_), .A3(G78gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n758_), .B2(G78gat), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n757_), .B1(new_n760_), .B2(new_n761_), .ZN(G1335gat));
  NOR3_X1   g561(.A1(new_n570_), .A2(new_n512_), .A3(new_n586_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n677_), .A2(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(G85gat), .B1(new_n764_), .B2(new_n402_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n688_), .A2(new_n569_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(new_n735_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n769_), .A2(new_n515_), .A3(new_n401_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n765_), .A2(new_n770_), .ZN(G1336gat));
  OAI21_X1  g570(.A(G92gat), .B1(new_n764_), .B2(new_n336_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n769_), .A2(new_n516_), .A3(new_n636_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(G1337gat));
  OR3_X1    g573(.A1(new_n768_), .A2(new_n480_), .A3(new_n520_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n677_), .A2(new_n440_), .A3(new_n763_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n776_), .A2(KEYINPUT115), .A3(G99gat), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT115), .B1(new_n776_), .B2(G99gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n775_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT51), .ZN(G1338gat));
  OR3_X1    g579(.A1(new_n768_), .A2(G106gat), .A3(new_n429_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n677_), .A2(new_n783_), .A3(new_n477_), .A4(new_n763_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n784_), .A2(G106gat), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n677_), .A2(new_n477_), .A3(new_n763_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT116), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n782_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n788_));
  AND4_X1   g587(.A1(new_n782_), .A2(new_n787_), .A3(G106gat), .A4(new_n784_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n781_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT53), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n792_), .B(new_n781_), .C1(new_n788_), .C2(new_n789_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(G1339gat));
  NAND2_X1  g593(.A1(new_n336_), .A2(new_n429_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n440_), .A2(new_n401_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n512_), .A2(new_n564_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n800_), .B1(new_n550_), .B2(new_n553_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n551_), .A2(new_n552_), .A3(KEYINPUT118), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n801_), .B(new_n803_), .C1(new_n800_), .C2(new_n550_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n550_), .A2(new_n800_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n563_), .B1(new_n805_), .B2(new_n802_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n804_), .A2(new_n806_), .A3(KEYINPUT56), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT56), .B1(new_n804_), .B2(new_n806_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n799_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n497_), .A2(new_n498_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n498_), .B1(new_n490_), .B2(new_n493_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n508_), .B1(new_n503_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n511_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n565_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n809_), .A2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n816_), .A2(new_n624_), .A3(KEYINPUT57), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n814_), .A2(new_n564_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n818_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  OAI221_X1 g620(.A(new_n818_), .B1(KEYINPUT120), .B2(KEYINPUT58), .C1(new_n807_), .C2(new_n808_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n821_), .A2(new_n822_), .A3(new_n667_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT57), .B1(new_n816_), .B2(new_n624_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n817_), .B(new_n823_), .C1(new_n824_), .C2(KEYINPUT119), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT119), .ZN(new_n826_));
  AOI211_X1 g625(.A(new_n826_), .B(KEYINPUT57), .C1(new_n816_), .C2(new_n624_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n630_), .B1(new_n825_), .B2(new_n827_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n725_), .B(KEYINPUT117), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n829_), .A2(new_n570_), .A3(new_n618_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(KEYINPUT54), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n798_), .B1(new_n828_), .B2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(G113gat), .B1(new_n832_), .B2(new_n512_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n798_), .A2(KEYINPUT59), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n817_), .A2(new_n823_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n824_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n586_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n830_), .B(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n834_), .B1(new_n837_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n832_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n841_), .B1(new_n842_), .B2(KEYINPUT59), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n512_), .A2(G113gat), .ZN(new_n844_));
  XOR2_X1   g643(.A(new_n844_), .B(KEYINPUT121), .Z(new_n845_));
  AOI21_X1  g644(.A(new_n833_), .B1(new_n843_), .B2(new_n845_), .ZN(G1340gat));
  NAND2_X1  g645(.A1(new_n843_), .A2(new_n569_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(G120gat), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT60), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n569_), .A2(new_n849_), .ZN(new_n850_));
  MUX2_X1   g649(.A(new_n850_), .B(new_n849_), .S(G120gat), .Z(new_n851_));
  OAI21_X1  g650(.A(new_n848_), .B1(new_n842_), .B2(new_n851_), .ZN(G1341gat));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n586_), .B(new_n840_), .C1(new_n832_), .C2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(G127gat), .ZN(new_n855_));
  INV_X1    g654(.A(G127gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n832_), .A2(new_n856_), .A3(new_n586_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n855_), .A2(KEYINPUT122), .A3(new_n857_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1342gat));
  NAND2_X1  g661(.A1(new_n843_), .A2(new_n667_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(G134gat), .ZN(new_n864_));
  OR2_X1    g663(.A1(new_n626_), .A2(G134gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n842_), .B2(new_n865_), .ZN(G1343gat));
  NAND2_X1  g665(.A1(new_n828_), .A2(new_n831_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NOR4_X1   g667(.A1(new_n636_), .A2(new_n429_), .A3(new_n402_), .A4(new_n440_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n868_), .A2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n512_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n569_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g674(.A1(new_n871_), .A2(new_n586_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(KEYINPUT61), .B(G155gat), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n876_), .B(new_n877_), .ZN(G1346gat));
  INV_X1    g677(.A(G162gat), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n867_), .A2(new_n879_), .A3(new_n627_), .A4(new_n869_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n868_), .A2(new_n618_), .A3(new_n870_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(new_n879_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(KEYINPUT123), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT123), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n880_), .B(new_n884_), .C1(new_n881_), .C2(new_n879_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(G1347gat));
  NOR2_X1   g685(.A1(new_n837_), .A2(new_n839_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n336_), .A2(new_n480_), .A3(new_n401_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n512_), .ZN(new_n889_));
  XOR2_X1   g688(.A(new_n889_), .B(KEYINPUT124), .Z(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n429_), .ZN(new_n891_));
  OAI21_X1  g690(.A(G169gat), .B1(new_n887_), .B2(new_n891_), .ZN(new_n892_));
  OR2_X1    g691(.A1(new_n892_), .A2(KEYINPUT125), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(KEYINPUT125), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n893_), .A2(KEYINPUT62), .A3(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n888_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n887_), .A2(new_n477_), .A3(new_n896_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n897_), .A2(new_n512_), .A3(new_n251_), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n895_), .B(new_n898_), .C1(KEYINPUT62), .C2(new_n894_), .ZN(G1348gat));
  AOI21_X1  g698(.A(G176gat), .B1(new_n897_), .B2(new_n569_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n569_), .A2(G176gat), .A3(new_n888_), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n868_), .A2(new_n477_), .A3(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT126), .ZN(new_n903_));
  OR3_X1    g702(.A1(new_n900_), .A2(new_n902_), .A3(new_n903_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n900_), .B2(new_n902_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1349gat));
  AOI21_X1  g705(.A(new_n630_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n867_), .A2(new_n429_), .A3(new_n586_), .A4(new_n888_), .ZN(new_n908_));
  AOI22_X1  g707(.A1(new_n897_), .A2(new_n907_), .B1(new_n908_), .B2(new_n233_), .ZN(G1350gat));
  NAND3_X1  g708(.A1(new_n897_), .A2(new_n232_), .A3(new_n627_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n228_), .B1(new_n897_), .B2(new_n667_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n911_), .A2(KEYINPUT127), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n911_), .A2(KEYINPUT127), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n910_), .B1(new_n912_), .B2(new_n913_), .ZN(G1351gat));
  AND4_X1   g713(.A1(new_n671_), .A2(new_n867_), .A3(new_n636_), .A4(new_n480_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n512_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g716(.A1(new_n915_), .A2(new_n569_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g718(.A(KEYINPUT63), .B(G211gat), .C1(new_n915_), .C2(new_n586_), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n915_), .A2(new_n586_), .ZN(new_n921_));
  XOR2_X1   g720(.A(KEYINPUT63), .B(G211gat), .Z(new_n922_));
  AOI21_X1  g721(.A(new_n920_), .B1(new_n921_), .B2(new_n922_), .ZN(G1354gat));
  NAND3_X1  g722(.A1(new_n915_), .A2(new_n213_), .A3(new_n627_), .ZN(new_n924_));
  AND2_X1   g723(.A1(new_n915_), .A2(new_n667_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n925_), .B2(new_n213_), .ZN(G1355gat));
endmodule


