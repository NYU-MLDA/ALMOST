//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0 1 0 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n685_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n763_, new_n764_,
    new_n765_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n780_, new_n781_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n939_, new_n940_, new_n941_,
    new_n943_, new_n944_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n952_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n959_, new_n960_, new_n961_;
  INV_X1    g000(.A(G190gat), .ZN(new_n202_));
  AND3_X1   g001(.A1(new_n202_), .A2(KEYINPUT80), .A3(KEYINPUT26), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT26), .B(G190gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT80), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n203_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(KEYINPUT79), .A2(G183gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT25), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT24), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G169gat), .B(G176gat), .ZN(new_n210_));
  OAI22_X1  g009(.A1(new_n206_), .A2(new_n208_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT81), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT23), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G183gat), .A3(G190gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  OAI221_X1 g017(.A(KEYINPUT81), .B1(new_n209_), .B2(new_n210_), .C1(new_n206_), .C2(new_n208_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n209_), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n213_), .A2(new_n218_), .A3(new_n219_), .A4(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT84), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n215_), .A2(new_n217_), .A3(new_n223_), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n216_), .A2(KEYINPUT84), .A3(G183gat), .A4(G190gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n224_), .A2(new_n225_), .A3(new_n227_), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n228_), .A2(KEYINPUT85), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(KEYINPUT85), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT82), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT22), .ZN(new_n232_));
  OAI21_X1  g031(.A(G169gat), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(G176gat), .ZN(new_n234_));
  INV_X1    g033(.A(G169gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(KEYINPUT82), .A3(KEYINPUT22), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n233_), .A2(new_n234_), .A3(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT83), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n235_), .A2(new_n234_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n240_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n229_), .A2(new_n230_), .A3(new_n239_), .A4(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n222_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G15gat), .B(G43gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT86), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT30), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n243_), .B(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G227gat), .A2(G233gat), .ZN(new_n248_));
  INV_X1    g047(.A(G71gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n247_), .B(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G127gat), .B(G134gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G113gat), .B(G120gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT87), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT31), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(G99gat), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n251_), .A2(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n251_), .A2(new_n258_), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G22gat), .B(G50gat), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(G155gat), .A2(G162gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT88), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G155gat), .A2(G162gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(G141gat), .ZN(new_n270_));
  INV_X1    g069(.A(G148gat), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT89), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT2), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT2), .ZN(new_n274_));
  OAI211_X1 g073(.A(KEYINPUT89), .B(new_n274_), .C1(new_n270_), .C2(new_n271_), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(G141gat), .A2(G148gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT3), .ZN(new_n278_));
  AOI21_X1  g077(.A(KEYINPUT90), .B1(new_n276_), .B2(new_n278_), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n278_), .A2(KEYINPUT90), .A3(new_n273_), .A4(new_n275_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n269_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT29), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n267_), .B(KEYINPUT1), .Z(new_n284_));
  NAND2_X1  g083(.A1(new_n266_), .A2(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(G141gat), .B(G148gat), .Z(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n282_), .A2(new_n283_), .A3(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT28), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n288_), .A2(KEYINPUT28), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n263_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n291_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(new_n289_), .A3(new_n262_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G78gat), .B(G106gat), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G228gat), .A2(G233gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n283_), .B1(new_n282_), .B2(new_n287_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G211gat), .B(G218gat), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT91), .ZN(new_n303_));
  INV_X1    g102(.A(G197gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(G204gat), .ZN(new_n305_));
  INV_X1    g104(.A(G204gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(G197gat), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT21), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n303_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n305_), .A2(new_n307_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n311_), .A2(KEYINPUT91), .A3(KEYINPUT21), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n302_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT92), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n314_), .B1(new_n306_), .B2(G197gat), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n304_), .A2(KEYINPUT92), .A3(G204gat), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n315_), .A2(new_n316_), .A3(new_n309_), .A4(new_n307_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT93), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n315_), .A2(new_n316_), .A3(new_n307_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n301_), .A2(new_n309_), .ZN(new_n320_));
  AOI22_X1  g119(.A1(new_n313_), .A2(new_n318_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n299_), .B1(new_n300_), .B2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n278_), .A2(new_n273_), .A3(new_n275_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT90), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n268_), .B1(new_n325_), .B2(new_n280_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n287_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT29), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n313_), .A2(new_n318_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n320_), .A2(new_n319_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n328_), .A2(new_n298_), .A3(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n297_), .B1(new_n322_), .B2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n295_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n322_), .A2(new_n332_), .A3(new_n297_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT95), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n335_), .B1(new_n333_), .B2(KEYINPUT94), .ZN(new_n338_));
  AND3_X1   g137(.A1(new_n328_), .A2(new_n298_), .A3(new_n331_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n298_), .B1(new_n328_), .B2(new_n331_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n296_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT94), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n295_), .B(new_n337_), .C1(new_n338_), .C2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n341_), .A2(new_n342_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n333_), .A2(KEYINPUT94), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n346_), .A2(new_n347_), .A3(new_n335_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n337_), .B1(new_n348_), .B2(new_n295_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n336_), .B1(new_n345_), .B2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n222_), .A2(new_n242_), .A3(new_n321_), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n351_), .A2(KEYINPUT20), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT103), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G226gat), .A2(G233gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT19), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(new_n220_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n358_), .A2(new_n225_), .A3(new_n224_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT97), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT25), .B(G183gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n204_), .A2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n362_), .B1(new_n357_), .B2(new_n210_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT97), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n358_), .A2(new_n224_), .A3(new_n365_), .A4(new_n225_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n360_), .A2(new_n364_), .A3(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT22), .B(G169gat), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n240_), .B1(new_n368_), .B2(new_n234_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n218_), .A2(new_n227_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n367_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n331_), .A2(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n352_), .A2(new_n353_), .A3(new_n356_), .A4(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT20), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n367_), .A2(new_n371_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n375_), .B1(new_n376_), .B2(new_n321_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n243_), .A2(new_n331_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(new_n355_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n351_), .A2(new_n373_), .A3(KEYINPUT20), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT103), .B1(new_n381_), .B2(new_n355_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n374_), .A2(new_n380_), .A3(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G8gat), .B(G36gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT18), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G64gat), .B(G92gat), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n385_), .B(new_n386_), .Z(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n383_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n381_), .A2(new_n355_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n377_), .A2(new_n378_), .A3(new_n356_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(new_n391_), .A3(new_n387_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n389_), .A2(KEYINPUT27), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT27), .ZN(new_n394_));
  INV_X1    g193(.A(new_n392_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n387_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n394_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n393_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G225gat), .A2(G233gat), .ZN(new_n400_));
  XOR2_X1   g199(.A(new_n400_), .B(KEYINPUT99), .Z(new_n401_));
  INV_X1    g200(.A(KEYINPUT4), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n256_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n282_), .A2(new_n287_), .A3(new_n254_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n402_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n282_), .A2(new_n287_), .ZN(new_n406_));
  AOI21_X1  g205(.A(KEYINPUT4), .B1(new_n406_), .B2(new_n256_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n401_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n254_), .B(KEYINPUT87), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n409_), .B1(new_n282_), .B2(new_n287_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n254_), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n326_), .A2(new_n327_), .A3(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n400_), .ZN(new_n413_));
  NOR3_X1   g212(.A1(new_n410_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G57gat), .B(G85gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT101), .ZN(new_n417_));
  INV_X1    g216(.A(G1gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT100), .B(KEYINPUT0), .ZN(new_n420_));
  INV_X1    g219(.A(G29gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n419_), .B(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n408_), .A2(new_n415_), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n424_), .B1(new_n408_), .B2(new_n415_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT105), .ZN(new_n428_));
  NOR3_X1   g227(.A1(new_n426_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n408_), .A2(new_n415_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n423_), .ZN(new_n431_));
  AOI21_X1  g230(.A(KEYINPUT105), .B1(new_n431_), .B2(new_n425_), .ZN(new_n432_));
  OR2_X1    g231(.A1(new_n429_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n350_), .A2(new_n399_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n390_), .A2(new_n391_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n387_), .A2(KEYINPUT32), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n438_), .B1(new_n431_), .B2(new_n425_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT104), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n383_), .A2(new_n440_), .A3(new_n437_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n440_), .B1(new_n383_), .B2(new_n437_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n439_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n425_), .A2(KEYINPUT33), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT33), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n408_), .A2(new_n415_), .A3(new_n445_), .A4(new_n424_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT98), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n448_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT102), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT4), .B1(new_n410_), .B2(new_n412_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n407_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n413_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n403_), .A2(new_n404_), .A3(new_n401_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n423_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n450_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n400_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n457_), .A2(KEYINPUT102), .A3(new_n423_), .A4(new_n454_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n435_), .A2(new_n388_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(KEYINPUT98), .A3(new_n392_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n447_), .A2(new_n449_), .A3(new_n459_), .A4(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n443_), .A2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n295_), .B1(new_n338_), .B2(new_n343_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT95), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n465_), .A2(new_n344_), .B1(new_n335_), .B2(new_n334_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n463_), .A2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n261_), .B1(new_n434_), .B2(new_n467_), .ZN(new_n468_));
  AND4_X1   g267(.A1(new_n466_), .A2(new_n399_), .A3(new_n433_), .A4(new_n261_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G190gat), .B(G218gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G134gat), .B(G162gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT36), .ZN(new_n474_));
  AND2_X1   g273(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n475_));
  NOR2_X1   g274(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(G106gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G99gat), .A2(G106gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT6), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT6), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(G99gat), .A3(G106gat), .ZN(new_n482_));
  AOI22_X1  g281(.A1(new_n477_), .A2(new_n478_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT9), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT64), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT64), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT9), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G85gat), .B(G92gat), .ZN(new_n489_));
  INV_X1    g288(.A(G92gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n484_), .A2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n488_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n492_));
  AND2_X1   g291(.A1(G85gat), .A2(G92gat), .ZN(new_n493_));
  NOR2_X1   g292(.A1(G85gat), .A2(G92gat), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n491_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n483_), .B1(new_n492_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT65), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n495_), .A2(new_n496_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n488_), .A2(new_n489_), .A3(new_n491_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT65), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(new_n503_), .A3(new_n483_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT7), .ZN(new_n505_));
  INV_X1    g304(.A(G99gat), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(new_n506_), .A3(new_n478_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT66), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n480_), .A2(new_n482_), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT66), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n511_), .A2(new_n505_), .A3(new_n506_), .A4(new_n478_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .A4(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n493_), .A2(new_n494_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT67), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT8), .B1(new_n514_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n515_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n513_), .A2(new_n514_), .A3(new_n517_), .ZN(new_n520_));
  AOI22_X1  g319(.A1(new_n499_), .A2(new_n504_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G29gat), .B(G36gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G43gat), .B(G50gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT35), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G232gat), .A2(G233gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT34), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n521_), .A2(new_n524_), .B1(new_n525_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT73), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT15), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n524_), .B(new_n531_), .ZN(new_n532_));
  NOR3_X1   g331(.A1(new_n521_), .A2(new_n530_), .A3(new_n532_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n502_), .A2(new_n503_), .A3(new_n483_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n503_), .B1(new_n502_), .B2(new_n483_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n520_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n517_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n537_));
  OAI22_X1  g336(.A1(new_n534_), .A2(new_n535_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n524_), .B(KEYINPUT15), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT73), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n529_), .B1(new_n533_), .B2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n528_), .A2(new_n525_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n473_), .A2(KEYINPUT36), .ZN(new_n544_));
  INV_X1    g343(.A(new_n542_), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n545_), .B(new_n529_), .C1(new_n533_), .C2(new_n540_), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n543_), .A2(new_n544_), .A3(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n544_), .B1(new_n543_), .B2(new_n546_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n474_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n470_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G1gat), .B(G8gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT76), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G15gat), .B(G22gat), .ZN(new_n553_));
  INV_X1    g352(.A(G8gat), .ZN(new_n554_));
  OAI21_X1  g353(.A(KEYINPUT14), .B1(new_n418_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n552_), .B(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G231gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT68), .B(G71gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(G78gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G57gat), .B(G64gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT11), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n562_), .A2(KEYINPUT11), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n561_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(G78gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n560_), .B(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(new_n563_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n566_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n559_), .B(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT17), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G127gat), .B(G155gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT16), .ZN(new_n574_));
  XOR2_X1   g373(.A(G183gat), .B(G211gat), .Z(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  NOR3_X1   g375(.A1(new_n571_), .A2(new_n572_), .A3(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(KEYINPUT17), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n577_), .B1(new_n571_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT13), .ZN(new_n580_));
  XOR2_X1   g379(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n581_));
  INV_X1    g380(.A(new_n570_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n581_), .B1(new_n521_), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G230gat), .A2(G233gat), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n538_), .A2(new_n570_), .A3(KEYINPUT12), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n521_), .A2(new_n582_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n583_), .A2(new_n584_), .A3(new_n585_), .A4(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n584_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n521_), .A2(new_n582_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n538_), .A2(new_n570_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n588_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(G120gat), .B(G148gat), .Z(new_n592_));
  XNOR2_X1  g391(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G176gat), .B(G204gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n587_), .A2(new_n591_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT71), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT71), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n587_), .A2(new_n591_), .A3(new_n600_), .A4(new_n597_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT72), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n587_), .A2(new_n591_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(new_n596_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n602_), .A2(new_n603_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n603_), .B1(new_n602_), .B2(new_n605_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n580_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n608_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(KEYINPUT13), .A3(new_n606_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G229gat), .A2(G233gat), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n557_), .A2(new_n524_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n557_), .A2(new_n524_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n613_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G113gat), .B(G141gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G169gat), .B(G197gat), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n618_), .B(new_n619_), .Z(new_n620_));
  NOR2_X1   g419(.A1(new_n532_), .A2(new_n557_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT77), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(KEYINPUT77), .B1(new_n532_), .B2(new_n557_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n613_), .B(KEYINPUT78), .Z(new_n626_));
  NAND2_X1  g425(.A1(new_n615_), .A2(new_n626_), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n617_), .B(new_n620_), .C1(new_n625_), .C2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n620_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n627_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n629_), .B1(new_n630_), .B2(new_n616_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n612_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n550_), .A2(new_n579_), .A3(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(G1gat), .B1(new_n635_), .B2(new_n433_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n350_), .A2(new_n398_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n637_), .A2(new_n433_), .A3(new_n261_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n429_), .A2(new_n432_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n465_), .A2(new_n344_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n639_), .B1(new_n640_), .B2(new_n336_), .ZN(new_n641_));
  AOI22_X1  g440(.A1(new_n641_), .A2(new_n399_), .B1(new_n466_), .B2(new_n463_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n638_), .B1(new_n642_), .B2(new_n261_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT37), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n543_), .A2(new_n544_), .A3(new_n546_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT74), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n644_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT75), .ZN(new_n649_));
  INV_X1    g448(.A(new_n546_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n530_), .B1(new_n521_), .B2(new_n532_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n538_), .A2(KEYINPUT73), .A3(new_n539_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n545_), .B1(new_n653_), .B2(new_n529_), .ZN(new_n654_));
  OAI22_X1  g453(.A1(new_n650_), .A2(new_n654_), .B1(KEYINPUT36), .B2(new_n473_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(new_n645_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n649_), .B1(new_n656_), .B2(new_n474_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n474_), .ZN(new_n658_));
  AOI211_X1 g457(.A(KEYINPUT75), .B(new_n658_), .C1(new_n655_), .C2(new_n645_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n648_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n549_), .A2(KEYINPUT75), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n656_), .A2(new_n649_), .A3(new_n474_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n661_), .A2(new_n647_), .A3(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n660_), .A2(new_n663_), .A3(new_n579_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n643_), .A2(new_n665_), .A3(new_n634_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT38), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n639_), .A2(new_n418_), .ZN(new_n668_));
  OR3_X1    g467(.A1(new_n666_), .A2(new_n667_), .A3(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n667_), .B1(new_n666_), .B2(new_n668_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n636_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT106), .ZN(G1324gat));
  OAI21_X1  g471(.A(G8gat), .B1(new_n635_), .B2(new_n399_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT39), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n666_), .A2(G8gat), .A3(new_n399_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n676_), .B(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n673_), .A2(new_n674_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n675_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT40), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n675_), .A2(new_n678_), .A3(KEYINPUT40), .A4(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1325gat));
  INV_X1    g483(.A(new_n261_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G15gat), .B1(new_n635_), .B2(new_n685_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT41), .Z(new_n687_));
  OR2_X1    g486(.A1(new_n685_), .A2(G15gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n687_), .B1(new_n666_), .B2(new_n688_), .ZN(G1326gat));
  OAI21_X1  g488(.A(G22gat), .B1(new_n635_), .B2(new_n466_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT42), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n466_), .A2(G22gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(new_n666_), .B2(new_n692_), .ZN(G1327gat));
  INV_X1    g492(.A(new_n549_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n694_), .A2(new_n579_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n643_), .A2(new_n634_), .A3(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(KEYINPUT108), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT108), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n643_), .A2(new_n698_), .A3(new_n634_), .A4(new_n695_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(G29gat), .B1(new_n700_), .B2(new_n639_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n612_), .A2(new_n579_), .A3(new_n633_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n657_), .A2(new_n659_), .A3(new_n648_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n647_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n703_), .B1(new_n643_), .B2(new_n707_), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n703_), .B(new_n707_), .C1(new_n468_), .C2(new_n469_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n702_), .B1(new_n708_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(KEYINPUT43), .B1(new_n470_), .B2(new_n706_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n709_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n715_), .A2(KEYINPUT44), .A3(new_n702_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n713_), .A2(new_n716_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n433_), .A2(new_n421_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n701_), .B1(new_n717_), .B2(new_n718_), .ZN(G1328gat));
  NAND3_X1  g518(.A1(new_n713_), .A2(new_n398_), .A3(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(G36gat), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT109), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT110), .B1(new_n722_), .B2(KEYINPUT46), .ZN(new_n723_));
  NOR2_X1   g522(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n399_), .A2(G36gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n697_), .A2(new_n699_), .A3(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT45), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT45), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n697_), .A2(new_n728_), .A3(new_n699_), .A4(new_n725_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n724_), .B1(new_n727_), .B2(new_n729_), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n721_), .A2(new_n723_), .A3(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n723_), .B1(new_n721_), .B2(new_n730_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1329gat));
  NAND4_X1  g532(.A1(new_n713_), .A2(new_n716_), .A3(G43gat), .A4(new_n261_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n697_), .A2(new_n261_), .A3(new_n699_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT111), .ZN(new_n736_));
  INV_X1    g535(.A(G43gat), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n735_), .A2(new_n736_), .A3(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n736_), .B1(new_n735_), .B2(new_n737_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n734_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT47), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT47), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n734_), .B(new_n742_), .C1(new_n738_), .C2(new_n739_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1330gat));
  AOI21_X1  g543(.A(G50gat), .B1(new_n700_), .B2(new_n350_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n350_), .A2(G50gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n717_), .B2(new_n746_), .ZN(G1331gat));
  NAND4_X1  g546(.A1(new_n550_), .A2(new_n579_), .A3(new_n633_), .A4(new_n612_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G57gat), .B1(new_n748_), .B2(new_n433_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n470_), .A2(new_n632_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n750_), .A2(new_n665_), .A3(new_n612_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n433_), .A2(G57gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n749_), .B1(new_n751_), .B2(new_n752_), .ZN(G1332gat));
  OAI21_X1  g552(.A(G64gat), .B1(new_n748_), .B2(new_n399_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT48), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n399_), .A2(G64gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n755_), .B1(new_n751_), .B2(new_n756_), .ZN(G1333gat));
  OAI21_X1  g556(.A(G71gat), .B1(new_n748_), .B2(new_n685_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT49), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n261_), .A2(new_n249_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT112), .Z(new_n761_));
  OAI21_X1  g560(.A(new_n759_), .B1(new_n751_), .B2(new_n761_), .ZN(G1334gat));
  OAI21_X1  g561(.A(G78gat), .B1(new_n748_), .B2(new_n466_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT50), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n350_), .A2(new_n567_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n751_), .B2(new_n765_), .ZN(G1335gat));
  AND2_X1   g565(.A1(new_n612_), .A2(new_n695_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n750_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(G85gat), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n770_), .A3(new_n639_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n579_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n612_), .A2(new_n772_), .A3(new_n633_), .ZN(new_n773_));
  OR2_X1    g572(.A1(new_n773_), .A2(KEYINPUT113), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(KEYINPUT113), .ZN(new_n775_));
  AOI22_X1  g574(.A1(new_n714_), .A2(new_n709_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT114), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n777_), .A2(new_n639_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n771_), .B1(new_n778_), .B2(new_n770_), .ZN(G1336gat));
  NAND3_X1  g578(.A1(new_n769_), .A2(new_n490_), .A3(new_n398_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n777_), .A2(new_n398_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(new_n490_), .ZN(G1337gat));
  NAND2_X1  g581(.A1(new_n261_), .A2(new_n477_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT51), .ZN(new_n784_));
  OAI22_X1  g583(.A1(new_n768_), .A2(new_n783_), .B1(KEYINPUT115), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n776_), .A2(new_n261_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n786_), .B2(G99gat), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n784_), .A2(KEYINPUT115), .ZN(new_n788_));
  XOR2_X1   g587(.A(new_n787_), .B(new_n788_), .Z(G1338gat));
  NAND3_X1  g588(.A1(new_n769_), .A2(new_n478_), .A3(new_n350_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n776_), .A2(new_n350_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(G106gat), .ZN(new_n793_));
  AOI211_X1 g592(.A(KEYINPUT52), .B(new_n478_), .C1(new_n776_), .C2(new_n350_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n790_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT53), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n797_), .B(new_n790_), .C1(new_n793_), .C2(new_n794_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(G1339gat));
  NOR2_X1   g598(.A1(new_n685_), .A2(new_n433_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n637_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n602_), .A2(new_n632_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT116), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n602_), .A2(new_n804_), .A3(new_n632_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n588_), .A2(KEYINPUT118), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n583_), .A2(new_n586_), .A3(new_n585_), .A4(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n584_), .A2(new_n809_), .ZN(new_n810_));
  AND4_X1   g609(.A1(new_n586_), .A2(new_n583_), .A3(new_n585_), .A4(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n808_), .B1(new_n811_), .B2(new_n807_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n587_), .A2(new_n809_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n587_), .A2(KEYINPUT117), .A3(new_n809_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n812_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT56), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT119), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n817_), .A2(new_n596_), .A3(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n817_), .B2(new_n596_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n803_), .B(new_n805_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n614_), .A2(new_n615_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n620_), .B1(new_n823_), .B2(new_n626_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n626_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n615_), .A2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n824_), .B1(new_n625_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n628_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n822_), .A2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(KEYINPUT57), .A3(new_n694_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT120), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n694_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n549_), .B1(new_n822_), .B2(new_n830_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(new_n838_), .A3(KEYINPUT57), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT58), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n817_), .A2(new_n818_), .A3(new_n596_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n828_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n818_), .B1(new_n817_), .B2(new_n596_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n840_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n844_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n846_), .A2(KEYINPUT58), .A3(new_n841_), .A4(new_n842_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n845_), .B(new_n847_), .C1(new_n704_), .C2(new_n705_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n833_), .A2(new_n836_), .A3(new_n839_), .A4(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n772_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT54), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n609_), .A2(new_n611_), .A3(new_n633_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n851_), .B1(new_n665_), .B2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n609_), .A2(new_n611_), .A3(new_n633_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n854_), .A2(new_n664_), .A3(KEYINPUT54), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n853_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n801_), .B1(new_n850_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(G113gat), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n858_), .A2(new_n859_), .A3(new_n632_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n861_));
  INV_X1    g660(.A(new_n801_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n848_), .B1(KEYINPUT57), .B2(new_n837_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n838_), .B1(new_n837_), .B2(KEYINPUT57), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n579_), .B1(new_n865_), .B2(new_n839_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n861_), .B(new_n862_), .C1(new_n866_), .C2(new_n856_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n858_), .A2(new_n861_), .A3(KEYINPUT59), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n633_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n860_), .B1(new_n871_), .B2(new_n859_), .ZN(G1340gat));
  INV_X1    g671(.A(G120gat), .ZN(new_n873_));
  INV_X1    g672(.A(new_n612_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n874_), .B2(KEYINPUT60), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n858_), .B(new_n875_), .C1(KEYINPUT60), .C2(new_n873_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n874_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n877_), .B2(new_n873_), .ZN(G1341gat));
  INV_X1    g677(.A(G127gat), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n858_), .A2(new_n879_), .A3(new_n579_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n772_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(new_n879_), .ZN(G1342gat));
  INV_X1    g681(.A(G134gat), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n706_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n885_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n886_));
  AOI21_X1  g685(.A(G134gat), .B1(new_n858_), .B2(new_n549_), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT122), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(KEYINPUT59), .B1(new_n858_), .B2(new_n861_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n856_), .B1(new_n849_), .B2(new_n772_), .ZN(new_n890_));
  NOR4_X1   g689(.A1(new_n890_), .A2(KEYINPUT121), .A3(new_n868_), .A4(new_n801_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n884_), .B1(new_n889_), .B2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n893_));
  INV_X1    g692(.A(new_n887_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n892_), .A2(new_n893_), .A3(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n888_), .A2(new_n895_), .ZN(G1343gat));
  NAND2_X1  g695(.A1(new_n850_), .A2(new_n857_), .ZN(new_n897_));
  NOR4_X1   g696(.A1(new_n466_), .A2(new_n433_), .A3(new_n261_), .A4(new_n398_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(new_n633_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(new_n270_), .ZN(G1344gat));
  NOR2_X1   g700(.A1(new_n899_), .A2(new_n874_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(new_n271_), .ZN(G1345gat));
  AND2_X1   g702(.A1(new_n897_), .A2(new_n898_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n904_), .A2(new_n905_), .A3(new_n579_), .ZN(new_n906_));
  OAI21_X1  g705(.A(KEYINPUT123), .B1(new_n899_), .B2(new_n772_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT61), .B(G155gat), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n906_), .A2(new_n907_), .A3(new_n909_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1346gat));
  OR3_X1    g712(.A1(new_n899_), .A2(G162gat), .A3(new_n694_), .ZN(new_n914_));
  OAI21_X1  g713(.A(G162gat), .B1(new_n899_), .B2(new_n706_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1347gat));
  NOR3_X1   g715(.A1(new_n685_), .A2(new_n639_), .A3(new_n399_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n633_), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n466_), .B(new_n919_), .C1(new_n866_), .C2(new_n856_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n920_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n890_), .A2(new_n350_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n922_), .A2(new_n368_), .A3(new_n919_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(KEYINPUT62), .B1(new_n920_), .B2(G169gat), .ZN(new_n925_));
  OAI21_X1  g724(.A(KEYINPUT124), .B1(new_n924_), .B2(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n925_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n928_));
  NAND4_X1  g727(.A1(new_n927_), .A2(new_n928_), .A3(new_n923_), .A4(new_n921_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n926_), .A2(new_n929_), .ZN(G1348gat));
  NAND2_X1  g729(.A1(new_n922_), .A2(new_n917_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n931_), .ZN(new_n932_));
  AOI21_X1  g731(.A(G176gat), .B1(new_n932_), .B2(new_n612_), .ZN(new_n933_));
  OR2_X1    g732(.A1(new_n922_), .A2(KEYINPUT125), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n922_), .A2(KEYINPUT125), .ZN(new_n935_));
  AND2_X1   g734(.A1(new_n934_), .A2(new_n935_), .ZN(new_n936_));
  NOR3_X1   g735(.A1(new_n918_), .A2(new_n234_), .A3(new_n874_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n933_), .B1(new_n936_), .B2(new_n937_), .ZN(G1349gat));
  NOR3_X1   g737(.A1(new_n931_), .A2(new_n772_), .A3(new_n361_), .ZN(new_n939_));
  NAND4_X1  g738(.A1(new_n934_), .A2(new_n579_), .A3(new_n917_), .A4(new_n935_), .ZN(new_n940_));
  INV_X1    g739(.A(G183gat), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n939_), .B1(new_n940_), .B2(new_n941_), .ZN(G1350gat));
  OAI21_X1  g741(.A(G190gat), .B1(new_n931_), .B2(new_n706_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n549_), .A2(new_n204_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n943_), .B1(new_n931_), .B2(new_n944_), .ZN(G1351gat));
  NAND2_X1  g744(.A1(new_n641_), .A2(new_n685_), .ZN(new_n946_));
  AND2_X1   g745(.A1(new_n946_), .A2(KEYINPUT126), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n398_), .B1(new_n946_), .B2(KEYINPUT126), .ZN(new_n948_));
  NOR3_X1   g747(.A1(new_n890_), .A2(new_n947_), .A3(new_n948_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n949_), .A2(new_n632_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g750(.A1(new_n949_), .A2(new_n612_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n952_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g752(.A1(new_n949_), .A2(new_n579_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n955_));
  AND2_X1   g754(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n956_));
  NOR3_X1   g755(.A1(new_n954_), .A2(new_n955_), .A3(new_n956_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n957_), .B1(new_n954_), .B2(new_n955_), .ZN(G1354gat));
  NAND2_X1  g757(.A1(new_n949_), .A2(new_n549_), .ZN(new_n959_));
  XNOR2_X1  g758(.A(KEYINPUT127), .B(G218gat), .ZN(new_n960_));
  NOR2_X1   g759(.A1(new_n706_), .A2(new_n960_), .ZN(new_n961_));
  AOI22_X1  g760(.A1(new_n959_), .A2(new_n960_), .B1(new_n949_), .B2(new_n961_), .ZN(G1355gat));
endmodule


