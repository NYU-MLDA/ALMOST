//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 0 1 1 0 1 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 1 0 0 0 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n809_, new_n810_, new_n811_, new_n813_, new_n814_,
    new_n815_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n836_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n880_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_;
  AND3_X1   g000(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n202_));
  AOI21_X1  g001(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G99gat), .ZN(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n205_), .A2(new_n206_), .A3(KEYINPUT69), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT7), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT7), .ZN(new_n209_));
  NAND4_X1  g008(.A1(new_n209_), .A2(new_n205_), .A3(new_n206_), .A4(KEYINPUT69), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n204_), .A2(new_n208_), .A3(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(G85gat), .ZN(new_n212_));
  INV_X1    g011(.A(G92gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G85gat), .A2(G92gat), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n211_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT70), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT70), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n211_), .A2(new_n219_), .A3(new_n216_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(KEYINPUT8), .A3(new_n220_), .ZN(new_n221_));
  AOI211_X1 g020(.A(new_n219_), .B(KEYINPUT8), .C1(new_n211_), .C2(new_n216_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G57gat), .B(G64gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT11), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G71gat), .B(G78gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n224_), .A2(KEYINPUT11), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n226_), .B1(KEYINPUT11), .B2(new_n224_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n228_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n202_), .A2(new_n203_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT10), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(new_n205_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n206_), .A3(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n235_), .A2(KEYINPUT66), .A3(new_n206_), .A4(new_n236_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n233_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n215_), .A2(KEYINPUT67), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT9), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT9), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n215_), .A2(KEYINPUT67), .A3(new_n244_), .ZN(new_n245_));
  AND4_X1   g044(.A1(KEYINPUT68), .A2(new_n243_), .A3(new_n214_), .A4(new_n245_), .ZN(new_n246_));
  AOI22_X1  g045(.A1(new_n242_), .A2(KEYINPUT9), .B1(new_n212_), .B2(new_n213_), .ZN(new_n247_));
  AOI21_X1  g046(.A(KEYINPUT68), .B1(new_n247_), .B2(new_n245_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n241_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n221_), .A2(new_n223_), .A3(new_n232_), .A4(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G230gat), .A2(G233gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n250_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n220_), .A2(KEYINPUT8), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n219_), .B1(new_n211_), .B2(new_n216_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n249_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n231_), .B1(new_n258_), .B2(new_n222_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT12), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT12), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n261_), .B(new_n231_), .C1(new_n258_), .C2(new_n222_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n255_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n254_), .B1(new_n259_), .B2(new_n250_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G120gat), .B(G148gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT5), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G176gat), .B(G204gat), .ZN(new_n267_));
  XOR2_X1   g066(.A(new_n266_), .B(new_n267_), .Z(new_n268_));
  OR3_X1    g067(.A1(new_n263_), .A2(new_n264_), .A3(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n268_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT13), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT72), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  OR3_X1    g073(.A1(new_n272_), .A2(KEYINPUT72), .A3(new_n273_), .ZN(new_n275_));
  AOI21_X1  g074(.A(KEYINPUT71), .B1(new_n272_), .B2(new_n273_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n272_), .A2(new_n273_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n274_), .B(new_n275_), .C1(new_n276_), .C2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(G1gat), .ZN(new_n281_));
  INV_X1    g080(.A(G8gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT14), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(KEYINPUT79), .B(G15gat), .Z(new_n284_));
  OAI21_X1  g083(.A(new_n283_), .B1(new_n284_), .B2(G22gat), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n285_), .B1(G22gat), .B2(new_n284_), .ZN(new_n286_));
  XOR2_X1   g085(.A(G1gat), .B(G8gat), .Z(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n286_), .B(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G29gat), .B(G36gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G43gat), .B(G50gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(new_n292_), .ZN(new_n293_));
  XOR2_X1   g092(.A(new_n292_), .B(KEYINPUT15), .Z(new_n294_));
  OAI21_X1  g093(.A(new_n293_), .B1(new_n294_), .B2(new_n289_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G229gat), .A2(G233gat), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n289_), .B(new_n292_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n298_), .A2(new_n296_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G113gat), .B(G141gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G169gat), .B(G197gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  OR3_X1    g102(.A1(new_n297_), .A2(new_n299_), .A3(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n303_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n280_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT20), .ZN(new_n308_));
  INV_X1    g107(.A(G183gat), .ZN(new_n309_));
  INV_X1    g108(.A(G190gat), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT23), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT80), .B(KEYINPUT23), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(new_n311_), .ZN(new_n315_));
  AOI22_X1  g114(.A1(new_n313_), .A2(new_n315_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n316_));
  INV_X1    g115(.A(G176gat), .ZN(new_n317_));
  INV_X1    g116(.A(G169gat), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT81), .B1(new_n318_), .B2(KEYINPUT22), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT22), .B(G169gat), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n317_), .B(new_n319_), .C1(new_n320_), .C2(KEYINPUT81), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT25), .B(G183gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT26), .B(G190gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(G169gat), .A2(G176gat), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n328_), .A2(KEYINPUT24), .A3(new_n322_), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n326_), .B(new_n329_), .C1(KEYINPUT24), .C2(new_n328_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n312_), .A2(new_n314_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n331_), .B1(new_n332_), .B2(new_n312_), .ZN(new_n333_));
  OAI22_X1  g132(.A1(new_n316_), .A2(new_n323_), .B1(new_n330_), .B2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G211gat), .B(G218gat), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT91), .ZN(new_n336_));
  INV_X1    g135(.A(G204gat), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n336_), .B1(new_n337_), .B2(G197gat), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n335_), .A2(KEYINPUT21), .A3(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G197gat), .B(G204gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n340_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n342_), .A2(KEYINPUT21), .A3(new_n335_), .A4(new_n338_), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n335_), .A2(KEYINPUT21), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n341_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n308_), .B1(new_n334_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G226gat), .A2(G233gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT19), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n313_), .A2(new_n315_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT95), .B(KEYINPUT24), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n324_), .A2(new_n325_), .B1(new_n352_), .B2(new_n327_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n322_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT96), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(new_n328_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n355_), .A2(new_n356_), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n351_), .B(new_n353_), .C1(new_n358_), .C2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n309_), .A2(new_n310_), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n331_), .B(new_n361_), .C1(new_n332_), .C2(new_n312_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT97), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n320_), .B(new_n363_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n362_), .B(new_n322_), .C1(new_n364_), .C2(G176gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n360_), .A2(new_n365_), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n347_), .B(new_n350_), .C1(new_n366_), .C2(new_n346_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G8gat), .B(G36gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT18), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G64gat), .B(G92gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n360_), .A2(new_n346_), .A3(new_n365_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n334_), .A2(new_n345_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n308_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n367_), .B(new_n372_), .C1(new_n375_), .C2(new_n350_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n376_), .A2(KEYINPUT98), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n376_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n367_), .B1(new_n375_), .B2(new_n350_), .ZN(new_n380_));
  AOI21_X1  g179(.A(KEYINPUT98), .B1(new_n380_), .B2(new_n371_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n378_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT27), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n345_), .B(KEYINPUT94), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n347_), .B1(new_n384_), .B2(new_n366_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n349_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n375_), .A2(new_n350_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n371_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n379_), .A2(new_n383_), .ZN(new_n390_));
  AOI22_X1  g189(.A1(new_n382_), .A2(new_n383_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G127gat), .B(G134gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G113gat), .B(G120gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G141gat), .A2(G148gat), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(G141gat), .A2(G148gat), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(G155gat), .ZN(new_n400_));
  INV_X1    g199(.A(G162gat), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n400_), .A2(new_n401_), .A3(KEYINPUT84), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT84), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n403_), .B1(G155gat), .B2(G162gat), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT86), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G155gat), .A2(G162gat), .ZN(new_n407_));
  AOI21_X1  g206(.A(KEYINPUT85), .B1(new_n407_), .B2(KEYINPUT1), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(KEYINPUT85), .A3(KEYINPUT1), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n405_), .A2(new_n406_), .A3(new_n409_), .A4(new_n410_), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n407_), .A2(KEYINPUT1), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n402_), .A2(new_n404_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n414_), .A2(new_n408_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n406_), .B1(new_n415_), .B2(new_n410_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n399_), .B1(new_n413_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n405_), .A2(new_n407_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n398_), .A2(KEYINPUT87), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT3), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n396_), .B(KEYINPUT2), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n419_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n395_), .B1(new_n418_), .B2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n405_), .A2(new_n410_), .A3(new_n409_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT86), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n424_), .B1(new_n428_), .B2(new_n399_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n394_), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n425_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G225gat), .A2(G233gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n429_), .A2(new_n394_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT4), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n432_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n425_), .A2(new_n430_), .A3(KEYINPUT4), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n433_), .A2(new_n438_), .ZN(new_n439_));
  XOR2_X1   g238(.A(G1gat), .B(G29gat), .Z(new_n440_));
  XNOR2_X1  g239(.A(G57gat), .B(G85gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n443_));
  XOR2_X1   g242(.A(new_n442_), .B(new_n443_), .Z(new_n444_));
  NAND2_X1  g243(.A1(new_n439_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n444_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n433_), .A2(new_n438_), .A3(KEYINPUT100), .A4(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  AOI22_X1  g247(.A1(new_n431_), .A2(new_n432_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n449_));
  AOI21_X1  g248(.A(KEYINPUT100), .B1(new_n449_), .B2(new_n446_), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT101), .B1(new_n448_), .B2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n433_), .A2(new_n438_), .A3(new_n446_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT100), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT101), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n454_), .A2(new_n445_), .A3(new_n455_), .A4(new_n447_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n391_), .A2(new_n451_), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT29), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n429_), .A2(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(G22gat), .B(G50gat), .Z(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT94), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n345_), .B(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n424_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n459_), .B1(new_n417_), .B2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n465_), .B1(new_n467_), .B2(KEYINPUT93), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT93), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n469_), .B1(new_n429_), .B2(new_n459_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  AND2_X1   g270(.A1(KEYINPUT89), .A2(G228gat), .ZN(new_n472_));
  NOR2_X1   g271(.A1(KEYINPUT89), .A2(G228gat), .ZN(new_n473_));
  OAI21_X1  g272(.A(G233gat), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT90), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n471_), .A2(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n345_), .A2(new_n475_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT92), .B1(new_n467_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT92), .ZN(new_n480_));
  OAI211_X1 g279(.A(new_n480_), .B(new_n477_), .C1(new_n429_), .C2(new_n459_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G78gat), .B(G106gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n476_), .A2(new_n483_), .A3(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n475_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n487_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n484_), .B1(new_n488_), .B2(new_n482_), .ZN(new_n489_));
  XOR2_X1   g288(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n490_));
  AND3_X1   g289(.A1(new_n486_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n490_), .B1(new_n486_), .B2(new_n489_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n463_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(new_n334_), .B(KEYINPUT30), .Z(new_n494_));
  XNOR2_X1  g293(.A(G71gat), .B(G99gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT83), .ZN(new_n496_));
  XOR2_X1   g295(.A(G15gat), .B(G43gat), .Z(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G227gat), .A2(G233gat), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n499_), .B(KEYINPUT82), .Z(new_n500_));
  XNOR2_X1  g299(.A(new_n498_), .B(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n494_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n334_), .B(KEYINPUT30), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n498_), .A2(new_n500_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n498_), .A2(new_n500_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT31), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n502_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n507_), .B1(new_n502_), .B2(new_n506_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n395_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n510_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n512_), .A2(new_n394_), .A3(new_n508_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n490_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n485_), .B1(new_n476_), .B2(new_n483_), .ZN(new_n516_));
  NOR3_X1   g315(.A1(new_n488_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n515_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n486_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(new_n462_), .A3(new_n519_), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n493_), .A2(new_n514_), .A3(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n514_), .B1(new_n493_), .B2(new_n520_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n458_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n511_), .A2(new_n513_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n388_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n372_), .A2(KEYINPUT32), .ZN(new_n526_));
  MUX2_X1   g325(.A(new_n525_), .B(new_n380_), .S(new_n526_), .Z(new_n527_));
  OAI21_X1  g326(.A(new_n527_), .B1(new_n448_), .B2(new_n450_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n380_), .A2(new_n371_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT98), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n377_), .B1(new_n531_), .B2(new_n376_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n425_), .A2(new_n430_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n437_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n432_), .B1(new_n425_), .B2(KEYINPUT4), .ZN(new_n535_));
  OAI221_X1 g334(.A(new_n444_), .B1(new_n533_), .B2(new_n432_), .C1(new_n534_), .C2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT33), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n452_), .A2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n449_), .A2(KEYINPUT33), .A3(new_n446_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n532_), .A2(new_n536_), .A3(new_n538_), .A4(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n524_), .B1(new_n528_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n493_), .A2(new_n520_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n307_), .B1(new_n523_), .B2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G190gat), .B(G218gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT74), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G134gat), .B(G162gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT36), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT77), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n258_), .A2(new_n222_), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n552_), .A2(new_n294_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n292_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G232gat), .A2(G233gat), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n555_), .B(KEYINPUT34), .Z(new_n556_));
  XOR2_X1   g355(.A(KEYINPUT73), .B(KEYINPUT35), .Z(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n553_), .A2(new_n554_), .A3(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n556_), .A2(new_n557_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n560_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n553_), .A2(new_n562_), .A3(new_n554_), .A4(new_n558_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n551_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT37), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n565_), .A2(KEYINPUT78), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n548_), .A2(new_n549_), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n568_), .B(KEYINPUT75), .Z(new_n569_));
  NAND3_X1  g368(.A1(new_n561_), .A2(new_n563_), .A3(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(KEYINPUT76), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT76), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n561_), .A2(new_n572_), .A3(new_n563_), .A4(new_n569_), .ZN(new_n573_));
  AOI211_X1 g372(.A(new_n564_), .B(new_n567_), .C1(new_n571_), .C2(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n564_), .B1(new_n571_), .B2(new_n573_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT78), .B(KEYINPUT37), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n574_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G231gat), .A2(G233gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n289_), .B(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(new_n232_), .ZN(new_n582_));
  XOR2_X1   g381(.A(G127gat), .B(G155gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT16), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G183gat), .B(G211gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT17), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n582_), .A2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n586_), .B(KEYINPUT17), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n589_), .B1(new_n582_), .B2(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n579_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n544_), .A2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT102), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n451_), .A2(new_n456_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n595_), .A2(new_n281_), .A3(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT38), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n575_), .B(KEYINPUT103), .Z(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n601_), .B1(new_n523_), .B2(new_n543_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n307_), .A2(new_n592_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(G1gat), .B1(new_n604_), .B2(new_n596_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n599_), .A2(new_n605_), .ZN(G1324gat));
  INV_X1    g405(.A(new_n391_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n595_), .A2(new_n282_), .A3(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(G8gat), .B1(new_n604_), .B2(new_n391_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT39), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g411(.A(G15gat), .B1(new_n604_), .B2(new_n514_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT41), .Z(new_n614_));
  INV_X1    g413(.A(G15gat), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n595_), .A2(new_n615_), .A3(new_n524_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT104), .Z(G1326gat));
  INV_X1    g417(.A(G22gat), .ZN(new_n619_));
  INV_X1    g418(.A(new_n542_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n595_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(G22gat), .B1(new_n604_), .B2(new_n542_), .ZN(new_n622_));
  XOR2_X1   g421(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n621_), .A2(new_n624_), .ZN(G1327gat));
  INV_X1    g424(.A(new_n307_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n523_), .A2(new_n543_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n592_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n576_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n626_), .A2(new_n627_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(G29gat), .B1(new_n631_), .B2(new_n597_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n491_), .A2(new_n492_), .A3(new_n463_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n462_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n524_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n493_), .A2(new_n520_), .A3(new_n514_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n457_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n541_), .A2(new_n542_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n579_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT43), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT43), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n579_), .B(new_n641_), .C1(new_n637_), .C2(new_n638_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n628_), .B1(new_n640_), .B2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n643_), .A2(KEYINPUT44), .A3(new_n626_), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n644_), .A2(G29gat), .A3(new_n597_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n641_), .B1(new_n627_), .B2(new_n579_), .ZN(new_n646_));
  AOI211_X1 g445(.A(KEYINPUT43), .B(new_n578_), .C1(new_n523_), .C2(new_n543_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n626_), .B(new_n592_), .C1(new_n646_), .C2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n632_), .B1(new_n645_), .B2(new_n650_), .ZN(G1328gat));
  OAI21_X1  g450(.A(new_n607_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n652_));
  AOI21_X1  g451(.A(KEYINPUT44), .B1(new_n643_), .B2(new_n626_), .ZN(new_n653_));
  OAI21_X1  g452(.A(G36gat), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT107), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n391_), .A2(G36gat), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(KEYINPUT45), .B1(new_n630_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT45), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n544_), .A2(new_n659_), .A3(new_n629_), .A4(new_n656_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n654_), .A2(new_n655_), .A3(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n655_), .B1(new_n654_), .B2(new_n661_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT106), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n664_), .A2(KEYINPUT46), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n662_), .A2(new_n663_), .A3(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(G36gat), .ZN(new_n668_));
  AOI211_X1 g467(.A(new_n307_), .B(new_n628_), .C1(new_n640_), .C2(new_n642_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n391_), .B1(new_n669_), .B2(KEYINPUT44), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n668_), .B1(new_n670_), .B2(new_n650_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n661_), .ZN(new_n672_));
  OAI21_X1  g471(.A(KEYINPUT107), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n654_), .A2(new_n655_), .A3(new_n661_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n665_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n667_), .A2(new_n675_), .ZN(G1329gat));
  NAND4_X1  g475(.A1(new_n650_), .A2(new_n644_), .A3(G43gat), .A4(new_n524_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n630_), .A2(new_n514_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n677_), .B1(G43gat), .B2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g479(.A1(new_n630_), .A2(G50gat), .A3(new_n542_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n650_), .A2(new_n644_), .A3(new_n620_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n682_), .A2(KEYINPUT108), .A3(G50gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT108), .B1(new_n682_), .B2(G50gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n681_), .B1(new_n683_), .B2(new_n684_), .ZN(G1331gat));
  INV_X1    g484(.A(new_n280_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n592_), .A2(new_n306_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n602_), .A2(new_n686_), .A3(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(G57gat), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n688_), .A2(new_n689_), .A3(new_n596_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n280_), .A2(new_n306_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n691_), .A2(new_n627_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(new_n593_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n596_), .B1(new_n693_), .B2(KEYINPUT109), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n694_), .B1(KEYINPUT109), .B2(new_n693_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n690_), .B1(new_n695_), .B2(new_n689_), .ZN(G1332gat));
  OAI21_X1  g495(.A(G64gat), .B1(new_n688_), .B2(new_n391_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT48), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n391_), .A2(G64gat), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n698_), .B1(new_n693_), .B2(new_n699_), .ZN(G1333gat));
  OAI21_X1  g499(.A(G71gat), .B1(new_n688_), .B2(new_n514_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT49), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n514_), .A2(G71gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n693_), .B2(new_n703_), .ZN(G1334gat));
  OAI21_X1  g503(.A(G78gat), .B1(new_n688_), .B2(new_n542_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT50), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n542_), .A2(G78gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n706_), .B1(new_n693_), .B2(new_n707_), .ZN(G1335gat));
  NAND2_X1  g507(.A1(new_n643_), .A2(new_n691_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G85gat), .B1(new_n709_), .B2(new_n596_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n692_), .A2(new_n629_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n711_), .A2(new_n212_), .A3(new_n597_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(G1336gat));
  OAI21_X1  g512(.A(G92gat), .B1(new_n709_), .B2(new_n391_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n711_), .A2(new_n213_), .A3(new_n607_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1337gat));
  OAI21_X1  g515(.A(G99gat), .B1(new_n709_), .B2(new_n514_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n711_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n524_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n717_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT51), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n721_), .A2(KEYINPUT110), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n720_), .B(new_n722_), .ZN(G1338gat));
  NAND3_X1  g522(.A1(new_n711_), .A2(new_n206_), .A3(new_n620_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n643_), .A2(new_n620_), .A3(new_n691_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT52), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n725_), .A2(new_n726_), .A3(G106gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n725_), .B2(G106gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n724_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g529(.A(KEYINPUT112), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT55), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n250_), .A2(new_n254_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n262_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n221_), .A2(new_n223_), .A3(new_n249_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n261_), .B1(new_n735_), .B2(new_n231_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n733_), .B1(new_n734_), .B2(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n250_), .B1(new_n734_), .B2(new_n736_), .ZN(new_n738_));
  AOI22_X1  g537(.A1(new_n732_), .A2(new_n737_), .B1(new_n738_), .B2(new_n253_), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n733_), .B(KEYINPUT55), .C1(new_n734_), .C2(new_n736_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n731_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n738_), .A2(new_n253_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n737_), .A2(new_n732_), .ZN(new_n743_));
  AND4_X1   g542(.A1(new_n731_), .A2(new_n742_), .A3(new_n743_), .A4(new_n740_), .ZN(new_n744_));
  OAI211_X1 g543(.A(KEYINPUT56), .B(new_n268_), .C1(new_n741_), .C2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT114), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n250_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n749_));
  OAI22_X1  g548(.A1(KEYINPUT55), .A2(new_n263_), .B1(new_n749_), .B2(new_n254_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n740_), .ZN(new_n751_));
  OAI21_X1  g550(.A(KEYINPUT112), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n742_), .A2(new_n743_), .A3(new_n731_), .A4(new_n740_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n754_), .A2(KEYINPUT114), .A3(KEYINPUT56), .A4(new_n268_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n268_), .B1(new_n741_), .B2(new_n744_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT56), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n747_), .A2(new_n755_), .A3(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n298_), .A2(new_n296_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n760_), .B(new_n302_), .C1(new_n296_), .C2(new_n295_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n305_), .A2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n269_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT113), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT113), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n762_), .A2(new_n765_), .A3(new_n269_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n759_), .A2(KEYINPUT58), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT115), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n759_), .A2(new_n767_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT58), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n759_), .A2(new_n773_), .A3(KEYINPUT58), .A4(new_n767_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n769_), .A2(new_n772_), .A3(new_n579_), .A4(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n306_), .A2(new_n269_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT56), .B1(new_n754_), .B2(new_n268_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n268_), .ZN(new_n779_));
  AOI211_X1 g578(.A(new_n757_), .B(new_n779_), .C1(new_n752_), .C2(new_n753_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n777_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n762_), .A2(new_n271_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT57), .B1(new_n783_), .B2(new_n576_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT57), .ZN(new_n785_));
  AOI211_X1 g584(.A(new_n785_), .B(new_n575_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n784_), .A2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n628_), .B1(new_n775_), .B2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n280_), .A2(new_n578_), .A3(new_n687_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(KEYINPUT111), .B(KEYINPUT54), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n789_), .B(new_n790_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n788_), .A2(new_n791_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n596_), .A2(new_n607_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n522_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n792_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(G113gat), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n796_), .A3(new_n306_), .ZN(new_n797_));
  OR2_X1    g596(.A1(new_n795_), .A2(KEYINPUT59), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n795_), .A2(KEYINPUT59), .ZN(new_n799_));
  AOI22_X1  g598(.A1(new_n798_), .A2(new_n799_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n797_), .B1(new_n800_), .B2(new_n796_), .ZN(G1340gat));
  INV_X1    g600(.A(KEYINPUT60), .ZN(new_n802_));
  INV_X1    g601(.A(G120gat), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n686_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n795_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n280_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(new_n803_), .ZN(G1341gat));
  INV_X1    g607(.A(G127gat), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n795_), .A2(new_n809_), .A3(new_n628_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n592_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n810_), .B1(new_n811_), .B2(new_n809_), .ZN(G1342gat));
  INV_X1    g611(.A(G134gat), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n795_), .A2(new_n813_), .A3(new_n601_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n578_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n814_), .B1(new_n815_), .B2(new_n813_), .ZN(G1343gat));
  NAND2_X1  g615(.A1(new_n793_), .A2(new_n521_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(KEYINPUT116), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n792_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n306_), .ZN(new_n820_));
  XOR2_X1   g619(.A(KEYINPUT117), .B(G141gat), .Z(new_n821_));
  XNOR2_X1  g620(.A(new_n820_), .B(new_n821_), .ZN(G1344gat));
  NAND2_X1  g621(.A1(new_n819_), .A2(new_n686_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g623(.A1(new_n819_), .A2(new_n628_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT118), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n819_), .A2(new_n827_), .A3(new_n628_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(KEYINPUT61), .B(G155gat), .ZN(new_n830_));
  XOR2_X1   g629(.A(new_n830_), .B(KEYINPUT119), .Z(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n829_), .A2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n826_), .A2(new_n828_), .A3(new_n831_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(G1346gat));
  NAND3_X1  g634(.A1(new_n819_), .A2(new_n401_), .A3(new_n601_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n819_), .A2(new_n579_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n836_), .B1(new_n838_), .B2(new_n401_), .ZN(G1347gat));
  INV_X1    g638(.A(new_n791_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n776_), .B1(new_n758_), .B2(new_n745_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n782_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n576_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n785_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n783_), .A2(KEYINPUT57), .A3(new_n576_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n772_), .A2(new_n579_), .A3(new_n774_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n847_), .B2(new_n769_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n840_), .B1(new_n848_), .B2(new_n628_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n596_), .A2(new_n524_), .A3(new_n607_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(KEYINPUT120), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n849_), .A2(KEYINPUT124), .A3(new_n542_), .A4(new_n851_), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n542_), .B(new_n851_), .C1(new_n788_), .C2(new_n791_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT124), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n852_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n364_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n856_), .A2(new_n857_), .A3(new_n306_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT62), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n851_), .A2(new_n860_), .A3(new_n306_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n851_), .B2(new_n306_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n863_), .B(new_n542_), .C1(new_n788_), .C2(new_n791_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n859_), .B1(new_n864_), .B2(G169gat), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(KEYINPUT123), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n864_), .A2(new_n859_), .A3(G169gat), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(KEYINPUT122), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n858_), .B1(new_n866_), .B2(new_n868_), .ZN(G1348gat));
  NOR3_X1   g668(.A1(new_n853_), .A2(new_n317_), .A3(new_n280_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT125), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n853_), .B(KEYINPUT124), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n871_), .B(new_n317_), .C1(new_n872_), .C2(new_n280_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n280_), .B1(new_n852_), .B2(new_n855_), .ZN(new_n874_));
  OAI21_X1  g673(.A(KEYINPUT125), .B1(new_n874_), .B2(G176gat), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n870_), .B1(new_n873_), .B2(new_n875_), .ZN(G1349gat));
  NOR2_X1   g675(.A1(new_n592_), .A2(new_n324_), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n853_), .A2(new_n592_), .ZN(new_n878_));
  AOI22_X1  g677(.A1(new_n856_), .A2(new_n877_), .B1(new_n878_), .B2(new_n309_), .ZN(G1350gat));
  OAI21_X1  g678(.A(G190gat), .B1(new_n872_), .B2(new_n578_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n856_), .A2(new_n601_), .A3(new_n325_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1351gat));
  NAND3_X1  g681(.A1(new_n521_), .A2(new_n596_), .A3(new_n607_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n792_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n306_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n686_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n888_));
  XOR2_X1   g687(.A(new_n887_), .B(new_n888_), .Z(G1353gat));
  NAND2_X1  g688(.A1(new_n884_), .A2(new_n628_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n890_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n891_));
  XOR2_X1   g690(.A(KEYINPUT63), .B(G211gat), .Z(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n890_), .B2(new_n892_), .ZN(G1354gat));
  NAND2_X1  g692(.A1(new_n884_), .A2(new_n579_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(G218gat), .ZN(new_n895_));
  INV_X1    g694(.A(G218gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n884_), .A2(new_n896_), .A3(new_n601_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT127), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n895_), .A2(KEYINPUT127), .A3(new_n897_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(G1355gat));
endmodule


