//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_;
  XOR2_X1   g000(.A(G211gat), .B(G218gat), .Z(new_n202_));
  INV_X1    g001(.A(KEYINPUT21), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204_));
  AOI21_X1  g003(.A(new_n202_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n204_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT21), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n202_), .A3(KEYINPUT21), .ZN(new_n209_));
  AND2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  AND2_X1   g009(.A1(G228gat), .A2(G233gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT91), .B(KEYINPUT2), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT89), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT89), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(G141gat), .A3(G148gat), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n217_), .B1(new_n219_), .B2(new_n221_), .ZN(new_n222_));
  OR3_X1    g021(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT92), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND4_X1  g025(.A1(KEYINPUT92), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n223_), .A2(new_n226_), .A3(new_n227_), .A4(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n216_), .B1(new_n222_), .B2(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n213_), .B1(new_n215_), .B2(KEYINPUT1), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n231_), .B1(KEYINPUT1), .B2(new_n213_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT90), .ZN(new_n233_));
  INV_X1    g032(.A(G141gat), .ZN(new_n234_));
  INV_X1    g033(.A(G148gat), .ZN(new_n235_));
  AOI22_X1  g034(.A1(new_n219_), .A2(new_n221_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n232_), .A2(new_n233_), .A3(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n233_), .B1(new_n232_), .B2(new_n236_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n230_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT93), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT93), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n242_), .B(new_n230_), .C1(new_n238_), .C2(new_n239_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT29), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n212_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n247_));
  NAND2_X1  g046(.A1(new_n240_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n208_), .A2(new_n209_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(new_n211_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G78gat), .B(G106gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n252_), .B(KEYINPUT96), .Z(new_n253_));
  AND3_X1   g052(.A1(new_n246_), .A2(new_n251_), .A3(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n253_), .B1(new_n246_), .B2(new_n251_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n244_), .A2(new_n245_), .ZN(new_n257_));
  XOR2_X1   g056(.A(KEYINPUT94), .B(KEYINPUT28), .Z(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(G22gat), .B(G50gat), .Z(new_n260_));
  INV_X1    g059(.A(new_n258_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n244_), .A2(new_n245_), .A3(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n259_), .A2(new_n260_), .A3(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n260_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n261_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n265_));
  AOI211_X1 g064(.A(KEYINPUT29), .B(new_n258_), .C1(new_n241_), .C2(new_n243_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n264_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n263_), .A2(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT97), .B1(new_n256_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n246_), .A2(new_n251_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n253_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n246_), .A2(new_n251_), .A3(new_n253_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT97), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n274_), .A2(new_n275_), .A3(new_n263_), .A4(new_n267_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n269_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n270_), .A2(new_n252_), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n278_), .A2(new_n273_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n268_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n277_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT24), .ZN(new_n282_));
  INV_X1    g081(.A(G169gat), .ZN(new_n283_));
  INV_X1    g082(.A(G176gat), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n283_), .A2(new_n284_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n285_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT25), .B(G183gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT26), .B(G190gat), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n288_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT23), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT85), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT23), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n292_), .B(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n294_), .B1(new_n296_), .B2(KEYINPUT85), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n291_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n292_), .B(KEYINPUT23), .ZN(new_n299_));
  OR2_X1    g098(.A1(G183gat), .A2(G190gat), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT22), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n302_));
  OAI21_X1  g101(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT98), .ZN(new_n305_));
  AOI22_X1  g104(.A1(new_n299_), .A2(new_n300_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n302_), .A2(KEYINPUT98), .A3(new_n303_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n298_), .A2(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT99), .B1(new_n309_), .B2(new_n249_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT99), .ZN(new_n311_));
  AOI22_X1  g110(.A1(new_n297_), .A2(new_n291_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n210_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n310_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G226gat), .A2(G233gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT19), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT20), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n288_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n299_), .ZN(new_n320_));
  XOR2_X1   g119(.A(KEYINPUT82), .B(G183gat), .Z(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT25), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT83), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT26), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n323_), .B1(new_n324_), .B2(G190gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(G190gat), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT25), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(G183gat), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n325_), .A2(new_n326_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT84), .ZN(new_n330_));
  INV_X1    g129(.A(G190gat), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n331_), .A2(KEYINPUT83), .A3(KEYINPUT26), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n322_), .A2(new_n329_), .A3(new_n330_), .A4(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT82), .B(G183gat), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n334_), .A2(new_n327_), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n325_), .A2(new_n332_), .A3(new_n326_), .A4(new_n328_), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT84), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n320_), .B1(new_n333_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n321_), .A2(new_n331_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n304_), .B1(new_n297_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n339_), .A2(KEYINPUT86), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT86), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n344_), .B1(new_n338_), .B2(new_n341_), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n314_), .B(new_n318_), .C1(new_n346_), .C2(new_n210_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n343_), .A2(new_n210_), .A3(new_n345_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n317_), .B1(new_n309_), .B2(new_n249_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n316_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G8gat), .B(G36gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT18), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G64gat), .B(G92gat), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n353_), .B(new_n354_), .Z(new_n355_));
  NAND3_X1  g154(.A1(new_n347_), .A2(new_n351_), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n210_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT102), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n309_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n312_), .A2(KEYINPUT102), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n359_), .A2(new_n360_), .A3(new_n210_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT20), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n316_), .B1(new_n357_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n316_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n348_), .A2(new_n364_), .A3(new_n349_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n355_), .ZN(new_n367_));
  AOI21_X1  g166(.A(KEYINPUT103), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT103), .ZN(new_n369_));
  AOI211_X1 g168(.A(new_n369_), .B(new_n355_), .C1(new_n363_), .C2(new_n365_), .ZN(new_n370_));
  OAI211_X1 g169(.A(KEYINPUT27), .B(new_n356_), .C1(new_n368_), .C2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n314_), .A2(new_n318_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n372_), .A2(new_n357_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n364_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n367_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT100), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n356_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT27), .ZN(new_n378_));
  OAI211_X1 g177(.A(KEYINPUT100), .B(new_n367_), .C1(new_n373_), .C2(new_n374_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n377_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n371_), .A2(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n281_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT4), .ZN(new_n383_));
  XOR2_X1   g182(.A(G127gat), .B(G134gat), .Z(new_n384_));
  XNOR2_X1  g183(.A(G113gat), .B(G120gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n241_), .A2(new_n243_), .A3(new_n386_), .ZN(new_n387_));
  OR2_X1    g186(.A1(new_n240_), .A2(new_n386_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n383_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G225gat), .A2(G233gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT101), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n387_), .A2(new_n383_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n390_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n392_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G1gat), .B(G29gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(G85gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT0), .B(G57gat), .ZN(new_n400_));
  XOR2_X1   g199(.A(new_n399_), .B(new_n400_), .Z(new_n401_));
  NAND2_X1  g200(.A1(new_n397_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n401_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n394_), .A2(new_n403_), .A3(new_n396_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G71gat), .B(G99gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(G43gat), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n343_), .A2(new_n345_), .A3(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n408_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G227gat), .A2(G233gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(G15gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(KEYINPUT30), .ZN(new_n413_));
  OR3_X1    g212(.A1(new_n409_), .A2(new_n410_), .A3(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n413_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(KEYINPUT88), .B1(new_n416_), .B2(KEYINPUT87), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n386_), .B(KEYINPUT31), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n416_), .A2(KEYINPUT88), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n418_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n420_), .B1(new_n417_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n382_), .A2(new_n406_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n355_), .A2(KEYINPUT32), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n347_), .A2(new_n351_), .A3(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n366_), .A2(KEYINPUT32), .A3(new_n355_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n405_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n377_), .A2(new_n379_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT33), .ZN(new_n431_));
  INV_X1    g230(.A(new_n393_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n432_), .A2(new_n389_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n395_), .B1(new_n433_), .B2(new_n392_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n431_), .B1(new_n434_), .B2(new_n403_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n397_), .A2(KEYINPUT33), .A3(new_n401_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n387_), .A2(new_n388_), .A3(new_n392_), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n403_), .B(new_n437_), .C1(new_n433_), .C2(new_n392_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n430_), .A2(new_n435_), .A3(new_n436_), .A4(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n429_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n281_), .ZN(new_n441_));
  AND2_X1   g240(.A1(new_n371_), .A2(new_n380_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n405_), .B1(new_n277_), .B2(new_n280_), .ZN(new_n443_));
  AOI22_X1  g242(.A1(new_n440_), .A2(new_n441_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n425_), .B1(new_n444_), .B2(new_n424_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT81), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G113gat), .B(G141gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G169gat), .B(G197gat), .ZN(new_n448_));
  XOR2_X1   g247(.A(new_n447_), .B(new_n448_), .Z(new_n449_));
  NAND2_X1  g248(.A1(G229gat), .A2(G233gat), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G1gat), .B(G8gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT76), .B(G15gat), .ZN(new_n453_));
  INV_X1    g252(.A(G22gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT77), .B(G8gat), .ZN(new_n456_));
  INV_X1    g255(.A(G1gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT14), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n452_), .B1(new_n455_), .B2(new_n458_), .ZN(new_n459_));
  XOR2_X1   g258(.A(KEYINPUT76), .B(G15gat), .Z(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n454_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n453_), .A2(G22gat), .ZN(new_n462_));
  AND4_X1   g261(.A1(new_n458_), .A2(new_n461_), .A3(new_n462_), .A4(new_n452_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G29gat), .B(G36gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G43gat), .B(G50gat), .ZN(new_n465_));
  OR2_X1    g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n465_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n459_), .A2(new_n463_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n468_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n452_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n461_), .A2(new_n462_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n458_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n471_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n455_), .A2(new_n458_), .A3(new_n452_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n470_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n451_), .B1(new_n469_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT80), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n468_), .B1(new_n459_), .B2(new_n463_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n474_), .A2(new_n475_), .A3(new_n470_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT80), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n481_), .A2(new_n482_), .A3(new_n451_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n478_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT15), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n468_), .A2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n466_), .A2(KEYINPUT15), .A3(new_n467_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n474_), .A2(new_n486_), .A3(new_n475_), .A4(new_n487_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n488_), .A2(new_n479_), .A3(new_n450_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n449_), .B1(new_n484_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n449_), .ZN(new_n492_));
  AOI211_X1 g291(.A(new_n489_), .B(new_n492_), .C1(new_n478_), .C2(new_n483_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n446_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n482_), .B1(new_n481_), .B2(new_n451_), .ZN(new_n495_));
  AOI211_X1 g294(.A(KEYINPUT80), .B(new_n450_), .C1(new_n479_), .C2(new_n480_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n490_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(new_n492_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n484_), .A2(new_n490_), .A3(new_n449_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n498_), .A2(new_n499_), .A3(KEYINPUT81), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n494_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n445_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G57gat), .B(G64gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G71gat), .B(G78gat), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n505_), .A3(KEYINPUT11), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(KEYINPUT11), .ZN(new_n507_));
  INV_X1    g306(.A(new_n505_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n504_), .A2(KEYINPUT11), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n506_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT12), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G85gat), .B(G92gat), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n514_), .A2(KEYINPUT64), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT9), .ZN(new_n516_));
  XOR2_X1   g315(.A(KEYINPUT10), .B(G99gat), .Z(new_n517_));
  INV_X1    g316(.A(G106gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(G85gat), .ZN(new_n520_));
  INV_X1    g319(.A(G92gat), .ZN(new_n521_));
  AOI21_X1  g320(.A(KEYINPUT9), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n522_), .B1(new_n514_), .B2(KEYINPUT64), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G99gat), .A2(G106gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT6), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT6), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n526_), .A2(G99gat), .A3(G106gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n516_), .A2(new_n519_), .A3(new_n523_), .A4(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT65), .ZN(new_n531_));
  INV_X1    g330(.A(G99gat), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(new_n532_), .A3(new_n518_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT7), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT7), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n531_), .A2(new_n535_), .A3(new_n532_), .A4(new_n518_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n534_), .A2(new_n528_), .A3(new_n536_), .ZN(new_n537_));
  AND2_X1   g336(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n514_), .A2(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n530_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n537_), .A2(new_n530_), .A3(new_n539_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n513_), .B1(new_n529_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  AND3_X1   g344(.A1(new_n537_), .A2(new_n530_), .A3(new_n539_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n529_), .B1(new_n546_), .B2(new_n540_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT67), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n529_), .B(KEYINPUT67), .C1(new_n546_), .C2(new_n540_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n511_), .A2(KEYINPUT68), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT68), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n552_), .B(new_n506_), .C1(new_n509_), .C2(new_n510_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n549_), .A2(new_n550_), .A3(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G230gat), .A2(G233gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n554_), .ZN(new_n559_));
  AOI21_X1  g358(.A(KEYINPUT67), .B1(new_n543_), .B2(new_n529_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n550_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n559_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(KEYINPUT71), .B1(new_n562_), .B2(new_n512_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n554_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT71), .ZN(new_n565_));
  NOR3_X1   g364(.A1(new_n564_), .A2(new_n565_), .A3(KEYINPUT12), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n545_), .B(new_n558_), .C1(new_n563_), .C2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G120gat), .B(G148gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT5), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G176gat), .B(G204gat), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n569_), .B(new_n570_), .Z(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n555_), .A2(KEYINPUT69), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT70), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT69), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n549_), .A2(new_n575_), .A3(new_n550_), .A4(new_n554_), .ZN(new_n576_));
  AND3_X1   g375(.A1(new_n573_), .A2(new_n574_), .A3(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n574_), .B1(new_n573_), .B2(new_n576_), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n577_), .A2(new_n578_), .A3(new_n564_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n567_), .B(new_n572_), .C1(new_n579_), .C2(new_n556_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT72), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n573_), .A2(new_n576_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT70), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n573_), .A2(new_n574_), .A3(new_n576_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n583_), .A2(new_n584_), .A3(new_n562_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n556_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT72), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n587_), .A2(new_n588_), .A3(new_n567_), .A4(new_n572_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n581_), .A2(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n564_), .B1(new_n582_), .B2(KEYINPUT70), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n556_), .B1(new_n591_), .B2(new_n584_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n562_), .A2(KEYINPUT71), .A3(new_n512_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n565_), .B1(new_n564_), .B2(KEYINPUT12), .ZN(new_n594_));
  AOI211_X1 g393(.A(new_n544_), .B(new_n557_), .C1(new_n593_), .C2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n571_), .B1(new_n592_), .B2(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n597_));
  NOR2_X1   g396(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n590_), .B(new_n596_), .C1(new_n597_), .C2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n590_), .A2(new_n596_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n599_), .B1(new_n601_), .B2(new_n598_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT37), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n549_), .A2(new_n468_), .A3(new_n550_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n547_), .A2(new_n487_), .A3(new_n486_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n606_));
  NAND2_X1  g405(.A1(G232gat), .A2(G233gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n604_), .B(new_n605_), .C1(KEYINPUT35), .C2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(KEYINPUT35), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n609_), .B(new_n610_), .Z(new_n611_));
  INV_X1    g410(.A(KEYINPUT75), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G190gat), .B(G218gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G134gat), .B(G162gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT36), .Z(new_n616_));
  NAND3_X1  g415(.A1(new_n611_), .A2(new_n612_), .A3(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n609_), .B(new_n610_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n615_), .A2(KEYINPUT36), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n612_), .B1(new_n611_), .B2(new_n616_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n603_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n474_), .A2(new_n475_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G231gat), .A2(G233gat), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n624_), .B(new_n625_), .Z(new_n626_));
  AND2_X1   g425(.A1(new_n626_), .A2(new_n511_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT17), .ZN(new_n628_));
  XOR2_X1   g427(.A(G127gat), .B(G155gat), .Z(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT79), .ZN(new_n630_));
  XOR2_X1   g429(.A(G183gat), .B(G211gat), .Z(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  XOR2_X1   g431(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n627_), .A2(new_n628_), .A3(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n635_), .B1(new_n511_), .B2(new_n626_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n634_), .B(KEYINPUT17), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n626_), .A2(new_n559_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n626_), .A2(new_n559_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n637_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n636_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n611_), .A2(new_n616_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n643_), .A2(KEYINPUT37), .A3(new_n620_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n623_), .A2(new_n642_), .A3(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n602_), .A2(new_n646_), .ZN(new_n647_));
  OR3_X1    g446(.A1(new_n503_), .A2(new_n647_), .A3(KEYINPUT104), .ZN(new_n648_));
  OAI21_X1  g447(.A(KEYINPUT104), .B1(new_n503_), .B2(new_n647_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n648_), .A2(new_n457_), .A3(new_n405_), .A4(new_n649_), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n650_), .A2(KEYINPUT105), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(KEYINPUT105), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT38), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n621_), .A2(new_n622_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n656_), .A2(new_n641_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n445_), .A2(new_n502_), .A3(new_n602_), .A4(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G1gat), .B1(new_n658_), .B2(new_n406_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n651_), .A2(KEYINPUT38), .A3(new_n652_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n655_), .A2(new_n659_), .A3(new_n660_), .ZN(G1324gat));
  AND2_X1   g460(.A1(new_n381_), .A2(new_n456_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n648_), .A2(new_n649_), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT106), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n648_), .A2(KEYINPUT106), .A3(new_n649_), .A4(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G8gat), .B1(new_n658_), .B2(new_n442_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT39), .ZN(new_n669_));
  XNOR2_X1  g468(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n667_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n667_), .B2(new_n669_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1325gat));
  AND2_X1   g472(.A1(new_n648_), .A2(new_n649_), .ZN(new_n674_));
  INV_X1    g473(.A(G15gat), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n674_), .A2(new_n675_), .A3(new_n424_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT108), .ZN(new_n677_));
  OAI21_X1  g476(.A(G15gat), .B1(new_n658_), .B2(new_n423_), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT41), .Z(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(G1326gat));
  NAND3_X1  g479(.A1(new_n674_), .A2(new_n454_), .A3(new_n281_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G22gat), .B1(new_n658_), .B2(new_n441_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT42), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(G1327gat));
  INV_X1    g483(.A(new_n602_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n685_), .A2(new_n501_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n623_), .A2(new_n644_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n445_), .A2(new_n687_), .A3(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n687_), .B1(new_n445_), .B2(new_n688_), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n641_), .B(new_n686_), .C1(new_n689_), .C2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n445_), .A2(new_n688_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT43), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n445_), .A2(new_n687_), .A3(new_n688_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n697_), .A2(KEYINPUT44), .A3(new_n641_), .A4(new_n686_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n693_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(G29gat), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n699_), .A2(new_n700_), .A3(new_n406_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n656_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n702_), .A2(new_n642_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n503_), .A2(new_n685_), .A3(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(G29gat), .B1(new_n705_), .B2(new_n405_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n701_), .A2(new_n706_), .ZN(G1328gat));
  NAND3_X1  g506(.A1(new_n693_), .A2(new_n698_), .A3(new_n381_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(G36gat), .ZN(new_n709_));
  INV_X1    g508(.A(G36gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n705_), .A2(new_n710_), .A3(new_n381_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT45), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n709_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT46), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n709_), .A2(KEYINPUT46), .A3(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1329gat));
  NAND2_X1  g516(.A1(new_n424_), .A2(G43gat), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n705_), .A2(new_n424_), .ZN(new_n719_));
  OAI22_X1  g518(.A1(new_n699_), .A2(new_n718_), .B1(G43gat), .B2(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g520(.A(G50gat), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n699_), .A2(new_n722_), .A3(new_n441_), .ZN(new_n723_));
  AOI21_X1  g522(.A(G50gat), .B1(new_n705_), .B2(new_n281_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1331gat));
  NAND2_X1  g524(.A1(new_n445_), .A2(new_n501_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT109), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n727_), .A2(new_n602_), .A3(new_n645_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n405_), .ZN(new_n729_));
  INV_X1    g528(.A(G57gat), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT110), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n729_), .A2(new_n733_), .A3(new_n730_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n685_), .A2(new_n501_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n445_), .A2(new_n657_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n406_), .A2(new_n730_), .ZN(new_n738_));
  AOI22_X1  g537(.A1(new_n732_), .A2(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(G1332gat));
  INV_X1    g538(.A(G64gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n737_), .B2(new_n381_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT48), .Z(new_n742_));
  NAND3_X1  g541(.A1(new_n728_), .A2(new_n740_), .A3(new_n381_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1333gat));
  INV_X1    g543(.A(G71gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n737_), .B2(new_n424_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT49), .Z(new_n747_));
  NAND3_X1  g546(.A1(new_n728_), .A2(new_n745_), .A3(new_n424_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1334gat));
  INV_X1    g548(.A(G78gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n750_), .B1(new_n737_), .B2(new_n281_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n751_), .B(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n728_), .A2(new_n750_), .A3(new_n281_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1335gat));
  NOR3_X1   g554(.A1(new_n727_), .A2(new_n602_), .A3(new_n704_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n756_), .A2(new_n520_), .A3(new_n405_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n735_), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n758_), .B(new_n641_), .C1(new_n689_), .C2(new_n690_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT112), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT112), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n697_), .A2(new_n761_), .A3(new_n641_), .A4(new_n758_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n760_), .A2(new_n762_), .A3(KEYINPUT113), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT113), .B1(new_n760_), .B2(new_n762_), .ZN(new_n764_));
  NOR3_X1   g563(.A1(new_n763_), .A2(new_n764_), .A3(new_n406_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n757_), .B1(new_n765_), .B2(new_n520_), .ZN(G1336gat));
  NAND3_X1  g565(.A1(new_n756_), .A2(new_n521_), .A3(new_n381_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n763_), .A2(new_n764_), .A3(new_n442_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(new_n521_), .ZN(G1337gat));
  NAND3_X1  g568(.A1(new_n756_), .A2(new_n424_), .A3(new_n517_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n423_), .B1(new_n760_), .B2(new_n762_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(new_n532_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT51), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n770_), .B(new_n774_), .C1(new_n771_), .C2(new_n532_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1338gat));
  NAND3_X1  g575(.A1(new_n756_), .A2(new_n518_), .A3(new_n281_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n778_), .B(G106gat), .C1(new_n759_), .C2(new_n441_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n697_), .A2(new_n281_), .A3(new_n641_), .A4(new_n758_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n778_), .B1(new_n781_), .B2(G106gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n777_), .B1(new_n780_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT53), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n777_), .B(new_n785_), .C1(new_n780_), .C2(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1339gat));
  NAND3_X1  g586(.A1(new_n382_), .A2(new_n405_), .A3(new_n424_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n623_), .A2(new_n644_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n567_), .A2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n544_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n792_), .A2(KEYINPUT55), .A3(new_n558_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n582_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n556_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n791_), .B(new_n793_), .C1(new_n795_), .C2(new_n796_), .ZN(new_n797_));
  AOI211_X1 g596(.A(KEYINPUT115), .B(new_n556_), .C1(new_n792_), .C2(new_n794_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n571_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT56), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT56), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n801_), .B(new_n571_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n481_), .A2(new_n450_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n488_), .A2(new_n479_), .A3(new_n451_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(new_n492_), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n499_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n806_), .B1(new_n581_), .B2(new_n589_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n800_), .A2(new_n802_), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT58), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n789_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n800_), .A2(KEYINPUT58), .A3(new_n802_), .A4(new_n807_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n806_), .B1(new_n590_), .B2(new_n596_), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n799_), .A2(KEYINPUT116), .A3(KEYINPUT56), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT56), .B1(new_n799_), .B2(KEYINPUT116), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT114), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n817_), .B1(new_n590_), .B2(new_n502_), .ZN(new_n818_));
  AOI211_X1 g617(.A(KEYINPUT114), .B(new_n501_), .C1(new_n581_), .C2(new_n589_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n813_), .B1(new_n816_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n656_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n812_), .B1(new_n821_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n799_), .A2(KEYINPUT116), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n801_), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n585_), .A2(new_n586_), .B1(new_n792_), .B2(new_n558_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n588_), .B1(new_n828_), .B2(new_n572_), .ZN(new_n829_));
  NOR4_X1   g628(.A1(new_n592_), .A2(new_n595_), .A3(KEYINPUT72), .A4(new_n571_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n502_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT114), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n590_), .A2(new_n817_), .A3(new_n502_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n799_), .A2(KEYINPUT116), .A3(KEYINPUT56), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n827_), .A2(new_n832_), .A3(new_n833_), .A4(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n813_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(KEYINPUT57), .B1(new_n837_), .B2(new_n702_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n641_), .B1(new_n825_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n840_));
  AND4_X1   g639(.A1(new_n840_), .A2(new_n602_), .A3(new_n646_), .A4(new_n501_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n600_), .B1(KEYINPUT73), .B2(KEYINPUT13), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n645_), .B1(new_n842_), .B2(new_n599_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n840_), .B1(new_n843_), .B2(new_n501_), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n841_), .A2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n788_), .B1(new_n839_), .B2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(G113gat), .B1(new_n846_), .B2(new_n502_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n848_));
  INV_X1    g647(.A(new_n788_), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n837_), .A2(new_n823_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n822_), .B1(new_n821_), .B2(new_n656_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n642_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n841_), .A2(new_n844_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n848_), .B(new_n849_), .C1(new_n852_), .C2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(KEYINPUT117), .B1(new_n846_), .B2(new_n848_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT117), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n850_), .A2(new_n851_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n853_), .B1(new_n858_), .B2(new_n641_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n857_), .B(KEYINPUT59), .C1(new_n859_), .C2(new_n788_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n855_), .B1(new_n856_), .B2(new_n860_), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n502_), .A2(G113gat), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n847_), .B1(new_n861_), .B2(new_n862_), .ZN(G1340gat));
  INV_X1    g662(.A(KEYINPUT60), .ZN(new_n864_));
  AOI21_X1  g663(.A(G120gat), .B1(new_n685_), .B2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT118), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n867_), .B1(new_n864_), .B2(G120gat), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n846_), .B(new_n866_), .C1(new_n865_), .C2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n854_), .A2(new_n685_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(new_n856_), .B2(new_n860_), .ZN(new_n871_));
  INV_X1    g670(.A(G120gat), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n869_), .B1(new_n871_), .B2(new_n872_), .ZN(G1341gat));
  AOI21_X1  g672(.A(G127gat), .B1(new_n846_), .B2(new_n642_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n642_), .A2(G127gat), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n861_), .B2(new_n875_), .ZN(G1342gat));
  AOI21_X1  g675(.A(G134gat), .B1(new_n846_), .B2(new_n656_), .ZN(new_n877_));
  XOR2_X1   g676(.A(KEYINPUT119), .B(G134gat), .Z(new_n878_));
  NOR2_X1   g677(.A1(new_n789_), .A2(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n877_), .B1(new_n861_), .B2(new_n879_), .ZN(G1343gat));
  NAND2_X1  g679(.A1(new_n839_), .A2(new_n845_), .ZN(new_n881_));
  NOR4_X1   g680(.A1(new_n424_), .A2(new_n441_), .A3(new_n406_), .A4(new_n381_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(new_n501_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(new_n234_), .ZN(G1344gat));
  NOR2_X1   g684(.A1(new_n883_), .A2(new_n602_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(new_n235_), .ZN(G1345gat));
  OAI211_X1 g686(.A(new_n642_), .B(new_n882_), .C1(new_n852_), .C2(new_n853_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(KEYINPUT120), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n881_), .A2(new_n890_), .A3(new_n642_), .A4(new_n882_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT61), .B(G155gat), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n889_), .A2(new_n891_), .A3(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n889_), .B2(new_n891_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1346gat));
  OAI21_X1  g694(.A(G162gat), .B1(new_n883_), .B2(new_n789_), .ZN(new_n896_));
  OR2_X1    g695(.A1(new_n702_), .A2(G162gat), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n883_), .B2(new_n897_), .ZN(G1347gat));
  NOR3_X1   g697(.A1(new_n442_), .A2(new_n423_), .A3(new_n405_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n502_), .ZN(new_n900_));
  XOR2_X1   g699(.A(new_n900_), .B(KEYINPUT121), .Z(new_n901_));
  NAND3_X1  g700(.A1(new_n881_), .A2(new_n441_), .A3(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT62), .ZN(new_n903_));
  AND3_X1   g702(.A1(new_n902_), .A2(new_n903_), .A3(G169gat), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n903_), .B1(new_n902_), .B2(G169gat), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n881_), .A2(new_n441_), .A3(new_n899_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT22), .B(G169gat), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n502_), .A2(new_n907_), .ZN(new_n908_));
  OAI22_X1  g707(.A1(new_n904_), .A2(new_n905_), .B1(new_n906_), .B2(new_n908_), .ZN(G1348gat));
  XOR2_X1   g708(.A(KEYINPUT122), .B(G176gat), .Z(new_n910_));
  OR3_X1    g709(.A1(new_n906_), .A2(new_n602_), .A3(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n906_), .B2(new_n602_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1349gat));
  NOR3_X1   g712(.A1(new_n906_), .A2(new_n289_), .A3(new_n641_), .ZN(new_n914_));
  OR2_X1    g713(.A1(new_n906_), .A2(new_n641_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n914_), .B1(new_n321_), .B2(new_n915_), .ZN(G1350gat));
  OAI21_X1  g715(.A(G190gat), .B1(new_n906_), .B2(new_n789_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n656_), .A2(new_n290_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n906_), .B2(new_n918_), .ZN(G1351gat));
  INV_X1    g718(.A(new_n443_), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n920_), .A2(new_n424_), .A3(new_n442_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n859_), .A2(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n502_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g724(.A1(new_n881_), .A2(new_n921_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n927_));
  OAI22_X1  g726(.A1(new_n926_), .A2(new_n602_), .B1(new_n927_), .B2(G204gat), .ZN(new_n928_));
  XOR2_X1   g727(.A(KEYINPUT123), .B(G204gat), .Z(new_n929_));
  NAND3_X1  g728(.A1(new_n923_), .A2(new_n685_), .A3(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n928_), .A2(new_n930_), .ZN(G1353gat));
  AOI21_X1  g730(.A(new_n641_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n881_), .A2(new_n921_), .A3(new_n932_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(KEYINPUT125), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n933_), .A2(new_n937_), .A3(new_n934_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT124), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n939_), .B1(new_n933_), .B2(new_n934_), .ZN(new_n940_));
  INV_X1    g739(.A(new_n934_), .ZN(new_n941_));
  NAND4_X1  g740(.A1(new_n923_), .A2(KEYINPUT124), .A3(new_n941_), .A4(new_n932_), .ZN(new_n942_));
  AOI22_X1  g741(.A1(new_n936_), .A2(new_n938_), .B1(new_n940_), .B2(new_n942_), .ZN(G1354gat));
  XNOR2_X1  g742(.A(KEYINPUT127), .B(G218gat), .ZN(new_n944_));
  NOR3_X1   g743(.A1(new_n926_), .A2(new_n789_), .A3(new_n944_), .ZN(new_n945_));
  INV_X1    g744(.A(KEYINPUT126), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n946_), .B1(new_n926_), .B2(new_n702_), .ZN(new_n947_));
  NAND4_X1  g746(.A1(new_n881_), .A2(KEYINPUT126), .A3(new_n656_), .A4(new_n921_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(new_n948_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n945_), .B1(new_n949_), .B2(new_n944_), .ZN(G1355gat));
endmodule


