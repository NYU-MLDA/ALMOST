//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 1 0 1 0 1 1 1 1 0 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n588_,
    new_n589_, new_n590_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n782_, new_n783_,
    new_n784_, new_n786_, new_n787_, new_n789_, new_n790_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n811_, new_n813_, new_n815_, new_n816_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n824_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n831_, new_n832_,
    new_n833_, new_n834_;
  INV_X1    g000(.A(KEYINPUT22), .ZN(new_n202_));
  INV_X1    g001(.A(G169gat), .ZN(new_n203_));
  NOR3_X1   g002(.A1(new_n202_), .A2(new_n203_), .A3(KEYINPUT80), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(G176gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT80), .B1(new_n203_), .B2(KEYINPUT81), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n206_), .A2(new_n202_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n202_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n205_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n211_), .A2(KEYINPUT23), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT79), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n211_), .B(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n212_), .B1(new_n214_), .B2(KEYINPUT23), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n209_), .B(new_n210_), .C1(new_n215_), .C2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n211_), .A2(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n219_), .B1(new_n214_), .B2(new_n218_), .ZN(new_n220_));
  INV_X1    g019(.A(G176gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n203_), .A2(new_n221_), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n222_), .A2(KEYINPUT24), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT77), .ZN(new_n224_));
  INV_X1    g023(.A(G190gat), .ZN(new_n225_));
  NOR3_X1   g024(.A1(new_n224_), .A2(new_n225_), .A3(KEYINPUT26), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT25), .B(G183gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT26), .B1(new_n224_), .B2(new_n225_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n220_), .B(new_n223_), .C1(new_n226_), .C2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n222_), .A2(KEYINPUT24), .A3(new_n210_), .ZN(new_n231_));
  XOR2_X1   g030(.A(new_n231_), .B(KEYINPUT78), .Z(new_n232_));
  OAI21_X1  g031(.A(new_n217_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G227gat), .A2(G233gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(KEYINPUT31), .B(G43gat), .Z(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G113gat), .B(G120gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT82), .ZN(new_n239_));
  XOR2_X1   g038(.A(G127gat), .B(G134gat), .Z(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XOR2_X1   g040(.A(KEYINPUT30), .B(G15gat), .Z(new_n242_));
  XNOR2_X1  g041(.A(G71gat), .B(G99gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n241_), .B(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n237_), .B(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(G155gat), .A2(G162gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT83), .ZN(new_n248_));
  INV_X1    g047(.A(G155gat), .ZN(new_n249_));
  INV_X1    g048(.A(G162gat), .ZN(new_n250_));
  INV_X1    g049(.A(G141gat), .ZN(new_n251_));
  INV_X1    g050(.A(G148gat), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  OR2_X1    g052(.A1(KEYINPUT85), .A2(KEYINPUT2), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT84), .ZN(new_n255_));
  AOI22_X1  g054(.A1(new_n253_), .A2(new_n254_), .B1(new_n255_), .B2(KEYINPUT3), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n251_), .A2(new_n252_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n257_), .B1(new_n255_), .B2(KEYINPUT3), .ZN(new_n258_));
  OR4_X1    g057(.A1(new_n255_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n256_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(KEYINPUT85), .A2(KEYINPUT2), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n253_), .B1(new_n254_), .B2(new_n261_), .ZN(new_n262_));
  OAI221_X1 g061(.A(new_n248_), .B1(new_n249_), .B2(new_n250_), .C1(new_n260_), .C2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT1), .B1(new_n249_), .B2(new_n250_), .ZN(new_n264_));
  OR3_X1    g063(.A1(new_n249_), .A2(new_n250_), .A3(KEYINPUT1), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n248_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n253_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n266_), .A2(new_n257_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n263_), .A2(new_n268_), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n269_), .A2(new_n241_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n241_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n270_), .A2(KEYINPUT4), .A3(new_n271_), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n271_), .A2(KEYINPUT4), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G225gat), .A2(G233gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n274_), .B(KEYINPUT94), .Z(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n272_), .A2(new_n273_), .A3(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n270_), .A2(new_n271_), .A3(new_n274_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G1gat), .B(G29gat), .ZN(new_n280_));
  INV_X1    g079(.A(G85gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT0), .B(G57gat), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n282_), .B(new_n283_), .Z(new_n284_));
  NAND2_X1  g083(.A1(new_n279_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n284_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n277_), .A2(new_n278_), .A3(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  AOI211_X1 g087(.A(new_n216_), .B(new_n219_), .C1(new_n214_), .C2(new_n218_), .ZN(new_n289_));
  XOR2_X1   g088(.A(KEYINPUT22), .B(G169gat), .Z(new_n290_));
  OAI21_X1  g089(.A(new_n210_), .B1(new_n290_), .B2(G176gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT26), .B(G190gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n227_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(new_n223_), .A3(new_n231_), .ZN(new_n294_));
  OAI22_X1  g093(.A1(new_n289_), .A2(new_n291_), .B1(new_n215_), .B2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G211gat), .B(G218gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT89), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G197gat), .B(G204gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT21), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n299_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n297_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n296_), .A2(KEYINPUT89), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n296_), .A2(KEYINPUT89), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(new_n300_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n295_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT90), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n307_), .B(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n308_), .B1(new_n310_), .B2(new_n233_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G226gat), .A2(G233gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT19), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n311_), .A2(KEYINPUT20), .A3(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(G64gat), .B(G92gat), .Z(new_n316_));
  XNOR2_X1  g115(.A(G8gat), .B(G36gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n318_), .B(new_n319_), .Z(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT32), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n295_), .A2(new_n307_), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n322_), .B(KEYINPUT20), .C1(new_n310_), .C2(new_n233_), .ZN(new_n323_));
  AND3_X1   g122(.A1(new_n323_), .A2(KEYINPUT92), .A3(new_n313_), .ZN(new_n324_));
  AOI21_X1  g123(.A(KEYINPUT92), .B1(new_n323_), .B2(new_n313_), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n315_), .B(new_n321_), .C1(new_n324_), .C2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT97), .B(KEYINPUT20), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n314_), .B1(new_n311_), .B2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n323_), .A2(new_n313_), .ZN(new_n329_));
  OAI211_X1 g128(.A(KEYINPUT32), .B(new_n320_), .C1(new_n328_), .C2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n288_), .A2(new_n326_), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT98), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT98), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n288_), .A2(new_n326_), .A3(new_n330_), .A4(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n315_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n320_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n320_), .B(new_n315_), .C1(new_n324_), .C2(new_n325_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(KEYINPUT95), .A2(KEYINPUT33), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n287_), .A2(new_n340_), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n287_), .A2(new_n340_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n270_), .A2(new_n271_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n284_), .B1(new_n343_), .B2(new_n275_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT96), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n272_), .A2(new_n274_), .A3(new_n273_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n344_), .A2(new_n345_), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n341_), .B(new_n342_), .C1(new_n348_), .C2(new_n349_), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n332_), .B(new_n334_), .C1(new_n339_), .C2(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n269_), .A2(KEYINPUT29), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G78gat), .B(G106gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n355_));
  XOR2_X1   g154(.A(new_n354_), .B(new_n355_), .Z(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n269_), .A2(KEYINPUT29), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G228gat), .A2(G233gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT88), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n310_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT91), .ZN(new_n362_));
  OR2_X1    g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n358_), .A2(new_n307_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n364_), .A2(G228gat), .A3(G233gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n361_), .A2(new_n362_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n363_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G22gat), .B(G50gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n368_), .B(KEYINPUT87), .Z(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n367_), .A2(new_n369_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n357_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n367_), .A2(new_n369_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n374_), .A2(new_n370_), .A3(new_n356_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n351_), .A2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n288_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT27), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n380_), .A2(KEYINPUT99), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(KEYINPUT99), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n339_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n328_), .A2(new_n329_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n338_), .B(KEYINPUT27), .C1(new_n320_), .C2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n379_), .A2(new_n383_), .A3(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n246_), .B1(new_n378_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n383_), .A2(new_n385_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n288_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n373_), .A2(new_n375_), .A3(new_n389_), .A4(new_n246_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  OR2_X1    g190(.A1(new_n387_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT13), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n393_), .A2(KEYINPUT69), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT68), .ZN(new_n395_));
  XOR2_X1   g194(.A(KEYINPUT67), .B(KEYINPUT5), .Z(new_n396_));
  XNOR2_X1  g195(.A(G120gat), .B(G148gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G176gat), .B(G204gat), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n398_), .B(new_n399_), .Z(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G230gat), .A2(G233gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G57gat), .A2(G64gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(G57gat), .A2(G64gat), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT11), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(G71gat), .B(G78gat), .Z(new_n407_));
  INV_X1    g206(.A(G57gat), .ZN(new_n408_));
  INV_X1    g207(.A(G64gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT11), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(new_n411_), .A3(new_n403_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n406_), .A2(new_n407_), .A3(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G71gat), .B(G78gat), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n414_), .B(KEYINPUT11), .C1(new_n405_), .C2(new_n404_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  XOR2_X1   g215(.A(KEYINPUT10), .B(G99gat), .Z(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT64), .B(G106gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT9), .ZN(new_n420_));
  INV_X1    g219(.A(G92gat), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n420_), .B1(new_n281_), .B2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT65), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n281_), .A2(new_n421_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT65), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n426_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n422_), .A2(new_n424_), .A3(new_n425_), .A4(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G99gat), .A2(G106gat), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT6), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n419_), .A2(new_n428_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT7), .ZN(new_n435_));
  INV_X1    g234(.A(G99gat), .ZN(new_n436_));
  INV_X1    g235(.A(G106gat), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n435_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n438_), .A2(new_n431_), .A3(new_n432_), .A4(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT8), .ZN(new_n441_));
  XOR2_X1   g240(.A(G85gat), .B(G92gat), .Z(new_n442_));
  AND3_X1   g241(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n441_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n416_), .B(new_n434_), .C1(new_n443_), .C2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT66), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n434_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n416_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n446_), .B1(new_n447_), .B2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n440_), .A2(new_n442_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT8), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n416_), .B1(new_n455_), .B2(new_n434_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT66), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n402_), .B1(new_n451_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n402_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n450_), .A2(KEYINPUT12), .A3(new_n445_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT12), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n448_), .A2(new_n461_), .A3(new_n449_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n459_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n401_), .B1(new_n458_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NOR3_X1   g264(.A1(new_n458_), .A2(new_n463_), .A3(new_n401_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n395_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n466_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(KEYINPUT68), .A3(new_n464_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n394_), .B1(new_n467_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n393_), .A2(KEYINPUT69), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n467_), .A2(new_n469_), .A3(KEYINPUT69), .A4(new_n393_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(G29gat), .B(G36gat), .Z(new_n475_));
  XNOR2_X1  g274(.A(G43gat), .B(G50gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(G43gat), .B(G50gat), .Z(new_n478_));
  XNOR2_X1  g277(.A(G29gat), .B(G36gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT15), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G15gat), .B(G22gat), .ZN(new_n484_));
  INV_X1    g283(.A(G1gat), .ZN(new_n485_));
  INV_X1    g284(.A(G8gat), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT14), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n484_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G1gat), .B(G8gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n483_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT75), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G229gat), .A2(G233gat), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n490_), .A2(new_n481_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n495_), .B1(new_n483_), .B2(new_n490_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n493_), .B(new_n494_), .C1(new_n492_), .C2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n490_), .B(new_n481_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(G229gat), .A3(G233gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G169gat), .B(G197gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT76), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G113gat), .B(G141gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n500_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n497_), .A2(new_n499_), .A3(new_n504_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n474_), .A2(new_n509_), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n392_), .A2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n449_), .B(new_n490_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G231gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G127gat), .B(G155gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(G211gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(KEYINPUT16), .B(G183gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(KEYINPUT73), .B(KEYINPUT17), .Z(new_n519_));
  AND2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n514_), .A2(KEYINPUT74), .A3(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(KEYINPUT74), .B1(new_n514_), .B2(new_n520_), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n518_), .B(KEYINPUT17), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n514_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n483_), .A2(new_n448_), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n448_), .A2(new_n481_), .ZN(new_n529_));
  XOR2_X1   g328(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n530_));
  NAND2_X1  g329(.A1(G232gat), .A2(G233gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT35), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n528_), .A2(new_n529_), .A3(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n532_), .A2(new_n533_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT36), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G190gat), .B(G218gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G134gat), .B(G162gat), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n539_), .B(new_n540_), .Z(new_n541_));
  NAND2_X1  g340(.A1(new_n535_), .A2(new_n536_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n537_), .A2(new_n538_), .A3(new_n541_), .A4(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(KEYINPUT71), .B(KEYINPUT37), .Z(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n536_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n535_), .B(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n541_), .B(KEYINPUT36), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n543_), .B(new_n545_), .C1(new_n547_), .C2(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n543_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n550_), .A2(KEYINPUT72), .B1(new_n551_), .B2(KEYINPUT37), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n547_), .A2(new_n549_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT72), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n553_), .A2(new_n543_), .A3(new_n554_), .A4(new_n545_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n527_), .B1(new_n552_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n511_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n288_), .A2(new_n485_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT38), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n551_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n527_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n511_), .A2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(G1gat), .B1(new_n564_), .B2(new_n389_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n565_), .A2(KEYINPUT100), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(KEYINPUT100), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n561_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT101), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT101), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n561_), .A2(new_n570_), .A3(new_n566_), .A4(new_n567_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(G1324gat));
  NAND4_X1  g371(.A1(new_n511_), .A2(new_n486_), .A3(new_n388_), .A4(new_n556_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n388_), .ZN(new_n574_));
  OAI21_X1  g373(.A(G8gat), .B1(new_n564_), .B2(new_n574_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n575_), .A2(KEYINPUT39), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(KEYINPUT39), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n573_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n578_), .B(new_n580_), .ZN(G1325gat));
  INV_X1    g380(.A(new_n246_), .ZN(new_n582_));
  OAI21_X1  g381(.A(G15gat), .B1(new_n564_), .B2(new_n582_), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n583_), .A2(KEYINPUT41), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(KEYINPUT41), .ZN(new_n585_));
  OR3_X1    g384(.A1(new_n557_), .A2(G15gat), .A3(new_n582_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n584_), .A2(new_n585_), .A3(new_n586_), .ZN(G1326gat));
  OAI21_X1  g386(.A(G22gat), .B1(new_n564_), .B2(new_n377_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT42), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n377_), .A2(G22gat), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n589_), .B1(new_n557_), .B2(new_n590_), .ZN(G1327gat));
  INV_X1    g390(.A(G29gat), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n550_), .A2(KEYINPUT72), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n551_), .A2(KEYINPUT37), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n593_), .A2(new_n555_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n596_), .B1(new_n387_), .B2(new_n391_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT43), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n598_), .B1(new_n596_), .B2(KEYINPUT103), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n597_), .A2(new_n600_), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n596_), .B(new_n599_), .C1(new_n387_), .C2(new_n391_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n601_), .A2(new_n510_), .A3(new_n527_), .A4(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT44), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n527_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n606_), .B1(new_n597_), .B2(new_n600_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n607_), .A2(KEYINPUT44), .A3(new_n510_), .A4(new_n602_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n605_), .A2(new_n288_), .A3(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT104), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n592_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n611_), .B1(new_n610_), .B2(new_n609_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n606_), .A2(new_n551_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n511_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n288_), .A2(new_n592_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n612_), .B1(new_n614_), .B2(new_n615_), .ZN(G1328gat));
  NAND3_X1  g415(.A1(new_n605_), .A2(new_n388_), .A3(new_n608_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT105), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n605_), .A2(KEYINPUT105), .A3(new_n388_), .A4(new_n608_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(G36gat), .A3(new_n620_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n574_), .A2(G36gat), .ZN(new_n622_));
  OR3_X1    g421(.A1(new_n614_), .A2(KEYINPUT45), .A3(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(KEYINPUT45), .B1(new_n614_), .B2(new_n622_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n621_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT46), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n621_), .A2(KEYINPUT46), .A3(new_n625_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1329gat));
  NAND4_X1  g429(.A1(new_n605_), .A2(G43gat), .A3(new_n246_), .A4(new_n608_), .ZN(new_n631_));
  XOR2_X1   g430(.A(KEYINPUT106), .B(G43gat), .Z(new_n632_));
  OAI21_X1  g431(.A(new_n632_), .B1(new_n614_), .B2(new_n582_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g434(.A1(new_n605_), .A2(new_n376_), .A3(new_n608_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(G50gat), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n377_), .A2(G50gat), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n637_), .B1(new_n614_), .B2(new_n638_), .ZN(G1331gat));
  INV_X1    g438(.A(new_n474_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n640_), .A2(new_n508_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n392_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(new_n563_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n643_), .A2(new_n408_), .A3(new_n389_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n556_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(new_n288_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n644_), .B1(new_n408_), .B2(new_n647_), .ZN(G1332gat));
  OAI21_X1  g447(.A(G64gat), .B1(new_n643_), .B2(new_n574_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT48), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n646_), .A2(new_n409_), .A3(new_n388_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1333gat));
  OAI21_X1  g451(.A(G71gat), .B1(new_n643_), .B2(new_n582_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT49), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n582_), .A2(G71gat), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n654_), .B1(new_n645_), .B2(new_n655_), .ZN(G1334gat));
  OAI21_X1  g455(.A(G78gat), .B1(new_n643_), .B2(new_n377_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT50), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n377_), .A2(G78gat), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n659_), .B(KEYINPUT107), .Z(new_n660_));
  OAI21_X1  g459(.A(new_n658_), .B1(new_n645_), .B2(new_n660_), .ZN(G1335gat));
  NAND3_X1  g460(.A1(new_n607_), .A2(new_n602_), .A3(new_n641_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n662_), .A2(new_n281_), .A3(new_n389_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n642_), .A2(new_n613_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(new_n288_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n663_), .B1(new_n666_), .B2(new_n281_), .ZN(G1336gat));
  NOR3_X1   g466(.A1(new_n662_), .A2(new_n421_), .A3(new_n574_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n665_), .A2(new_n388_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n669_), .B2(new_n421_), .ZN(G1337gat));
  OAI21_X1  g469(.A(G99gat), .B1(new_n662_), .B2(new_n582_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n246_), .A2(new_n417_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(new_n664_), .B2(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g473(.A(KEYINPUT52), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n607_), .A2(new_n376_), .A3(new_n602_), .A4(new_n641_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT108), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n676_), .A2(new_n677_), .A3(G106gat), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n677_), .B1(new_n676_), .B2(G106gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n675_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n680_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n682_), .A2(KEYINPUT52), .A3(new_n678_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n665_), .A2(new_n418_), .A3(new_n376_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n681_), .A2(new_n683_), .A3(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT53), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT53), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n681_), .A2(new_n683_), .A3(new_n687_), .A4(new_n684_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(G1339gat));
  NOR3_X1   g488(.A1(new_n388_), .A2(new_n376_), .A3(new_n582_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT58), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n460_), .A2(new_n459_), .A3(new_n462_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(KEYINPUT111), .B(KEYINPUT55), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(new_n463_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT55), .ZN(new_n695_));
  AOI211_X1 g494(.A(new_n695_), .B(new_n459_), .C1(new_n460_), .C2(new_n462_), .ZN(new_n696_));
  OAI21_X1  g495(.A(KEYINPUT112), .B1(new_n694_), .B2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n445_), .A2(KEYINPUT12), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n698_), .A2(new_n456_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n462_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n402_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n693_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT112), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n463_), .A2(KEYINPUT55), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n703_), .A2(new_n704_), .A3(new_n705_), .A4(new_n692_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n697_), .A2(new_n706_), .A3(new_n401_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT56), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n697_), .A2(new_n706_), .A3(KEYINPUT56), .A4(new_n401_), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n709_), .A2(KEYINPUT113), .A3(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n504_), .B1(new_n498_), .B2(new_n494_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n493_), .B1(new_n492_), .B2(new_n496_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(new_n494_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n507_), .A2(new_n714_), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n468_), .B(new_n715_), .C1(new_n710_), .C2(KEYINPUT113), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n691_), .B1(new_n711_), .B2(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n717_), .A2(KEYINPUT114), .A3(new_n596_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT114), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n715_), .A2(new_n468_), .ZN(new_n720_));
  AND4_X1   g519(.A1(KEYINPUT56), .A2(new_n697_), .A3(new_n401_), .A4(new_n706_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT113), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n720_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n709_), .A2(KEYINPUT113), .A3(new_n710_), .ZN(new_n724_));
  AOI21_X1  g523(.A(KEYINPUT58), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n719_), .B1(new_n725_), .B2(new_n595_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n723_), .A2(new_n724_), .A3(KEYINPUT58), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n718_), .A2(new_n726_), .A3(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n508_), .A2(new_n468_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n729_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n467_), .A2(new_n469_), .A3(new_n715_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n551_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT57), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n606_), .B1(new_n728_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n556_), .A2(new_n509_), .A3(new_n473_), .A4(new_n472_), .ZN(new_n736_));
  XOR2_X1   g535(.A(KEYINPUT109), .B(KEYINPUT54), .Z(new_n737_));
  OAI21_X1  g536(.A(new_n735_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n595_), .A2(new_n509_), .A3(new_n606_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n737_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n640_), .A2(new_n739_), .A3(KEYINPUT110), .A4(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n736_), .A2(new_n737_), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n738_), .A2(new_n741_), .A3(new_n742_), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n288_), .B(new_n690_), .C1(new_n734_), .C2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT115), .ZN(new_n745_));
  AOI21_X1  g544(.A(G113gat), .B1(new_n745_), .B2(new_n508_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT116), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n728_), .A2(new_n733_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(new_n527_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n738_), .A2(new_n741_), .A3(new_n742_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n389_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT59), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n751_), .A2(KEYINPUT117), .A3(new_n752_), .A4(new_n690_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT117), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n754_), .B1(new_n744_), .B2(KEYINPUT59), .ZN(new_n755_));
  AOI22_X1  g554(.A1(new_n753_), .A2(new_n755_), .B1(KEYINPUT59), .B2(new_n744_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT118), .Z(new_n757_));
  AND2_X1   g556(.A1(new_n508_), .A2(G113gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n747_), .B1(new_n757_), .B2(new_n758_), .ZN(G1340gat));
  INV_X1    g558(.A(KEYINPUT119), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT115), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n744_), .B(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(G120gat), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n763_), .A2(KEYINPUT60), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n640_), .A2(KEYINPUT60), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(new_n763_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n760_), .B1(new_n762_), .B2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n745_), .A2(KEYINPUT119), .A3(new_n766_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n753_), .A2(new_n755_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT120), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n640_), .B1(new_n744_), .B2(KEYINPUT59), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n771_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(G120gat), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n772_), .B1(new_n771_), .B2(new_n773_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n770_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT121), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n770_), .B(KEYINPUT121), .C1(new_n775_), .C2(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(G1341gat));
  AOI21_X1  g580(.A(G127gat), .B1(new_n745_), .B2(new_n606_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n527_), .A2(KEYINPUT122), .ZN(new_n783_));
  MUX2_X1   g582(.A(KEYINPUT122), .B(new_n783_), .S(G127gat), .Z(new_n784_));
  AOI21_X1  g583(.A(new_n782_), .B1(new_n757_), .B2(new_n784_), .ZN(G1342gat));
  AOI21_X1  g584(.A(G134gat), .B1(new_n745_), .B2(new_n562_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n596_), .A2(G134gat), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n757_), .B2(new_n787_), .ZN(G1343gat));
  NAND4_X1  g587(.A1(new_n751_), .A2(new_n376_), .A3(new_n574_), .A4(new_n582_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n789_), .A2(new_n509_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(new_n251_), .ZN(G1344gat));
  NOR2_X1   g590(.A1(new_n789_), .A2(new_n640_), .ZN(new_n792_));
  XOR2_X1   g591(.A(KEYINPUT123), .B(G148gat), .Z(new_n793_));
  XNOR2_X1  g592(.A(new_n792_), .B(new_n793_), .ZN(G1345gat));
  NOR2_X1   g593(.A1(new_n789_), .A2(new_n527_), .ZN(new_n795_));
  XOR2_X1   g594(.A(KEYINPUT61), .B(G155gat), .Z(new_n796_));
  XNOR2_X1  g595(.A(new_n795_), .B(new_n796_), .ZN(G1346gat));
  INV_X1    g596(.A(new_n789_), .ZN(new_n798_));
  AOI21_X1  g597(.A(G162gat), .B1(new_n798_), .B2(new_n562_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n595_), .A2(new_n250_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(KEYINPUT124), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n799_), .B1(new_n798_), .B2(new_n801_), .ZN(G1347gat));
  AOI21_X1  g601(.A(new_n574_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n390_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(G169gat), .B1(new_n805_), .B2(new_n509_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(KEYINPUT62), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n509_), .A2(new_n290_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT125), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n807_), .B1(new_n805_), .B2(new_n809_), .ZN(G1348gat));
  NOR2_X1   g609(.A1(new_n805_), .A2(new_n640_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(new_n221_), .ZN(G1349gat));
  NOR2_X1   g611(.A1(new_n805_), .A2(new_n527_), .ZN(new_n813_));
  MUX2_X1   g612(.A(G183gat), .B(new_n227_), .S(new_n813_), .Z(G1350gat));
  OAI21_X1  g613(.A(G190gat), .B1(new_n805_), .B2(new_n595_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n562_), .A2(new_n292_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n815_), .B1(new_n805_), .B2(new_n816_), .ZN(G1351gat));
  NAND2_X1  g616(.A1(new_n379_), .A2(new_n582_), .ZN(new_n818_));
  XOR2_X1   g617(.A(new_n818_), .B(KEYINPUT126), .Z(new_n819_));
  NAND2_X1  g618(.A1(new_n803_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n508_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n474_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g624(.A1(new_n821_), .A2(new_n606_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n827_));
  AND2_X1   g626(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n826_), .A2(new_n827_), .A3(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n829_), .B1(new_n826_), .B2(new_n827_), .ZN(G1354gat));
  XOR2_X1   g629(.A(KEYINPUT127), .B(G218gat), .Z(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n820_), .A2(new_n595_), .A3(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n821_), .A2(new_n562_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n834_), .B2(new_n832_), .ZN(G1355gat));
endmodule


