//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n607_, new_n608_, new_n609_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n823_, new_n824_, new_n825_, new_n826_, new_n828_,
    new_n829_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n875_, new_n876_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_;
  INV_X1    g000(.A(KEYINPUT66), .ZN(new_n202_));
  OR3_X1    g001(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT65), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n207_), .B1(G99gat), .B2(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n209_), .A2(KEYINPUT6), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n206_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(KEYINPUT6), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n207_), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n212_), .A2(new_n213_), .A3(KEYINPUT65), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n205_), .B1(new_n211_), .B2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G85gat), .B(G92gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n216_), .A2(KEYINPUT8), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n202_), .B1(new_n215_), .B2(new_n218_), .ZN(new_n219_));
  AND3_X1   g018(.A1(new_n212_), .A2(new_n213_), .A3(KEYINPUT65), .ZN(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT65), .B1(new_n212_), .B2(new_n213_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  OAI211_X1 g021(.A(KEYINPUT66), .B(new_n217_), .C1(new_n222_), .C2(new_n205_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n216_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n208_), .A2(new_n210_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n224_), .B1(new_n225_), .B2(new_n205_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT8), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n219_), .A2(new_n223_), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(G85gat), .ZN(new_n229_));
  INV_X1    g028(.A(G92gat), .ZN(new_n230_));
  NOR3_X1   g029(.A1(new_n229_), .A2(new_n230_), .A3(KEYINPUT9), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n231_), .B1(new_n224_), .B2(KEYINPUT9), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT10), .B(G99gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT64), .ZN(new_n234_));
  OAI221_X1 g033(.A(new_n232_), .B1(new_n220_), .B2(new_n221_), .C1(new_n234_), .C2(G106gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n228_), .A2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G29gat), .B(G36gat), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n237_), .A2(KEYINPUT71), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(KEYINPUT71), .ZN(new_n239_));
  XOR2_X1   g038(.A(G43gat), .B(G50gat), .Z(new_n240_));
  OR3_X1    g039(.A1(new_n238_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n240_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n242_));
  AND2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n236_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G232gat), .A2(G233gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT34), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n246_), .A2(KEYINPUT35), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n244_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n236_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n241_), .A2(new_n242_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT15), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n241_), .A2(new_n242_), .A3(KEYINPUT15), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n228_), .A2(KEYINPUT67), .A3(new_n235_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n250_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n248_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(KEYINPUT35), .A3(new_n246_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n246_), .A2(KEYINPUT35), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n248_), .A2(new_n257_), .A3(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(KEYINPUT72), .B(KEYINPUT36), .Z(new_n262_));
  NAND3_X1  g061(.A1(new_n259_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G190gat), .B(G218gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G134gat), .B(G162gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n259_), .A2(new_n261_), .ZN(new_n267_));
  XOR2_X1   g066(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n268_));
  AOI21_X1  g067(.A(new_n266_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n266_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n268_), .ZN(new_n271_));
  AOI211_X1 g070(.A(new_n270_), .B(new_n271_), .C1(new_n259_), .C2(new_n261_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n263_), .B1(new_n269_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT37), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT37), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n263_), .B(new_n275_), .C1(new_n269_), .C2(new_n272_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G127gat), .B(G155gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT16), .ZN(new_n279_));
  XOR2_X1   g078(.A(G183gat), .B(G211gat), .Z(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G57gat), .B(G64gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT11), .ZN(new_n283_));
  XOR2_X1   g082(.A(G71gat), .B(G78gat), .Z(new_n284_));
  OR2_X1    g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n282_), .A2(KEYINPUT11), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n283_), .A2(new_n284_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n285_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G231gat), .A2(G233gat), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n288_), .B(new_n289_), .Z(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT74), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G15gat), .B(G22gat), .ZN(new_n292_));
  INV_X1    g091(.A(G1gat), .ZN(new_n293_));
  INV_X1    g092(.A(G8gat), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT14), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n292_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G1gat), .B(G8gat), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n296_), .B(new_n297_), .Z(new_n298_));
  XNOR2_X1  g097(.A(new_n291_), .B(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT75), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n281_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT17), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT17), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n303_), .B1(new_n299_), .B2(new_n281_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n302_), .B1(new_n301_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n277_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT76), .ZN(new_n308_));
  INV_X1    g107(.A(new_n298_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n243_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n251_), .A2(new_n298_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G229gat), .A2(G233gat), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n253_), .A2(new_n254_), .A3(new_n309_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n311_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n315_), .B1(new_n317_), .B2(new_n314_), .ZN(new_n318_));
  XOR2_X1   g117(.A(G113gat), .B(G141gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT77), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G169gat), .B(G197gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n318_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n322_), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n315_), .B(new_n324_), .C1(new_n317_), .C2(new_n314_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n326_), .B(KEYINPUT78), .Z(new_n327_));
  INV_X1    g126(.A(KEYINPUT12), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n288_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n250_), .A2(new_n256_), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT68), .ZN(new_n332_));
  INV_X1    g131(.A(new_n236_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n328_), .B1(new_n333_), .B2(new_n288_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT68), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n250_), .A2(new_n335_), .A3(new_n256_), .A4(new_n330_), .ZN(new_n336_));
  AND2_X1   g135(.A1(G230gat), .A2(G233gat), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n337_), .B1(new_n333_), .B2(new_n288_), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n332_), .A2(new_n334_), .A3(new_n336_), .A4(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n333_), .A2(new_n288_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n333_), .A2(new_n288_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n337_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n339_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G176gat), .B(G204gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT70), .ZN(new_n346_));
  XOR2_X1   g145(.A(G120gat), .B(G148gat), .Z(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n344_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n344_), .A2(new_n350_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT13), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n351_), .A2(KEYINPUT13), .A3(new_n352_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(G204gat), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n358_), .A2(G197gat), .ZN(new_n359_));
  INV_X1    g158(.A(G197gat), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n360_), .A2(G204gat), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT21), .B1(new_n359_), .B2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G211gat), .B(G218gat), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT91), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n361_), .B1(new_n364_), .B2(new_n359_), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT91), .B1(new_n358_), .B2(G197gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n362_), .B(new_n363_), .C1(new_n367_), .C2(KEYINPUT21), .ZN(new_n368_));
  INV_X1    g167(.A(new_n363_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n367_), .A2(KEYINPUT21), .A3(new_n369_), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  OR2_X1    g170(.A1(KEYINPUT79), .A2(G183gat), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT80), .ZN(new_n373_));
  NAND2_X1  g172(.A1(KEYINPUT79), .A2(G183gat), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n372_), .B(KEYINPUT25), .C1(new_n373_), .C2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT25), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n376_), .A2(KEYINPUT80), .A3(G183gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT26), .B(G190gat), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n375_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT81), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT81), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n375_), .A2(new_n381_), .A3(new_n377_), .A4(new_n378_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G183gat), .A2(G190gat), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n384_), .A2(KEYINPUT23), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(KEYINPUT23), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(G169gat), .ZN(new_n390_));
  INV_X1    g189(.A(G176gat), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n389_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  OR3_X1    g191(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n383_), .A2(new_n387_), .A3(new_n394_), .ZN(new_n395_));
  OR2_X1    g194(.A1(new_n385_), .A2(KEYINPUT82), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n385_), .A2(KEYINPUT82), .A3(new_n386_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n372_), .A2(new_n374_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n396_), .B(new_n397_), .C1(G190gat), .C2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(G169gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n371_), .B1(new_n395_), .B2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G226gat), .A2(G233gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n387_), .B1(G183gat), .B2(G190gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n401_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT25), .B(G183gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n378_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n410_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n396_), .A2(new_n397_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n408_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n368_), .A2(new_n370_), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT20), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NOR3_X1   g214(.A1(new_n403_), .A2(new_n406_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n406_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n395_), .A2(new_n371_), .A3(new_n402_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT20), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n419_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n417_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n416_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G8gat), .B(G36gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT18), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G64gat), .B(G92gat), .ZN(new_n425_));
  XOR2_X1   g224(.A(new_n424_), .B(new_n425_), .Z(new_n426_));
  NAND2_X1  g225(.A1(new_n422_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n426_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n428_), .B1(new_n416_), .B2(new_n421_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT27), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n431_), .B1(new_n422_), .B2(new_n426_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n406_), .B1(new_n403_), .B2(new_n415_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n418_), .A2(new_n417_), .A3(new_n420_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n426_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT95), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  AOI211_X1 g237(.A(KEYINPUT95), .B(new_n426_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n433_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n432_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G155gat), .A2(G162gat), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT85), .ZN(new_n443_));
  OR3_X1    g242(.A1(new_n442_), .A2(new_n443_), .A3(KEYINPUT1), .ZN(new_n444_));
  OR2_X1    g243(.A1(G155gat), .A2(G162gat), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n443_), .B1(new_n442_), .B2(KEYINPUT1), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n442_), .A2(KEYINPUT1), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n444_), .A2(new_n445_), .A3(new_n446_), .A4(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(G141gat), .ZN(new_n449_));
  INV_X1    g248(.A(G148gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G141gat), .A2(G148gat), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n448_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(KEYINPUT2), .ZN(new_n454_));
  AND2_X1   g253(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n455_));
  NOR2_X1   g254(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n449_), .B(new_n450_), .C1(new_n455_), .C2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT87), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n451_), .A2(KEYINPUT87), .A3(KEYINPUT3), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n454_), .A2(new_n457_), .A3(new_n460_), .A4(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT88), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n445_), .A2(new_n442_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n463_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n453_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT89), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  OAI211_X1 g269(.A(KEYINPUT89), .B(new_n453_), .C1(new_n466_), .C2(new_n467_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G127gat), .B(G134gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G113gat), .B(G120gat), .ZN(new_n473_));
  XOR2_X1   g272(.A(new_n472_), .B(new_n473_), .Z(new_n474_));
  NAND3_X1  g273(.A1(new_n470_), .A2(new_n471_), .A3(new_n474_), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n468_), .A2(new_n474_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G225gat), .A2(G233gat), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G1gat), .B(G29gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(G85gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT0), .B(G57gat), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n480_), .B(new_n481_), .Z(new_n482_));
  AND3_X1   g281(.A1(new_n475_), .A2(KEYINPUT4), .A3(new_n476_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n477_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n484_), .B1(new_n475_), .B2(KEYINPUT4), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n478_), .B(new_n482_), .C1(new_n483_), .C2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT94), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n475_), .A2(KEYINPUT4), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n475_), .A2(KEYINPUT4), .A3(new_n476_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(new_n484_), .A3(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n482_), .B1(new_n490_), .B2(new_n478_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n487_), .A2(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n478_), .B1(new_n483_), .B2(new_n485_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n482_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n495_), .A2(KEYINPUT94), .A3(new_n486_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n441_), .B1(new_n492_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT84), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G71gat), .B(G99gat), .ZN(new_n499_));
  INV_X1    g298(.A(G43gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n394_), .A2(new_n387_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n502_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n399_), .A2(new_n401_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n501_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G227gat), .A2(G233gat), .ZN(new_n506_));
  INV_X1    g305(.A(G15gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT30), .ZN(new_n509_));
  INV_X1    g308(.A(new_n501_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n395_), .A2(new_n510_), .A3(new_n402_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n505_), .A2(new_n509_), .A3(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n509_), .B1(new_n505_), .B2(new_n511_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n498_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n474_), .B(KEYINPUT31), .ZN(new_n516_));
  INV_X1    g315(.A(new_n509_), .ZN(new_n517_));
  NOR3_X1   g316(.A1(new_n503_), .A2(new_n504_), .A3(new_n501_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n510_), .B1(new_n395_), .B2(new_n402_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n517_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(KEYINPUT83), .B1(new_n520_), .B2(new_n512_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n515_), .B(new_n516_), .C1(new_n521_), .C2(new_n498_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n516_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n513_), .A2(new_n514_), .ZN(new_n524_));
  OAI211_X1 g323(.A(KEYINPUT84), .B(new_n523_), .C1(new_n524_), .C2(KEYINPUT83), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n522_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n470_), .A2(KEYINPUT29), .A3(new_n471_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G228gat), .A2(G233gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT90), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n371_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n453_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n467_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n531_), .B1(new_n532_), .B2(new_n465_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT29), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n414_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n528_), .ZN(new_n536_));
  AOI22_X1  g335(.A1(new_n527_), .A2(new_n530_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT28), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n470_), .A2(new_n471_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n538_), .B1(new_n539_), .B2(new_n534_), .ZN(new_n540_));
  AOI211_X1 g339(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n470_), .C2(new_n471_), .ZN(new_n541_));
  NOR3_X1   g340(.A1(new_n537_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n537_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G78gat), .B(G106gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G22gat), .B(G50gat), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n545_), .B(new_n546_), .Z(new_n547_));
  NAND3_X1  g346(.A1(new_n543_), .A2(new_n544_), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n547_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n544_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n549_), .B1(new_n550_), .B2(new_n542_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n526_), .A2(new_n548_), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n526_), .B1(new_n551_), .B2(new_n548_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n497_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n426_), .A2(KEYINPUT32), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n556_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n422_), .A2(new_n556_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(KEYINPUT93), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT93), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n422_), .A2(new_n560_), .A3(new_n556_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n557_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n492_), .A2(new_n496_), .A3(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n475_), .A2(new_n476_), .A3(new_n484_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n564_), .A2(new_n494_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n488_), .A2(new_n477_), .A3(new_n489_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n430_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT33), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n486_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n486_), .A2(new_n568_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n567_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n563_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n522_), .A2(new_n525_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n548_), .A2(new_n551_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  AOI211_X1 g375(.A(new_n327_), .B(new_n357_), .C1(new_n555_), .C2(new_n576_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n308_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n492_), .A2(new_n496_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n578_), .A2(new_n293_), .A3(new_n580_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n355_), .A2(new_n356_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(new_n326_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n436_), .B(new_n437_), .ZN(new_n584_));
  AOI22_X1  g383(.A1(new_n584_), .A2(new_n433_), .B1(new_n431_), .B2(new_n430_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n487_), .A2(new_n491_), .ZN(new_n586_));
  AOI211_X1 g385(.A(KEYINPUT94), .B(new_n482_), .C1(new_n490_), .C2(new_n478_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n585_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n551_), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n550_), .A2(new_n542_), .A3(new_n549_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n573_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n588_), .B1(new_n591_), .B2(new_n552_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n574_), .B1(new_n563_), .B2(new_n571_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NOR4_X1   g393(.A1(new_n583_), .A2(new_n594_), .A3(new_n273_), .A4(new_n306_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n595_), .A2(new_n580_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n581_), .B1(new_n293_), .B2(new_n596_), .ZN(new_n597_));
  MUX2_X1   g396(.A(new_n581_), .B(new_n597_), .S(KEYINPUT38), .Z(G1324gat));
  NAND3_X1  g397(.A1(new_n578_), .A2(new_n294_), .A3(new_n441_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n595_), .A2(new_n441_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(G8gat), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n601_), .A2(KEYINPUT39), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(KEYINPUT39), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n599_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT40), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(G1325gat));
  AOI21_X1  g405(.A(new_n507_), .B1(new_n595_), .B2(new_n526_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT41), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n578_), .A2(new_n507_), .A3(new_n526_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(G1326gat));
  INV_X1    g409(.A(G22gat), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n589_), .A2(new_n590_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n611_), .B1(new_n595_), .B2(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n614_), .B(KEYINPUT42), .Z(new_n615_));
  NAND3_X1  g414(.A1(new_n578_), .A2(new_n611_), .A3(new_n613_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(G1327gat));
  NOR2_X1   g416(.A1(KEYINPUT98), .A2(KEYINPUT44), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n583_), .A2(new_n305_), .A3(new_n618_), .ZN(new_n619_));
  AOI22_X1  g418(.A1(new_n555_), .A2(new_n576_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT43), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n620_), .A2(KEYINPUT96), .A3(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n277_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT96), .ZN(new_n624_));
  AOI21_X1  g423(.A(KEYINPUT43), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n619_), .B1(new_n622_), .B2(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(KEYINPUT98), .B1(KEYINPUT97), .B2(KEYINPUT44), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n621_), .B1(new_n620_), .B2(KEYINPUT96), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n623_), .A2(new_n624_), .A3(KEYINPUT43), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(new_n619_), .A3(new_n627_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n579_), .B1(new_n629_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(G29gat), .ZN(new_n635_));
  INV_X1    g434(.A(new_n273_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n305_), .A2(new_n636_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n577_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n580_), .A2(new_n635_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT99), .ZN(new_n641_));
  OAI22_X1  g440(.A1(new_n634_), .A2(new_n635_), .B1(new_n639_), .B2(new_n641_), .ZN(G1328gat));
  INV_X1    g441(.A(new_n633_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n627_), .B1(new_n632_), .B2(new_n619_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n441_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(G36gat), .ZN(new_n646_));
  INV_X1    g445(.A(G36gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n638_), .A2(new_n647_), .A3(new_n441_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT45), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT46), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n646_), .A2(new_n649_), .A3(KEYINPUT100), .A4(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(KEYINPUT100), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n650_), .A2(KEYINPUT100), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n629_), .A2(new_n633_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n647_), .B1(new_n654_), .B2(new_n441_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT45), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n648_), .B(new_n656_), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n652_), .B(new_n653_), .C1(new_n655_), .C2(new_n657_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n651_), .A2(new_n658_), .ZN(G1329gat));
  NAND3_X1  g458(.A1(new_n638_), .A2(new_n500_), .A3(new_n526_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n573_), .B1(new_n629_), .B2(new_n633_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n660_), .B1(new_n661_), .B2(new_n500_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT47), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(G1330gat));
  AOI21_X1  g463(.A(G50gat), .B1(new_n638_), .B2(new_n613_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n613_), .A2(G50gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n654_), .B2(new_n666_), .ZN(G1331gat));
  NOR3_X1   g466(.A1(new_n594_), .A2(new_n326_), .A3(new_n582_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n308_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(G57gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(new_n670_), .A3(new_n580_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n594_), .A2(new_n273_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n327_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n306_), .A2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n672_), .A2(new_n357_), .A3(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G57gat), .B1(new_n675_), .B2(new_n579_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n671_), .A2(new_n676_), .ZN(G1332gat));
  OAI21_X1  g476(.A(G64gat), .B1(new_n675_), .B2(new_n585_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT48), .ZN(new_n679_));
  INV_X1    g478(.A(G64gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n669_), .A2(new_n680_), .A3(new_n441_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(G1333gat));
  OAI21_X1  g481(.A(G71gat), .B1(new_n675_), .B2(new_n573_), .ZN(new_n683_));
  XOR2_X1   g482(.A(KEYINPUT101), .B(KEYINPUT49), .Z(new_n684_));
  XNOR2_X1  g483(.A(new_n683_), .B(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n573_), .A2(G71gat), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT102), .Z(new_n687_));
  NAND2_X1  g486(.A1(new_n669_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n685_), .A2(new_n688_), .ZN(G1334gat));
  OAI21_X1  g488(.A(G78gat), .B1(new_n675_), .B2(new_n612_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT50), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n612_), .A2(G78gat), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT103), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n669_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n691_), .A2(new_n694_), .ZN(G1335gat));
  AND2_X1   g494(.A1(new_n668_), .A2(new_n637_), .ZN(new_n696_));
  AOI21_X1  g495(.A(G85gat), .B1(new_n696_), .B2(new_n580_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n326_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n357_), .A2(new_n306_), .A3(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n357_), .A2(new_n306_), .A3(KEYINPUT104), .A4(new_n698_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n632_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n580_), .A2(G85gat), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT105), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n697_), .B1(new_n704_), .B2(new_n706_), .ZN(G1336gat));
  NAND3_X1  g506(.A1(new_n696_), .A2(new_n230_), .A3(new_n441_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n704_), .A2(new_n441_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(new_n709_), .B2(new_n230_), .ZN(G1337gat));
  INV_X1    g509(.A(new_n234_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n696_), .A2(new_n711_), .A3(new_n526_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n632_), .A2(new_n526_), .A3(new_n703_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n713_), .A2(KEYINPUT106), .A3(G99gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(KEYINPUT106), .B1(new_n713_), .B2(G99gat), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n712_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g516(.A(G106gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n696_), .A2(new_n718_), .A3(new_n613_), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n613_), .B(new_n703_), .C1(new_n622_), .C2(new_n625_), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT108), .B1(new_n720_), .B2(G106gat), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n720_), .A2(KEYINPUT108), .A3(G106gat), .ZN(new_n722_));
  XOR2_X1   g521(.A(KEYINPUT107), .B(KEYINPUT52), .Z(new_n723_));
  AOI21_X1  g522(.A(new_n721_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n723_), .ZN(new_n725_));
  AOI211_X1 g524(.A(KEYINPUT108), .B(new_n725_), .C1(new_n720_), .C2(G106gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n719_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT53), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT53), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n729_), .B(new_n719_), .C1(new_n724_), .C2(new_n726_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1339gat));
  AND2_X1   g530(.A1(new_n351_), .A2(new_n326_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n332_), .A2(new_n340_), .A3(new_n334_), .A4(new_n336_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(new_n337_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT55), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n339_), .A2(new_n735_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n336_), .A2(new_n334_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n737_), .A2(KEYINPUT55), .A3(new_n332_), .A4(new_n338_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n734_), .A2(new_n736_), .A3(new_n738_), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n739_), .A2(KEYINPUT56), .A3(new_n350_), .ZN(new_n740_));
  AOI21_X1  g539(.A(KEYINPUT56), .B1(new_n739_), .B2(new_n350_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n732_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n312_), .A2(new_n313_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(new_n322_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n316_), .B2(new_n311_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n746_), .A2(new_n313_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n316_), .A2(new_n745_), .A3(new_n311_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n325_), .ZN(new_n750_));
  OAI21_X1  g549(.A(KEYINPUT111), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n752_));
  INV_X1    g551(.A(new_n748_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n753_), .A2(new_n313_), .A3(new_n746_), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n752_), .B(new_n325_), .C1(new_n754_), .C2(new_n744_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n751_), .A2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n273_), .B1(new_n742_), .B2(new_n758_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(KEYINPUT112), .B(KEYINPUT57), .ZN(new_n760_));
  OAI21_X1  g559(.A(KEYINPUT113), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n762_));
  INV_X1    g561(.A(new_n760_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n739_), .A2(new_n350_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT56), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n739_), .A2(KEYINPUT56), .A3(new_n350_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n757_), .B1(new_n768_), .B2(new_n732_), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n762_), .B(new_n763_), .C1(new_n769_), .C2(new_n273_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n759_), .A2(KEYINPUT57), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n351_), .A2(new_n751_), .A3(new_n755_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n772_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(KEYINPUT114), .A2(KEYINPUT58), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n774_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n768_), .A2(new_n772_), .A3(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n775_), .A2(new_n277_), .A3(new_n777_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n761_), .A2(new_n770_), .A3(new_n771_), .A4(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n306_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n277_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n674_), .A2(new_n781_), .A3(new_n582_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(KEYINPUT109), .B(KEYINPUT54), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n674_), .A2(new_n781_), .A3(new_n582_), .A4(new_n783_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n780_), .A2(new_n787_), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n552_), .A2(new_n579_), .A3(new_n441_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(G113gat), .B1(new_n791_), .B2(new_n326_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n771_), .A2(new_n778_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n759_), .A2(new_n760_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n306_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n787_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT59), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n789_), .A2(new_n797_), .ZN(new_n798_));
  AOI22_X1  g597(.A1(new_n790_), .A2(KEYINPUT59), .B1(new_n796_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n673_), .A2(G113gat), .ZN(new_n800_));
  XOR2_X1   g599(.A(new_n800_), .B(KEYINPUT115), .Z(new_n801_));
  AOI21_X1  g600(.A(new_n792_), .B1(new_n799_), .B2(new_n801_), .ZN(G1340gat));
  NAND2_X1  g601(.A1(new_n796_), .A2(new_n798_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n357_), .B(new_n803_), .C1(new_n791_), .C2(new_n797_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(G120gat), .ZN(new_n805_));
  INV_X1    g604(.A(G120gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n806_), .B1(new_n582_), .B2(KEYINPUT60), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n791_), .B(new_n807_), .C1(KEYINPUT60), .C2(new_n806_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n805_), .A2(new_n808_), .ZN(G1341gat));
  AOI21_X1  g608(.A(G127gat), .B1(new_n791_), .B2(new_n305_), .ZN(new_n810_));
  INV_X1    g609(.A(G127gat), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n305_), .B2(KEYINPUT116), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(KEYINPUT116), .B2(new_n811_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n810_), .B1(new_n799_), .B2(new_n813_), .ZN(G1342gat));
  INV_X1    g613(.A(G134gat), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n790_), .B2(new_n636_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT117), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT117), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n818_), .B(new_n815_), .C1(new_n790_), .C2(new_n636_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n277_), .A2(G134gat), .ZN(new_n820_));
  XOR2_X1   g619(.A(new_n820_), .B(KEYINPUT118), .Z(new_n821_));
  AOI22_X1  g620(.A1(new_n817_), .A2(new_n819_), .B1(new_n799_), .B2(new_n821_), .ZN(G1343gat));
  AOI22_X1  g621(.A1(new_n779_), .A2(new_n306_), .B1(new_n786_), .B2(new_n785_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n823_), .A2(new_n591_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n579_), .A2(new_n441_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n824_), .A2(new_n326_), .A3(new_n825_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g626(.A1(new_n824_), .A2(new_n357_), .A3(new_n825_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(KEYINPUT119), .B(G148gat), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n828_), .B(new_n829_), .ZN(G1345gat));
  NAND4_X1  g629(.A1(new_n788_), .A2(new_n554_), .A3(new_n305_), .A4(new_n825_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT120), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT120), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n824_), .A2(new_n833_), .A3(new_n305_), .A4(new_n825_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(KEYINPUT61), .B(G155gat), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n832_), .A2(new_n834_), .A3(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n832_), .B2(new_n834_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(G1346gat));
  NAND2_X1  g637(.A1(new_n824_), .A2(new_n825_), .ZN(new_n839_));
  OAI21_X1  g638(.A(G162gat), .B1(new_n839_), .B2(new_n781_), .ZN(new_n840_));
  OR2_X1    g639(.A1(new_n636_), .A2(G162gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n839_), .B2(new_n841_), .ZN(G1347gat));
  NOR2_X1   g641(.A1(new_n580_), .A2(new_n585_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n844_), .A2(new_n573_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT121), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n846_), .A2(new_n847_), .A3(new_n698_), .ZN(new_n848_));
  AOI21_X1  g647(.A(KEYINPUT121), .B1(new_n845_), .B2(new_n326_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n848_), .A2(new_n613_), .A3(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n390_), .B1(new_n796_), .B2(new_n850_), .ZN(new_n851_));
  AND2_X1   g650(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n613_), .B1(new_n795_), .B2(new_n787_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(KEYINPUT22), .B(G169gat), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n854_), .A2(new_n326_), .A3(new_n845_), .A4(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n853_), .A2(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n852_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n851_), .A2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT123), .B1(new_n857_), .B2(new_n861_), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n851_), .A2(new_n860_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT123), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n863_), .A2(new_n864_), .A3(new_n853_), .A4(new_n856_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n862_), .A2(new_n865_), .ZN(G1348gat));
  NOR4_X1   g665(.A1(new_n823_), .A2(new_n613_), .A3(new_n582_), .A4(new_n846_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n854_), .A2(new_n845_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n357_), .A2(new_n391_), .ZN(new_n869_));
  OAI22_X1  g668(.A1(new_n867_), .A2(new_n391_), .B1(new_n868_), .B2(new_n869_), .ZN(G1349gat));
  NAND4_X1  g669(.A1(new_n788_), .A2(new_n612_), .A3(new_n305_), .A4(new_n845_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n398_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n846_), .A2(new_n409_), .A3(new_n306_), .ZN(new_n873_));
  AOI22_X1  g672(.A1(new_n871_), .A2(new_n872_), .B1(new_n854_), .B2(new_n873_), .ZN(G1350gat));
  OAI21_X1  g673(.A(G190gat), .B1(new_n868_), .B2(new_n781_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n273_), .A2(new_n378_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n868_), .B2(new_n876_), .ZN(G1351gat));
  NAND3_X1  g676(.A1(new_n824_), .A2(new_n326_), .A3(new_n843_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(G197gat), .ZN(G1352gat));
  NOR4_X1   g678(.A1(new_n823_), .A2(new_n591_), .A3(new_n582_), .A4(new_n844_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n358_), .A2(KEYINPUT124), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n358_), .A2(KEYINPUT124), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n880_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n880_), .B2(new_n882_), .ZN(G1353gat));
  NAND3_X1  g683(.A1(new_n824_), .A2(new_n305_), .A3(new_n843_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT63), .B(G211gat), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n885_), .B2(new_n888_), .ZN(G1354gat));
  XOR2_X1   g688(.A(KEYINPUT125), .B(G218gat), .Z(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n277_), .A2(new_n891_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(KEYINPUT126), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n824_), .A2(new_n843_), .A3(new_n893_), .ZN(new_n894_));
  NOR4_X1   g693(.A1(new_n823_), .A2(new_n636_), .A3(new_n591_), .A4(new_n844_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(new_n891_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(KEYINPUT127), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT127), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n894_), .B(new_n898_), .C1(new_n895_), .C2(new_n891_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n899_), .ZN(G1355gat));
endmodule


