//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 0 1 0 1 1 1 1 0 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n765_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n919_, new_n921_, new_n922_, new_n924_, new_n925_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n948_, new_n949_, new_n950_, new_n952_, new_n953_, new_n954_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_,
    new_n989_, new_n990_, new_n991_;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  AOI21_X1  g003(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT86), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT3), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n202_), .B(new_n204_), .C1(new_n207_), .C2(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n203_), .B1(KEYINPUT1), .B2(new_n202_), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n202_), .A2(KEYINPUT1), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  AND2_X1   g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n218_), .A2(new_n208_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n214_), .A2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT28), .B1(new_n221_), .B2(KEYINPUT29), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT28), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT29), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n214_), .A2(new_n223_), .A3(new_n224_), .A4(new_n220_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G22gat), .B(G50gat), .ZN(new_n226_));
  AND3_X1   g025(.A1(new_n222_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n226_), .B1(new_n222_), .B2(new_n225_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  OR2_X1    g028(.A1(G197gat), .A2(G204gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G197gat), .A2(G204gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT21), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n230_), .A2(KEYINPUT21), .A3(new_n231_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G211gat), .B(G218gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n234_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT88), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n235_), .A2(new_n236_), .ZN(new_n239_));
  AND3_X1   g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n238_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n204_), .A2(new_n202_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n205_), .B(KEYINPUT86), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n243_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  AOI211_X1 g045(.A(new_n218_), .B(new_n208_), .C1(new_n215_), .C2(new_n216_), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT29), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n251_));
  OAI21_X1  g050(.A(G228gat), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n242_), .A2(new_n248_), .A3(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n237_), .A2(new_n239_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n248_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n252_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G78gat), .B(G106gat), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n253_), .A2(new_n257_), .A3(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n241_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n262_));
  AND4_X1   g061(.A1(new_n261_), .A2(new_n248_), .A3(new_n262_), .A4(new_n252_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n252_), .B1(new_n248_), .B2(new_n254_), .ZN(new_n264_));
  OAI211_X1 g063(.A(KEYINPUT89), .B(new_n258_), .C1(new_n263_), .C2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n229_), .A2(new_n260_), .A3(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n253_), .A2(new_n257_), .ZN(new_n267_));
  AOI21_X1  g066(.A(KEYINPUT89), .B1(new_n267_), .B2(new_n258_), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT90), .B1(new_n266_), .B2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n222_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n222_), .A2(new_n225_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n226_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  AND3_X1   g072(.A1(new_n260_), .A2(new_n270_), .A3(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n267_), .A2(new_n258_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT89), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT90), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n274_), .A2(new_n277_), .A3(new_n278_), .A4(new_n265_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n269_), .A2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n229_), .B1(new_n260_), .B2(new_n275_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT27), .ZN(new_n284_));
  INV_X1    g083(.A(G169gat), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT22), .B1(new_n285_), .B2(KEYINPUT84), .ZN(new_n286_));
  INV_X1    g085(.A(G176gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT22), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(G169gat), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n286_), .B(new_n287_), .C1(KEYINPUT84), .C2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT23), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n293_), .B(new_n294_), .C1(G183gat), .C2(G190gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT83), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n290_), .A2(new_n295_), .A3(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n285_), .A2(new_n287_), .A3(KEYINPUT82), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT82), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n301_), .B1(G169gat), .B2(G176gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT24), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT25), .B(G183gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT26), .B(G190gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n291_), .B(KEYINPUT23), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n305_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n296_), .B(KEYINPUT83), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n300_), .A2(new_n302_), .A3(KEYINPUT24), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n299_), .B1(new_n310_), .B2(new_n313_), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n261_), .A2(new_n314_), .A3(new_n262_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n312_), .B1(G169gat), .B2(G176gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n285_), .A2(KEYINPUT22), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n289_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT91), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n289_), .A2(new_n317_), .A3(KEYINPUT91), .ZN(new_n321_));
  AOI21_X1  g120(.A(G176gat), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n295_), .A2(new_n298_), .ZN(new_n323_));
  OAI22_X1  g122(.A1(new_n310_), .A2(new_n316_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT20), .B1(new_n324_), .B2(new_n254_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G226gat), .A2(G233gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT19), .ZN(new_n327_));
  NOR3_X1   g126(.A1(new_n315_), .A2(new_n325_), .A3(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n327_), .ZN(new_n329_));
  OR2_X1    g128(.A1(new_n310_), .A2(new_n313_), .ZN(new_n330_));
  OAI211_X1 g129(.A(new_n330_), .B(new_n299_), .C1(new_n240_), .C2(new_n241_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT20), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n332_), .B1(new_n324_), .B2(new_n254_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n329_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(G8gat), .B(G36gat), .Z(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT18), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G64gat), .B(G92gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NOR3_X1   g138(.A1(new_n328_), .A2(new_n334_), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n331_), .A2(new_n333_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(new_n327_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n325_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n242_), .A2(new_n314_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n343_), .A2(new_n329_), .A3(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n338_), .B1(new_n342_), .B2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n284_), .B1(new_n340_), .B2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n327_), .B1(new_n315_), .B2(new_n325_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n331_), .A2(new_n333_), .A3(new_n329_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n339_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n342_), .A2(new_n345_), .A3(new_n338_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(KEYINPUT27), .A3(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n347_), .A2(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n283_), .A2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G71gat), .B(G99gat), .ZN(new_n356_));
  INV_X1    g155(.A(G43gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT30), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G227gat), .A2(G233gat), .ZN(new_n360_));
  INV_X1    g159(.A(G15gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n359_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n359_), .A2(new_n362_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n314_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n365_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n314_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n367_), .A2(new_n363_), .A3(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT85), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n366_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT31), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G127gat), .B(G134gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G113gat), .B(G120gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT31), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n366_), .A2(new_n369_), .A3(new_n370_), .A4(new_n377_), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n372_), .A2(new_n376_), .A3(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n376_), .B1(new_n372_), .B2(new_n378_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G225gat), .A2(G233gat), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n376_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n214_), .A2(new_n220_), .A3(new_n375_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(new_n383_), .A3(KEYINPUT4), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT4), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n221_), .A2(new_n385_), .A3(new_n376_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n381_), .B1(new_n384_), .B2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G1gat), .B(G29gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT92), .B(KEYINPUT0), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G57gat), .B(G85gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n381_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n393_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n394_));
  OR3_X1    g193(.A1(new_n387_), .A2(new_n392_), .A3(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n392_), .B1(new_n387_), .B2(new_n394_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NOR3_X1   g196(.A1(new_n379_), .A2(new_n380_), .A3(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n355_), .A2(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n354_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n397_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n396_), .A2(KEYINPUT93), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT33), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n340_), .A2(new_n346_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT33), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n396_), .A2(KEYINPUT93), .A3(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n384_), .A2(new_n381_), .A3(new_n386_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n392_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n382_), .A2(new_n383_), .A3(new_n393_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n403_), .A2(new_n404_), .A3(new_n406_), .A4(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n338_), .A2(KEYINPUT32), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n412_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n328_), .A2(new_n334_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n413_), .B1(new_n414_), .B2(new_n412_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n397_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n411_), .A2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n281_), .B1(new_n269_), .B2(new_n279_), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n400_), .A2(new_n401_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n379_), .A2(new_n380_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n399_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT13), .ZN(new_n422_));
  AND2_X1   g221(.A1(G230gat), .A2(G233gat), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT10), .ZN(new_n424_));
  INV_X1    g223(.A(G99gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT64), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n426_), .A2(KEYINPUT64), .A3(new_n427_), .ZN(new_n431_));
  AOI21_X1  g230(.A(G106gat), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  OAI211_X1 g231(.A(G85gat), .B(G92gat), .C1(KEYINPUT65), .C2(KEYINPUT9), .ZN(new_n433_));
  OAI211_X1 g232(.A(KEYINPUT65), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(KEYINPUT65), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G99gat), .A2(G106gat), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT6), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n437_), .A2(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n432_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n438_), .ZN(new_n446_));
  AND2_X1   g245(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n447_));
  NOR2_X1   g246(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n446_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT66), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n439_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n451_), .A2(new_n438_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT7), .ZN(new_n454_));
  INV_X1    g253(.A(G106gat), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(new_n425_), .A3(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n449_), .A2(new_n453_), .A3(new_n456_), .A4(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(G85gat), .A2(G92gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G85gat), .A2(G92gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n458_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT8), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT8), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n456_), .A2(new_n457_), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n462_), .B(new_n465_), .C1(new_n466_), .C2(new_n442_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n445_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT67), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G57gat), .B(G64gat), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n469_), .B1(new_n470_), .B2(KEYINPUT11), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  OR2_X1    g271(.A1(new_n470_), .A2(KEYINPUT11), .ZN(new_n473_));
  XOR2_X1   g272(.A(G71gat), .B(G78gat), .Z(new_n474_));
  NAND3_X1  g273(.A1(new_n470_), .A2(new_n469_), .A3(KEYINPUT11), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .A4(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n474_), .B1(KEYINPUT11), .B2(new_n470_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n475_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n477_), .B1(new_n478_), .B2(new_n471_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n476_), .A2(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n423_), .B1(new_n468_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n431_), .ZN(new_n482_));
  AOI21_X1  g281(.A(KEYINPUT64), .B1(new_n426_), .B2(new_n427_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n455_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n442_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n465_), .B1(new_n458_), .B2(new_n462_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n466_), .A2(new_n442_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n459_), .A2(new_n465_), .A3(new_n460_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n486_), .B1(new_n487_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n476_), .A2(new_n479_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n438_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n496_), .A2(new_n466_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n461_), .B1(new_n497_), .B2(new_n453_), .ZN(new_n498_));
  OAI211_X1 g297(.A(KEYINPUT68), .B(new_n467_), .C1(new_n498_), .C2(new_n465_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT68), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n500_), .B1(new_n487_), .B2(new_n490_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n445_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n492_), .A2(KEYINPUT12), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n481_), .B(new_n495_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n468_), .A2(new_n480_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n493_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n423_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G120gat), .B(G148gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT5), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G176gat), .B(G204gat), .ZN(new_n510_));
  XOR2_X1   g309(.A(new_n509_), .B(new_n510_), .Z(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n504_), .A2(new_n507_), .A3(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n512_), .B1(new_n504_), .B2(new_n507_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n422_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n515_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(KEYINPUT13), .A3(new_n513_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G113gat), .B(G141gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G169gat), .B(G197gat), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n520_), .B(new_n521_), .Z(new_n522_));
  NAND2_X1  g321(.A1(G229gat), .A2(G233gat), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G1gat), .B(G8gat), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT76), .ZN(new_n527_));
  INV_X1    g326(.A(G8gat), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT74), .ZN(new_n529_));
  INV_X1    g328(.A(G1gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(KEYINPUT74), .A2(G1gat), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n528_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT14), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT75), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  AND2_X1   g334(.A1(KEYINPUT74), .A2(G1gat), .ZN(new_n536_));
  NOR2_X1   g335(.A1(KEYINPUT74), .A2(G1gat), .ZN(new_n537_));
  OAI21_X1  g336(.A(G8gat), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT75), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n538_), .A2(new_n539_), .A3(KEYINPUT14), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n535_), .A2(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(G15gat), .B(G22gat), .Z(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n527_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n544_));
  AOI211_X1 g343(.A(KEYINPUT76), .B(new_n542_), .C1(new_n535_), .C2(new_n540_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n526_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NOR3_X1   g345(.A1(new_n533_), .A2(KEYINPUT75), .A3(new_n534_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n539_), .B1(new_n538_), .B2(KEYINPUT14), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n543_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT76), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n541_), .A2(new_n527_), .A3(new_n543_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(new_n551_), .A3(new_n525_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G29gat), .B(G36gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G43gat), .B(G50gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n546_), .A2(new_n552_), .A3(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n556_), .B1(new_n546_), .B2(new_n552_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n524_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NOR3_X1   g358(.A1(new_n544_), .A2(new_n545_), .A3(new_n526_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n525_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n555_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT15), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n555_), .B(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n546_), .A2(new_n565_), .A3(new_n552_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n562_), .A2(new_n523_), .A3(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n522_), .B1(new_n559_), .B2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n559_), .A2(new_n567_), .A3(new_n522_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT81), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT81), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n559_), .A2(new_n567_), .A3(new_n571_), .A4(new_n522_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n568_), .B1(new_n570_), .B2(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n519_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n421_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G232gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT34), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT35), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n578_), .B(KEYINPUT70), .Z(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n499_), .A2(new_n501_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n564_), .B1(new_n581_), .B2(new_n486_), .ZN(new_n582_));
  OAI22_X1  g381(.A1(new_n491_), .A2(new_n556_), .B1(KEYINPUT35), .B2(new_n577_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n580_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n577_), .A2(KEYINPUT35), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(new_n468_), .B2(new_n555_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n586_), .B(new_n579_), .C1(new_n564_), .C2(new_n502_), .ZN(new_n587_));
  XOR2_X1   g386(.A(G134gat), .B(G162gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(G190gat), .B(G218gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT36), .ZN(new_n591_));
  AND3_X1   g390(.A1(new_n584_), .A2(new_n587_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT36), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n590_), .A2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT71), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n595_), .B1(new_n584_), .B2(new_n587_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n592_), .A2(new_n596_), .A3(KEYINPUT72), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n584_), .A2(new_n587_), .A3(new_n591_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT72), .ZN(new_n599_));
  OAI21_X1  g398(.A(KEYINPUT37), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(KEYINPUT73), .B1(new_n597_), .B2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n592_), .A2(new_n596_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT37), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n584_), .A2(new_n587_), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n599_), .B(new_n598_), .C1(new_n605_), .C2(new_n595_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n603_), .B1(new_n592_), .B2(KEYINPUT72), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT73), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n606_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n601_), .A2(new_n604_), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT80), .ZN(new_n612_));
  INV_X1    g411(.A(G231gat), .ZN(new_n613_));
  INV_X1    g412(.A(G233gat), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n616_), .B1(new_n546_), .B2(new_n552_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n546_), .A2(new_n552_), .A3(new_n616_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n618_), .A2(new_n480_), .A3(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n619_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n492_), .B1(new_n621_), .B2(new_n617_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT17), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G127gat), .B(G155gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G183gat), .B(G211gat), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n626_), .A2(new_n627_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n623_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n626_), .A2(new_n627_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(KEYINPUT17), .A3(new_n628_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT79), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n620_), .A2(new_n622_), .A3(new_n635_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n633_), .B(KEYINPUT78), .Z(new_n637_));
  AOI21_X1  g436(.A(new_n637_), .B1(new_n620_), .B2(new_n622_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n612_), .B1(new_n636_), .B2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n620_), .A2(new_n622_), .A3(new_n635_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n620_), .A2(new_n622_), .ZN(new_n641_));
  OAI211_X1 g440(.A(KEYINPUT80), .B(new_n640_), .C1(new_n641_), .C2(new_n637_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n639_), .A2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n611_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(KEYINPUT94), .B1(new_n575_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT94), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n644_), .A2(new_n421_), .A3(new_n647_), .A4(new_n574_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n397_), .B(KEYINPUT95), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n651_), .A2(new_n537_), .A3(new_n536_), .ZN(new_n652_));
  XOR2_X1   g451(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n653_));
  NAND3_X1  g452(.A1(new_n649_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n420_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n339_), .B1(new_n328_), .B2(new_n334_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n656_), .A2(new_n352_), .A3(new_n410_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n405_), .B1(new_n396_), .B2(KEYINPUT93), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  AOI22_X1  g458(.A1(new_n659_), .A2(new_n406_), .B1(new_n397_), .B2(new_n415_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n660_), .A2(new_n283_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n418_), .A2(new_n397_), .A3(new_n354_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n655_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n602_), .B1(new_n663_), .B2(new_n399_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n636_), .A2(new_n638_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n574_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT97), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT97), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n574_), .A2(new_n668_), .A3(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n664_), .A2(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(G1gat), .B1(new_n671_), .B2(new_n401_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n654_), .A2(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n653_), .B1(new_n649_), .B2(new_n652_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT98), .ZN(G1324gat));
  INV_X1    g475(.A(KEYINPUT101), .ZN(new_n677_));
  INV_X1    g476(.A(new_n602_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n670_), .A2(new_n678_), .A3(new_n421_), .A4(new_n354_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT99), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n664_), .A2(KEYINPUT99), .A3(new_n670_), .A4(new_n354_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(G8gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(KEYINPUT39), .B1(new_n682_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT39), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n681_), .A2(new_n686_), .A3(G8gat), .A4(new_n683_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n354_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n689_), .A2(G8gat), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n646_), .A2(new_n648_), .A3(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n677_), .B1(new_n688_), .B2(new_n692_), .ZN(new_n693_));
  AOI211_X1 g492(.A(KEYINPUT101), .B(new_n691_), .C1(new_n685_), .C2(new_n687_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n693_), .A2(new_n694_), .A3(new_n696_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n683_), .A2(G8gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n686_), .B1(new_n698_), .B2(new_n681_), .ZN(new_n699_));
  AND4_X1   g498(.A1(new_n686_), .A2(new_n681_), .A3(G8gat), .A4(new_n683_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n692_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT101), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n688_), .A2(new_n677_), .A3(new_n692_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n695_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n697_), .A2(new_n704_), .ZN(G1325gat));
  OAI21_X1  g504(.A(G15gat), .B1(new_n671_), .B2(new_n655_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(KEYINPUT102), .B(KEYINPUT41), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n707_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n575_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(new_n644_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n420_), .A2(new_n361_), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n708_), .B(new_n709_), .C1(new_n711_), .C2(new_n712_), .ZN(G1326gat));
  XNOR2_X1  g512(.A(new_n418_), .B(KEYINPUT103), .ZN(new_n714_));
  OAI21_X1  g513(.A(G22gat), .B1(new_n671_), .B2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT42), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n714_), .A2(G22gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n711_), .B2(new_n717_), .ZN(G1327gat));
  INV_X1    g517(.A(new_n643_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n719_), .A2(new_n678_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n421_), .A2(new_n574_), .A3(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n421_), .A2(KEYINPUT105), .A3(new_n574_), .A4(new_n720_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(G29gat), .B1(new_n726_), .B2(new_n397_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n421_), .A2(new_n611_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT43), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n421_), .A2(new_n731_), .A3(new_n611_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n574_), .A2(new_n643_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n728_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n733_), .A2(new_n734_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n736_), .B2(KEYINPUT44), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n650_), .A2(G29gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n727_), .B1(new_n737_), .B2(new_n738_), .ZN(G1328gat));
  INV_X1    g538(.A(KEYINPUT46), .ZN(new_n740_));
  INV_X1    g539(.A(G36gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n737_), .B2(new_n354_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n689_), .A2(G36gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n723_), .A2(new_n724_), .A3(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT106), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT106), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n723_), .A2(new_n747_), .A3(new_n724_), .A4(new_n743_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n745_), .A2(new_n746_), .A3(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n746_), .B1(new_n745_), .B2(new_n748_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n740_), .B1(new_n742_), .B2(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n733_), .A2(KEYINPUT44), .A3(new_n734_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n753_), .B1(new_n736_), .B2(new_n728_), .ZN(new_n754_));
  OAI21_X1  g553(.A(G36gat), .B1(new_n754_), .B2(new_n689_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n755_), .B(KEYINPUT46), .C1(new_n750_), .C2(new_n749_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n752_), .A2(new_n756_), .ZN(G1329gat));
  NAND3_X1  g556(.A1(new_n737_), .A2(G43gat), .A3(new_n420_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n357_), .B1(new_n725_), .B2(new_n655_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT47), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT47), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n758_), .A2(new_n762_), .A3(new_n759_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1330gat));
  INV_X1    g563(.A(new_n714_), .ZN(new_n765_));
  AOI21_X1  g564(.A(G50gat), .B1(new_n726_), .B2(new_n765_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n283_), .A2(G50gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n737_), .B2(new_n767_), .ZN(G1331gat));
  INV_X1    g567(.A(new_n519_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n573_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n421_), .A2(new_n771_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n772_), .A2(new_n644_), .ZN(new_n773_));
  INV_X1    g572(.A(G57gat), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n773_), .A2(new_n774_), .A3(new_n650_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n664_), .A2(new_n719_), .A3(new_n573_), .A4(new_n519_), .ZN(new_n776_));
  OAI21_X1  g575(.A(G57gat), .B1(new_n776_), .B2(new_n401_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(new_n778_));
  XOR2_X1   g577(.A(new_n778_), .B(KEYINPUT107), .Z(G1332gat));
  OAI21_X1  g578(.A(G64gat), .B1(new_n776_), .B2(new_n689_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT48), .ZN(new_n781_));
  INV_X1    g580(.A(G64gat), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n773_), .A2(new_n782_), .A3(new_n354_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(G1333gat));
  OAI21_X1  g583(.A(G71gat), .B1(new_n776_), .B2(new_n655_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT49), .ZN(new_n786_));
  INV_X1    g585(.A(G71gat), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n773_), .A2(new_n787_), .A3(new_n420_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(G1334gat));
  OAI21_X1  g588(.A(G78gat), .B1(new_n776_), .B2(new_n714_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT50), .ZN(new_n791_));
  INV_X1    g590(.A(G78gat), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n773_), .A2(new_n792_), .A3(new_n765_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(G1335gat));
  NAND2_X1  g593(.A1(new_n772_), .A2(new_n720_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(G85gat), .B1(new_n796_), .B2(new_n650_), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n733_), .A2(new_n643_), .A3(new_n771_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n397_), .A2(G85gat), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT108), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n797_), .B1(new_n798_), .B2(new_n800_), .ZN(G1336gat));
  INV_X1    g600(.A(G92gat), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n796_), .A2(new_n802_), .A3(new_n354_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n798_), .A2(new_n354_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n803_), .B1(new_n804_), .B2(new_n802_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT109), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n805_), .B(new_n806_), .ZN(G1337gat));
  OAI211_X1 g606(.A(new_n796_), .B(new_n420_), .C1(new_n482_), .C2(new_n483_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n733_), .A2(new_n643_), .A3(new_n420_), .A4(new_n771_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT110), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n809_), .A2(new_n810_), .A3(G99gat), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n810_), .B1(new_n809_), .B2(G99gat), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n808_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g613(.A1(new_n796_), .A2(new_n455_), .A3(new_n283_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n733_), .A2(new_n643_), .A3(new_n283_), .A4(new_n771_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n816_), .A2(new_n817_), .A3(G106gat), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n817_), .B1(new_n816_), .B2(G106gat), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n815_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n820_), .B(new_n822_), .ZN(G1339gat));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n523_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n522_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n562_), .A2(new_n524_), .A3(new_n566_), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n825_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n828_), .B1(new_n570_), .B2(new_n572_), .ZN(new_n829_));
  XOR2_X1   g628(.A(KEYINPUT113), .B(KEYINPUT55), .Z(new_n830_));
  NAND2_X1  g629(.A1(new_n504_), .A2(new_n830_), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n495_), .B(new_n505_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n423_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n581_), .A2(new_n486_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n503_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n836_), .A2(KEYINPUT55), .A3(new_n495_), .A4(new_n481_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n831_), .A2(new_n833_), .A3(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n838_), .A2(KEYINPUT56), .A3(new_n511_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT56), .B1(new_n838_), .B2(new_n511_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n829_), .B(new_n513_), .C1(new_n840_), .C2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT58), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n824_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  AOI211_X1 g643(.A(new_n514_), .B(new_n828_), .C1(new_n570_), .C2(new_n572_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n838_), .A2(new_n511_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT56), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n839_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n845_), .A2(new_n849_), .A3(KEYINPUT115), .A4(KEYINPUT58), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n842_), .A2(new_n843_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n844_), .A2(new_n611_), .A3(new_n850_), .A4(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT57), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT114), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n570_), .A2(new_n572_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n568_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n514_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n849_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n517_), .A2(new_n513_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n829_), .A2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n855_), .B1(new_n862_), .B2(new_n678_), .ZN(new_n863_));
  AOI22_X1  g662(.A1(new_n858_), .A2(new_n849_), .B1(new_n860_), .B2(new_n829_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n864_), .A2(new_n602_), .A3(new_n854_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n852_), .B1(new_n863_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n665_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n573_), .A2(new_n639_), .A3(new_n642_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT112), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n573_), .A2(new_n639_), .A3(new_n642_), .A4(KEYINPUT112), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n871_), .A2(new_n610_), .A3(new_n769_), .A4(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(KEYINPUT54), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n872_), .A2(new_n769_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n875_), .A2(new_n876_), .A3(new_n610_), .A4(new_n871_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n874_), .A2(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n868_), .A2(KEYINPUT116), .A3(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT116), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n862_), .A2(new_n678_), .A3(new_n855_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n854_), .B1(new_n864_), .B2(new_n602_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n665_), .B1(new_n883_), .B2(new_n852_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n874_), .A2(new_n877_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n880_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n355_), .A2(new_n420_), .A3(new_n650_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n879_), .A2(new_n886_), .A3(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(G113gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n890_), .A2(new_n891_), .A3(new_n770_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n719_), .B1(new_n883_), .B2(new_n852_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n893_), .A2(new_n885_), .ZN(new_n894_));
  XOR2_X1   g693(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n895_));
  NOR3_X1   g694(.A1(new_n894_), .A2(new_n887_), .A3(new_n895_), .ZN(new_n896_));
  AOI211_X1 g695(.A(new_n573_), .B(new_n896_), .C1(KEYINPUT59), .C2(new_n889_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n892_), .B1(new_n897_), .B2(new_n891_), .ZN(G1340gat));
  AOI211_X1 g697(.A(new_n769_), .B(new_n896_), .C1(KEYINPUT59), .C2(new_n889_), .ZN(new_n899_));
  INV_X1    g698(.A(G120gat), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n769_), .A2(KEYINPUT60), .ZN(new_n901_));
  MUX2_X1   g700(.A(KEYINPUT60), .B(new_n901_), .S(new_n900_), .Z(new_n902_));
  AND3_X1   g701(.A1(new_n890_), .A2(KEYINPUT118), .A3(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(KEYINPUT118), .B1(new_n890_), .B2(new_n902_), .ZN(new_n904_));
  OAI22_X1  g703(.A1(new_n899_), .A2(new_n900_), .B1(new_n903_), .B2(new_n904_), .ZN(G1341gat));
  INV_X1    g704(.A(G127gat), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n890_), .A2(new_n906_), .A3(new_n719_), .ZN(new_n907_));
  AOI211_X1 g706(.A(new_n867_), .B(new_n896_), .C1(KEYINPUT59), .C2(new_n889_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(new_n906_), .ZN(G1342gat));
  INV_X1    g708(.A(G134gat), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n890_), .A2(new_n910_), .A3(new_n602_), .ZN(new_n911_));
  AOI211_X1 g710(.A(new_n610_), .B(new_n896_), .C1(KEYINPUT59), .C2(new_n889_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n912_), .B2(new_n910_), .ZN(G1343gat));
  NAND2_X1  g712(.A1(new_n879_), .A2(new_n886_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n655_), .A2(new_n400_), .A3(new_n650_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n770_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g717(.A1(new_n916_), .A2(new_n519_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g719(.A1(new_n916_), .A2(new_n719_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(KEYINPUT61), .B(G155gat), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n921_), .B(new_n922_), .ZN(G1346gat));
  INV_X1    g722(.A(G162gat), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n916_), .A2(new_n924_), .A3(new_n602_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n914_), .A2(new_n610_), .A3(new_n915_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n925_), .B1(new_n924_), .B2(new_n926_), .ZN(G1347gat));
  NAND3_X1  g726(.A1(new_n651_), .A2(new_n354_), .A3(new_n420_), .ZN(new_n928_));
  OR3_X1    g727(.A1(new_n894_), .A2(new_n765_), .A3(new_n928_), .ZN(new_n929_));
  OAI21_X1  g728(.A(G169gat), .B1(new_n929_), .B2(new_n573_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(KEYINPUT119), .B(KEYINPUT62), .ZN(new_n931_));
  OR2_X1    g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  INV_X1    g731(.A(new_n929_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n320_), .A2(new_n321_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n933_), .A2(new_n934_), .A3(new_n770_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n930_), .A2(new_n931_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n932_), .A2(new_n935_), .A3(new_n936_), .ZN(G1348gat));
  AOI21_X1  g736(.A(KEYINPUT116), .B1(new_n868_), .B2(new_n878_), .ZN(new_n938_));
  NOR3_X1   g737(.A1(new_n884_), .A2(new_n885_), .A3(new_n880_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n928_), .A2(new_n283_), .ZN(new_n941_));
  NAND4_X1  g740(.A1(new_n940_), .A2(G176gat), .A3(new_n519_), .A4(new_n941_), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT120), .ZN(new_n943_));
  AND2_X1   g742(.A1(new_n942_), .A2(new_n943_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n942_), .A2(new_n943_), .ZN(new_n945_));
  AOI21_X1  g744(.A(G176gat), .B1(new_n933_), .B2(new_n519_), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n944_), .A2(new_n945_), .A3(new_n946_), .ZN(G1349gat));
  NAND3_X1  g746(.A1(new_n940_), .A2(new_n719_), .A3(new_n941_), .ZN(new_n948_));
  INV_X1    g747(.A(G183gat), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n867_), .A2(new_n306_), .ZN(new_n950_));
  AOI22_X1  g749(.A1(new_n948_), .A2(new_n949_), .B1(new_n933_), .B2(new_n950_), .ZN(G1350gat));
  OAI21_X1  g750(.A(G190gat), .B1(new_n929_), .B2(new_n610_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n602_), .A2(new_n307_), .ZN(new_n953_));
  XOR2_X1   g752(.A(new_n953_), .B(KEYINPUT121), .Z(new_n954_));
  OAI21_X1  g753(.A(new_n952_), .B1(new_n929_), .B2(new_n954_), .ZN(G1351gat));
  NOR3_X1   g754(.A1(new_n420_), .A2(new_n397_), .A3(new_n418_), .ZN(new_n956_));
  AND2_X1   g755(.A1(new_n956_), .A2(KEYINPUT122), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n956_), .A2(KEYINPUT122), .ZN(new_n958_));
  NOR3_X1   g757(.A1(new_n957_), .A2(new_n958_), .A3(new_n689_), .ZN(new_n959_));
  AND3_X1   g758(.A1(new_n879_), .A2(new_n886_), .A3(new_n959_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n960_), .A2(new_n770_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n961_), .B(G197gat), .ZN(G1352gat));
  NAND4_X1  g761(.A1(new_n879_), .A2(new_n886_), .A3(new_n519_), .A4(new_n959_), .ZN(new_n963_));
  OR3_X1    g762(.A1(new_n963_), .A2(KEYINPUT125), .A3(G204gat), .ZN(new_n964_));
  OAI21_X1  g763(.A(KEYINPUT125), .B1(new_n963_), .B2(G204gat), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n964_), .A2(new_n965_), .ZN(new_n966_));
  INV_X1    g765(.A(G204gat), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n967_), .B1(new_n963_), .B2(KEYINPUT123), .ZN(new_n968_));
  INV_X1    g767(.A(KEYINPUT123), .ZN(new_n969_));
  NAND4_X1  g768(.A1(new_n940_), .A2(new_n969_), .A3(new_n519_), .A4(new_n959_), .ZN(new_n970_));
  AND3_X1   g769(.A1(new_n968_), .A2(new_n970_), .A3(KEYINPUT124), .ZN(new_n971_));
  AOI21_X1  g770(.A(KEYINPUT124), .B1(new_n968_), .B2(new_n970_), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n966_), .B1(new_n971_), .B2(new_n972_), .ZN(G1353gat));
  AOI21_X1  g772(.A(new_n867_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n974_));
  NAND4_X1  g773(.A1(new_n879_), .A2(new_n886_), .A3(new_n959_), .A4(new_n974_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n975_), .A2(KEYINPUT126), .ZN(new_n976_));
  INV_X1    g775(.A(new_n976_), .ZN(new_n977_));
  NOR2_X1   g776(.A1(new_n975_), .A2(KEYINPUT126), .ZN(new_n978_));
  OAI22_X1  g777(.A1(new_n977_), .A2(new_n978_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n979_));
  INV_X1    g778(.A(new_n978_), .ZN(new_n980_));
  NOR2_X1   g779(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n981_));
  NAND3_X1  g780(.A1(new_n980_), .A2(new_n981_), .A3(new_n976_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n979_), .A2(new_n982_), .ZN(G1354gat));
  INV_X1    g782(.A(G218gat), .ZN(new_n984_));
  NAND3_X1  g783(.A1(new_n960_), .A2(new_n984_), .A3(new_n602_), .ZN(new_n985_));
  NAND4_X1  g784(.A1(new_n879_), .A2(new_n886_), .A3(new_n611_), .A4(new_n959_), .ZN(new_n986_));
  NAND2_X1  g785(.A1(new_n986_), .A2(G218gat), .ZN(new_n987_));
  NAND2_X1  g786(.A1(new_n985_), .A2(new_n987_), .ZN(new_n988_));
  NAND2_X1  g787(.A1(new_n988_), .A2(KEYINPUT127), .ZN(new_n989_));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n990_));
  NAND3_X1  g789(.A1(new_n985_), .A2(new_n990_), .A3(new_n987_), .ZN(new_n991_));
  NAND2_X1  g790(.A1(new_n989_), .A2(new_n991_), .ZN(G1355gat));
endmodule


