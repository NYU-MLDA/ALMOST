//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n874_, new_n875_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_;
  XNOR2_X1  g000(.A(KEYINPUT10), .B(G99gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  AND2_X1   g002(.A1(new_n203_), .A2(KEYINPUT6), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(KEYINPUT6), .ZN(new_n205_));
  OAI22_X1  g004(.A1(new_n202_), .A2(G106gat), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT9), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n208_), .A2(KEYINPUT64), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n209_), .B1(new_n208_), .B2(KEYINPUT64), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G85gat), .ZN(new_n214_));
  INV_X1    g013(.A(G92gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(KEYINPUT65), .B1(new_n213_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n208_), .A2(KEYINPUT64), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT9), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n219_), .A2(new_n216_), .A3(new_n210_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n207_), .B1(new_n217_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n226_));
  OR3_X1    g025(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n226_), .B(new_n227_), .C1(new_n204_), .C2(new_n205_), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n216_), .A2(new_n208_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT8), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT8), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n228_), .A2(new_n232_), .A3(new_n229_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n213_), .A2(KEYINPUT65), .A3(new_n216_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n220_), .A2(new_n221_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n206_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT66), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n225_), .A2(new_n234_), .A3(new_n238_), .ZN(new_n239_));
  XOR2_X1   g038(.A(G71gat), .B(G78gat), .Z(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G57gat), .B(G64gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT11), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n242_), .A2(KEYINPUT11), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n240_), .A2(KEYINPUT11), .A3(new_n242_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n244_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n239_), .A2(KEYINPUT12), .A3(new_n247_), .ZN(new_n248_));
  AND2_X1   g047(.A1(G230gat), .A2(G233gat), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n228_), .A2(new_n232_), .A3(new_n229_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n232_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n252_), .A2(new_n237_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n247_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n249_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n254_), .B1(new_n234_), .B2(new_n223_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n257_));
  NOR3_X1   g056(.A1(new_n256_), .A2(new_n257_), .A3(KEYINPUT12), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n247_), .B1(new_n252_), .B2(new_n237_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT12), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT67), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n248_), .B(new_n255_), .C1(new_n258_), .C2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n253_), .A2(new_n254_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(new_n259_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(new_n249_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G176gat), .B(G204gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G120gat), .B(G148gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n266_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n266_), .A2(new_n271_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT13), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n273_), .A2(KEYINPUT13), .A3(new_n274_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(G141gat), .A2(G148gat), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT3), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G141gat), .A2(G148gat), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT2), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n282_), .A2(new_n285_), .A3(new_n286_), .A4(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G155gat), .A2(G162gat), .ZN(new_n289_));
  AND2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT86), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n292_), .A2(KEYINPUT87), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT87), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n294_), .A2(KEYINPUT86), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n291_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(KEYINPUT86), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n292_), .A2(KEYINPUT87), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n297_), .B(new_n298_), .C1(G155gat), .C2(G162gat), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT1), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n289_), .B(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n296_), .A2(new_n302_), .A3(new_n299_), .ZN(new_n303_));
  XOR2_X1   g102(.A(G141gat), .B(G148gat), .Z(new_n304_));
  AOI22_X1  g103(.A1(new_n290_), .A2(new_n300_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT29), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT92), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT21), .ZN(new_n308_));
  INV_X1    g107(.A(G197gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n309_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT90), .ZN(new_n311_));
  INV_X1    g110(.A(G204gat), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n311_), .B1(G197gat), .B2(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n312_), .A2(G197gat), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n308_), .B(new_n310_), .C1(new_n313_), .C2(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(G211gat), .B(G218gat), .Z(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n309_), .A2(G204gat), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT21), .B1(new_n314_), .B2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n315_), .A2(new_n317_), .A3(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n310_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n321_), .A2(KEYINPUT21), .A3(new_n316_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n303_), .A2(new_n304_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n288_), .A2(new_n296_), .A3(new_n299_), .A4(new_n289_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT92), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n326_), .A2(new_n327_), .A3(KEYINPUT29), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n307_), .A2(new_n323_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT93), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G228gat), .A2(G233gat), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n329_), .A2(new_n330_), .A3(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n330_), .B1(new_n329_), .B2(new_n332_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT88), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n324_), .A2(new_n336_), .A3(new_n325_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n336_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT29), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n339_), .A2(new_n323_), .A3(new_n331_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT91), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n340_), .A2(new_n341_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n333_), .B(new_n335_), .C1(new_n342_), .C2(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(G78gat), .B(G106gat), .Z(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(KEYINPUT94), .B1(new_n344_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n305_), .A2(new_n336_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n326_), .A2(KEYINPUT88), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(new_n349_), .A3(new_n306_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G22gat), .B(G50gat), .Z(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n350_), .B(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n344_), .A2(new_n346_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n340_), .B(new_n341_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n333_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n358_), .A2(new_n334_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n345_), .B1(new_n357_), .B2(new_n359_), .ZN(new_n360_));
  OAI22_X1  g159(.A1(new_n347_), .A2(new_n355_), .B1(new_n356_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n360_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n357_), .A2(new_n359_), .A3(new_n345_), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n362_), .A2(new_n363_), .A3(KEYINPUT94), .A4(new_n354_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n361_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT103), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n367_), .B(KEYINPUT101), .Z(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT4), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT85), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G127gat), .B(G134gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G113gat), .B(G120gat), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n371_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n372_), .B(new_n373_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n374_), .B1(new_n375_), .B2(new_n371_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n376_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n305_), .A2(new_n375_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n370_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n348_), .A2(new_n349_), .ZN(new_n380_));
  AOI21_X1  g179(.A(KEYINPUT4), .B1(new_n380_), .B2(new_n376_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n369_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n377_), .A2(new_n378_), .A3(new_n367_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G1gat), .B(G29gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(G85gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT0), .ZN(new_n386_));
  INV_X1    g185(.A(G57gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n382_), .A2(new_n383_), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n388_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n366_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n382_), .A2(new_n383_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n388_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n395_), .A2(KEYINPUT103), .A3(new_n389_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n392_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT23), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n398_), .B1(G183gat), .B2(G190gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(KEYINPUT83), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT83), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT23), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G183gat), .A2(G190gat), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n399_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n406_));
  NOR3_X1   g205(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT96), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT26), .B(G190gat), .ZN(new_n409_));
  INV_X1    g208(.A(G183gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT25), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT25), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(G183gat), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n411_), .A2(new_n413_), .A3(KEYINPUT95), .ZN(new_n414_));
  AOI21_X1  g213(.A(KEYINPUT95), .B1(new_n411_), .B2(new_n413_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n409_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G169gat), .A2(G176gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT96), .ZN(new_n421_));
  INV_X1    g220(.A(new_n407_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n404_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n421_), .B(new_n422_), .C1(new_n423_), .C2(new_n399_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n408_), .A2(new_n416_), .A3(new_n420_), .A4(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n323_), .ZN(new_n426_));
  OR2_X1    g225(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n428_));
  AOI21_X1  g227(.A(G176gat), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(KEYINPUT82), .A2(G169gat), .A3(G176gat), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(KEYINPUT82), .B1(G169gat), .B2(G176gat), .ZN(new_n433_));
  NOR3_X1   g232(.A1(new_n432_), .A2(new_n433_), .A3(KEYINPUT97), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT97), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT82), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n419_), .A2(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n435_), .B1(new_n437_), .B2(new_n431_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n430_), .B1(new_n434_), .B2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n400_), .A2(new_n402_), .A3(new_n404_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n405_), .A2(new_n398_), .ZN(new_n441_));
  INV_X1    g240(.A(G190gat), .ZN(new_n442_));
  AOI22_X1  g241(.A1(new_n440_), .A2(new_n441_), .B1(new_n410_), .B2(new_n442_), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n439_), .A2(new_n443_), .A3(KEYINPUT98), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT98), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT97), .B1(new_n432_), .B2(new_n433_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n437_), .A2(new_n435_), .A3(new_n431_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n429_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n440_), .A2(new_n441_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n410_), .A2(new_n442_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n445_), .B1(new_n448_), .B2(new_n451_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n425_), .B(new_n426_), .C1(new_n444_), .C2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT99), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n437_), .A2(new_n431_), .ZN(new_n457_));
  AOI22_X1  g256(.A1(new_n440_), .A2(new_n441_), .B1(new_n457_), .B2(new_n418_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT80), .ZN(new_n459_));
  NAND2_X1  g258(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n459_), .B(G183gat), .C1(new_n461_), .C2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT26), .ZN(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT81), .B(G190gat), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n463_), .B(new_n411_), .C1(new_n464_), .C2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n462_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n410_), .B1(new_n467_), .B2(new_n460_), .ZN(new_n468_));
  OAI22_X1  g267(.A1(new_n468_), .A2(new_n459_), .B1(KEYINPUT26), .B2(new_n442_), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n458_), .B(new_n422_), .C1(new_n466_), .C2(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n465_), .A2(G183gat), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n457_), .B(new_n430_), .C1(new_n406_), .C2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n456_), .B1(new_n473_), .B2(new_n323_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT98), .B1(new_n439_), .B2(new_n443_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n448_), .A2(new_n451_), .A3(new_n445_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n477_), .A2(KEYINPUT99), .A3(new_n426_), .A4(new_n425_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n455_), .A2(new_n474_), .A3(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G226gat), .A2(G233gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT19), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n479_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n477_), .A2(new_n425_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n323_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n470_), .A2(new_n426_), .A3(new_n472_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n485_), .A2(new_n486_), .A3(KEYINPUT20), .A4(new_n481_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n483_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G8gat), .B(G36gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G64gat), .B(G92gat), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n491_), .B(new_n492_), .Z(new_n493_));
  NAND2_X1  g292(.A1(new_n488_), .A2(new_n493_), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n425_), .B(new_n426_), .C1(new_n443_), .C2(new_n439_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n482_), .B1(new_n474_), .B2(new_n495_), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n485_), .A2(KEYINPUT20), .A3(new_n486_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n496_), .B1(new_n497_), .B2(new_n482_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n494_), .B(KEYINPUT27), .C1(new_n493_), .C2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n493_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n483_), .A2(new_n487_), .A3(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n494_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT27), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT104), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n483_), .A2(new_n487_), .A3(new_n500_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n500_), .B1(new_n483_), .B2(new_n487_), .ZN(new_n506_));
  OAI211_X1 g305(.A(KEYINPUT104), .B(new_n503_), .C1(new_n505_), .C2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n397_), .B(new_n499_), .C1(new_n504_), .C2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n365_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n361_), .A2(new_n364_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT33), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n389_), .A2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n502_), .A2(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n367_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n377_), .A2(new_n378_), .A3(new_n369_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n515_), .A2(new_n394_), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT102), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n390_), .A2(new_n518_), .A3(KEYINPUT33), .ZN(new_n519_));
  AOI21_X1  g318(.A(KEYINPUT102), .B1(new_n389_), .B2(new_n512_), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n514_), .B(new_n517_), .C1(new_n519_), .C2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n493_), .A2(KEYINPUT32), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n488_), .A2(new_n522_), .ZN(new_n523_));
  OAI221_X1 g322(.A(new_n523_), .B1(new_n498_), .B2(new_n522_), .C1(new_n390_), .C2(new_n391_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n511_), .A2(new_n521_), .A3(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G15gat), .B(G71gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n376_), .B(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G227gat), .A2(G233gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT30), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n527_), .B(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(KEYINPUT84), .B(G43gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT31), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(G99gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n473_), .B(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n530_), .B(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n510_), .A2(new_n525_), .A3(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n499_), .B1(new_n504_), .B2(new_n508_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT105), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  OAI211_X1 g339(.A(KEYINPUT105), .B(new_n499_), .C1(new_n504_), .C2(new_n508_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n397_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n542_), .A2(new_n536_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n540_), .A2(new_n511_), .A3(new_n541_), .A4(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n279_), .B1(new_n537_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G229gat), .A2(G233gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G29gat), .B(G36gat), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT71), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(G43gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(G50gat), .ZN(new_n551_));
  INV_X1    g350(.A(G43gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n549_), .B(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(G50gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n551_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G15gat), .B(G22gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT72), .ZN(new_n558_));
  INV_X1    g357(.A(G1gat), .ZN(new_n559_));
  INV_X1    g358(.A(G8gat), .ZN(new_n560_));
  OAI21_X1  g359(.A(KEYINPUT14), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT73), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n558_), .A2(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(G1gat), .B(G8gat), .Z(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n556_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT15), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n556_), .B(new_n567_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n546_), .B(new_n566_), .C1(new_n568_), .C2(new_n565_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n546_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n566_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n556_), .A2(new_n565_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n570_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G113gat), .B(G141gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT77), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(G169gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(new_n309_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n569_), .A2(new_n573_), .A3(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n578_), .B1(new_n569_), .B2(new_n573_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT78), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT78), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n583_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n545_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(G134gat), .ZN(new_n589_));
  INV_X1    g388(.A(G162gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT36), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G232gat), .A2(G233gat), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT69), .Z(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT34), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n596_), .A2(KEYINPUT35), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n556_), .A2(new_n253_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n239_), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n597_), .B(new_n598_), .C1(new_n568_), .C2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n596_), .A2(KEYINPUT35), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT70), .Z(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n556_), .B(KEYINPUT15), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(new_n239_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n602_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n605_), .A2(new_n606_), .A3(new_n597_), .A4(new_n598_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n593_), .B1(new_n603_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT37), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT36), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n591_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n603_), .A2(new_n607_), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n609_), .B(new_n610_), .C1(new_n612_), .C2(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n612_), .ZN(new_n615_));
  OAI21_X1  g414(.A(KEYINPUT37), .B1(new_n615_), .B2(new_n608_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n565_), .B(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(new_n254_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G183gat), .B(G211gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G127gat), .B(G155gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n621_), .B1(KEYINPUT17), .B2(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n627_), .B1(KEYINPUT17), .B2(new_n626_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n626_), .A2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT76), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n621_), .A2(new_n631_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n628_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n618_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n587_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT106), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n638_), .A2(new_n559_), .A3(new_n542_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT38), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT107), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n639_), .A2(new_n640_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n639_), .A2(KEYINPUT107), .A3(new_n640_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n615_), .A2(new_n608_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n646_), .B1(new_n537_), .B2(new_n544_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n279_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n581_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n650_), .A2(new_n634_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n647_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(new_n542_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(G1gat), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n643_), .A2(new_n644_), .A3(new_n645_), .A4(new_n654_), .ZN(G1324gat));
  NAND2_X1  g454(.A1(new_n540_), .A2(new_n541_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n647_), .A2(new_n656_), .A3(new_n651_), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n657_), .A2(KEYINPUT108), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(KEYINPUT108), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n658_), .A2(G8gat), .A3(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT109), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n658_), .A2(KEYINPUT109), .A3(G8gat), .A4(new_n659_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n662_), .A2(KEYINPUT39), .A3(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n638_), .A2(new_n560_), .A3(new_n656_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT39), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n660_), .A2(new_n661_), .A3(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n664_), .A2(new_n665_), .A3(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT40), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n664_), .A2(new_n665_), .A3(KEYINPUT40), .A4(new_n667_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1325gat));
  INV_X1    g471(.A(G15gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n638_), .A2(new_n673_), .A3(new_n535_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n652_), .B2(new_n535_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT41), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(G1326gat));
  INV_X1    g476(.A(G22gat), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n638_), .A2(new_n678_), .A3(new_n365_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n678_), .B1(new_n652_), .B2(new_n365_), .ZN(new_n680_));
  XOR2_X1   g479(.A(KEYINPUT110), .B(KEYINPUT42), .Z(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n679_), .A2(new_n682_), .ZN(G1327gat));
  INV_X1    g482(.A(new_n646_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n684_), .A2(new_n633_), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n545_), .A2(new_n586_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(G29gat), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n686_), .A2(new_n687_), .A3(new_n542_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n537_), .A2(new_n544_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n618_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT43), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n689_), .A2(new_n692_), .A3(new_n618_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT111), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT44), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n695_), .A2(KEYINPUT44), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n650_), .A2(new_n633_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n694_), .A2(new_n696_), .A3(new_n697_), .A4(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n692_), .B1(new_n689_), .B2(new_n618_), .ZN(new_n700_));
  AOI211_X1 g499(.A(KEYINPUT43), .B(new_n617_), .C1(new_n537_), .C2(new_n544_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n698_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n702_), .A2(new_n695_), .A3(KEYINPUT44), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n699_), .A2(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n687_), .B1(new_n704_), .B2(new_n542_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT112), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n705_), .A2(new_n706_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n688_), .B1(new_n707_), .B2(new_n708_), .ZN(G1328gat));
  INV_X1    g508(.A(G36gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n710_), .B1(new_n704_), .B2(new_n656_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n686_), .A2(new_n710_), .A3(new_n656_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT113), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT113), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n686_), .A2(new_n715_), .A3(new_n710_), .A4(new_n656_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n714_), .A2(KEYINPUT45), .A3(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n714_), .A2(new_n716_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n712_), .A2(KEYINPUT46), .A3(new_n717_), .A4(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT46), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n717_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(new_n723_), .B2(new_n711_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n721_), .A2(new_n724_), .ZN(G1329gat));
  AOI21_X1  g524(.A(new_n552_), .B1(new_n704_), .B2(new_n535_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n686_), .A2(new_n552_), .A3(new_n535_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  OR3_X1    g527(.A1(new_n726_), .A2(KEYINPUT47), .A3(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT47), .B1(new_n726_), .B2(new_n728_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1330gat));
  AOI21_X1  g530(.A(new_n554_), .B1(new_n704_), .B2(new_n365_), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n686_), .A2(new_n554_), .A3(new_n365_), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1331gat));
  NAND4_X1  g533(.A1(new_n647_), .A2(new_n633_), .A3(new_n585_), .A4(new_n279_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n735_), .A2(new_n387_), .A3(new_n397_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT114), .Z(new_n737_));
  NOR2_X1   g536(.A1(new_n648_), .A2(new_n649_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n537_), .B2(new_n544_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(new_n635_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n387_), .B1(new_n741_), .B2(new_n397_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n737_), .A2(new_n742_), .ZN(G1332gat));
  INV_X1    g542(.A(new_n656_), .ZN(new_n744_));
  OAI21_X1  g543(.A(G64gat), .B1(new_n735_), .B2(new_n744_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(KEYINPUT115), .B(KEYINPUT48), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n745_), .B(new_n746_), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n744_), .A2(G64gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n741_), .B2(new_n748_), .ZN(G1333gat));
  OAI21_X1  g548(.A(G71gat), .B1(new_n735_), .B2(new_n536_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT49), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n536_), .A2(G71gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n741_), .B2(new_n752_), .ZN(G1334gat));
  OAI21_X1  g552(.A(G78gat), .B1(new_n735_), .B2(new_n511_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT50), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n511_), .A2(G78gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n755_), .B1(new_n741_), .B2(new_n756_), .ZN(G1335gat));
  AND2_X1   g556(.A1(new_n740_), .A2(new_n685_), .ZN(new_n758_));
  AOI21_X1  g557(.A(G85gat), .B1(new_n758_), .B2(new_n542_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n739_), .A2(new_n633_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n694_), .A2(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n397_), .A2(new_n214_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n759_), .B1(new_n761_), .B2(new_n762_), .ZN(G1336gat));
  AOI21_X1  g562(.A(G92gat), .B1(new_n758_), .B2(new_n656_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n744_), .A2(new_n215_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n761_), .B2(new_n765_), .ZN(G1337gat));
  NAND2_X1  g565(.A1(new_n761_), .A2(new_n535_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(G99gat), .ZN(new_n768_));
  INV_X1    g567(.A(new_n202_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n758_), .A2(new_n769_), .A3(new_n535_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g571(.A(KEYINPUT116), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n694_), .A2(new_n773_), .A3(new_n365_), .A4(new_n760_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n365_), .B(new_n760_), .C1(new_n700_), .C2(new_n701_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT116), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n774_), .A2(new_n776_), .A3(G106gat), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT52), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n774_), .A2(new_n776_), .A3(new_n779_), .A4(G106gat), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(G106gat), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n758_), .A2(new_n782_), .A3(new_n365_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT53), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n781_), .A2(new_n786_), .A3(new_n783_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(G1339gat));
  INV_X1    g587(.A(KEYINPUT117), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n633_), .A2(new_n582_), .A3(new_n584_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n789_), .B1(new_n790_), .B2(new_n279_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n585_), .A2(KEYINPUT117), .A3(new_n633_), .A4(new_n648_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n792_), .A3(new_n617_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT54), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n248_), .B(new_n263_), .C1(new_n258_), .C2(new_n261_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n249_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n262_), .A2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n257_), .B1(new_n256_), .B2(KEYINPUT12), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n259_), .A2(KEYINPUT67), .A3(new_n260_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n801_), .A2(KEYINPUT55), .A3(new_n255_), .A4(new_n248_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n796_), .A2(new_n798_), .A3(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n803_), .A2(KEYINPUT56), .A3(new_n271_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n271_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT56), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT118), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT118), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n806_), .A2(new_n810_), .A3(new_n807_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n805_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n649_), .A2(new_n273_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT119), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n570_), .B(new_n566_), .C1(new_n568_), .C2(new_n565_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n546_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n579_), .B1(new_n577_), .B2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n275_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n810_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n820_));
  AOI211_X1 g619(.A(KEYINPUT118), .B(KEYINPUT56), .C1(new_n803_), .C2(new_n271_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n804_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT119), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n822_), .A2(new_n823_), .A3(new_n649_), .A4(new_n273_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n814_), .A2(new_n819_), .A3(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT120), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n826_), .A2(KEYINPUT57), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  AND3_X1   g627(.A1(new_n825_), .A2(new_n684_), .A3(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n825_), .B2(new_n684_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n808_), .A2(new_n804_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n818_), .A2(new_n831_), .A3(new_n273_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT58), .ZN(new_n833_));
  OR2_X1    g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n833_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n834_), .A2(new_n618_), .A3(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n829_), .A2(new_n830_), .A3(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n794_), .B1(new_n838_), .B2(new_n633_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n744_), .A2(new_n511_), .A3(new_n535_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n839_), .A2(new_n542_), .A3(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(G113gat), .B1(new_n843_), .B2(new_n649_), .ZN(new_n844_));
  AND2_X1   g643(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n845_));
  NOR2_X1   g644(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n842_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n825_), .A2(new_n684_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n827_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n825_), .A2(new_n684_), .A3(new_n828_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n850_), .A2(new_n836_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n634_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n397_), .B1(new_n853_), .B2(new_n794_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n854_), .A2(new_n841_), .A3(new_n845_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n585_), .B1(new_n848_), .B2(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n844_), .B1(new_n856_), .B2(G113gat), .ZN(G1340gat));
  XOR2_X1   g656(.A(KEYINPUT122), .B(G120gat), .Z(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n648_), .B2(KEYINPUT60), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n843_), .B(new_n859_), .C1(KEYINPUT60), .C2(new_n858_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n648_), .B1(new_n848_), .B2(new_n855_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(new_n858_), .ZN(G1341gat));
  AOI21_X1  g661(.A(G127gat), .B1(new_n843_), .B2(new_n633_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n634_), .B1(new_n848_), .B2(new_n855_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g664(.A(G134gat), .B1(new_n843_), .B2(new_n646_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n617_), .B1(new_n848_), .B2(new_n855_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(G134gat), .ZN(G1343gat));
  NOR2_X1   g667(.A1(new_n511_), .A2(new_n535_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n839_), .A2(new_n542_), .A3(new_n744_), .A4(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n870_), .A2(new_n581_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(KEYINPUT123), .B(G141gat), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(G1344gat));
  NOR2_X1   g672(.A1(new_n870_), .A2(new_n648_), .ZN(new_n874_));
  INV_X1    g673(.A(G148gat), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1345gat));
  NOR2_X1   g675(.A1(new_n870_), .A2(new_n634_), .ZN(new_n877_));
  XOR2_X1   g676(.A(KEYINPUT61), .B(G155gat), .Z(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1346gat));
  NOR3_X1   g678(.A1(new_n870_), .A2(new_n590_), .A3(new_n617_), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n870_), .A2(new_n684_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(new_n590_), .ZN(G1347gat));
  AOI21_X1  g681(.A(new_n744_), .B1(new_n853_), .B2(new_n794_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n543_), .A2(new_n511_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n883_), .A2(new_n649_), .A3(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n886_), .A2(new_n887_), .A3(G169gat), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n886_), .B2(G169gat), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n883_), .A2(new_n885_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n581_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n891_));
  XOR2_X1   g690(.A(new_n891_), .B(KEYINPUT124), .Z(new_n892_));
  OAI22_X1  g691(.A1(new_n888_), .A2(new_n889_), .B1(new_n890_), .B2(new_n892_), .ZN(G1348gat));
  NAND3_X1  g692(.A1(new_n883_), .A2(new_n279_), .A3(new_n885_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(G176gat), .ZN(G1349gat));
  OAI22_X1  g694(.A1(new_n414_), .A2(new_n415_), .B1(KEYINPUT125), .B2(G183gat), .ZN(new_n896_));
  OR3_X1    g695(.A1(new_n890_), .A2(new_n634_), .A3(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n890_), .A2(new_n634_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n410_), .A2(KEYINPUT125), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n897_), .B1(new_n898_), .B2(new_n899_), .ZN(G1350gat));
  OAI21_X1  g699(.A(G190gat), .B1(new_n890_), .B2(new_n617_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n646_), .A2(new_n409_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n890_), .B2(new_n902_), .ZN(G1351gat));
  NAND2_X1  g702(.A1(new_n869_), .A2(new_n397_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(KEYINPUT126), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n883_), .A2(new_n649_), .A3(new_n906_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G197gat), .ZN(G1352gat));
  AND2_X1   g707(.A1(new_n883_), .A2(new_n906_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(new_n279_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(G204gat), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n909_), .A2(new_n312_), .A3(new_n279_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1353gat));
  NAND4_X1  g712(.A1(new_n839_), .A2(new_n633_), .A3(new_n656_), .A4(new_n906_), .ZN(new_n914_));
  OR2_X1    g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT127), .ZN(new_n917_));
  XNOR2_X1  g716(.A(KEYINPUT63), .B(G211gat), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n883_), .A2(new_n633_), .A3(new_n906_), .A4(new_n918_), .ZN(new_n919_));
  AND3_X1   g718(.A1(new_n916_), .A2(new_n917_), .A3(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n917_), .B1(new_n916_), .B2(new_n919_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n920_), .A2(new_n921_), .ZN(G1354gat));
  AOI21_X1  g721(.A(G218gat), .B1(new_n909_), .B2(new_n646_), .ZN(new_n923_));
  AND2_X1   g722(.A1(new_n618_), .A2(G218gat), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n923_), .B1(new_n909_), .B2(new_n924_), .ZN(G1355gat));
endmodule


