//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 0 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1 0 0 1 0 0 0 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_, new_n931_, new_n932_, new_n933_, new_n935_, new_n937_,
    new_n938_, new_n940_, new_n941_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n959_,
    new_n960_, new_n961_, new_n963_, new_n964_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n972_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n980_, new_n981_;
  XNOR2_X1  g000(.A(G22gat), .B(G50gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G228gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT94), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT29), .ZN(new_n206_));
  AND2_X1   g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208_));
  NOR3_X1   g007(.A1(new_n207_), .A2(new_n208_), .A3(KEYINPUT1), .ZN(new_n209_));
  OR2_X1    g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT92), .B1(new_n209_), .B2(new_n213_), .ZN(new_n214_));
  OR2_X1    g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n212_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT92), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n218_), .A2(new_n221_), .A3(new_n222_), .A4(new_n211_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n214_), .A2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n207_), .A2(new_n208_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n220_), .A2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n227_), .B(new_n228_), .C1(KEYINPUT2), .C2(new_n219_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT93), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n225_), .B1(new_n229_), .B2(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n206_), .B1(new_n224_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(G211gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n236_), .A2(G218gat), .ZN(new_n237_));
  INV_X1    g036(.A(G218gat), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n238_), .A2(G211gat), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT98), .B1(new_n237_), .B2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(G211gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n236_), .A2(G218gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT98), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(G197gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G204gat), .ZN(new_n246_));
  INV_X1    g045(.A(G204gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(G197gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  AOI22_X1  g048(.A1(new_n240_), .A2(new_n244_), .B1(KEYINPUT21), .B2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT96), .B1(new_n247_), .B2(G197gat), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT96), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n252_), .A2(new_n245_), .A3(G204gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT21), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n251_), .A2(new_n253_), .A3(new_n254_), .A4(new_n248_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT97), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n255_), .A2(KEYINPUT97), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n250_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n251_), .A2(new_n253_), .A3(new_n248_), .ZN(new_n260_));
  AND4_X1   g059(.A1(KEYINPUT21), .A2(new_n240_), .A3(new_n260_), .A4(new_n244_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n259_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT95), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n235_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT99), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NOR3_X1   g066(.A1(new_n247_), .A2(KEYINPUT96), .A3(G197gat), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n245_), .A2(G204gat), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT97), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n270_), .A2(new_n271_), .A3(new_n254_), .A4(new_n251_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n256_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n261_), .B1(new_n273_), .B2(new_n250_), .ZN(new_n274_));
  NOR3_X1   g073(.A1(new_n274_), .A2(new_n234_), .A3(new_n266_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n205_), .B1(new_n267_), .B2(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n274_), .A2(new_n234_), .ZN(new_n278_));
  AOI21_X1  g077(.A(KEYINPUT99), .B1(new_n278_), .B2(new_n264_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n279_), .A2(new_n204_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n202_), .B1(new_n277_), .B2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n224_), .A2(new_n233_), .A3(new_n206_), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n282_), .A2(KEYINPUT28), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(KEYINPUT28), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G78gat), .B(G106gat), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n283_), .A2(new_n284_), .A3(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n286_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n204_), .B1(new_n279_), .B2(new_n275_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n267_), .A2(new_n205_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n202_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  AND3_X1   g092(.A1(new_n281_), .A2(new_n289_), .A3(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n289_), .B1(new_n281_), .B2(new_n293_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G1gat), .B(G29gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(G85gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT0), .B(G57gat), .ZN(new_n299_));
  XOR2_X1   g098(.A(new_n298_), .B(new_n299_), .Z(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n224_), .A2(new_n233_), .ZN(new_n302_));
  XOR2_X1   g101(.A(G113gat), .B(G120gat), .Z(new_n303_));
  INV_X1    g102(.A(G134gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(G127gat), .ZN(new_n305_));
  INV_X1    g104(.A(G127gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(G134gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT89), .ZN(new_n308_));
  AND3_X1   g107(.A1(new_n305_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n308_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n303_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n306_), .A2(G134gat), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n304_), .A2(G127gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT89), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n305_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G113gat), .B(G120gat), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  AND3_X1   g116(.A1(new_n311_), .A2(KEYINPUT90), .A3(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(KEYINPUT90), .B1(new_n311_), .B2(new_n317_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n302_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G225gat), .A2(G233gat), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n224_), .A2(new_n233_), .A3(new_n317_), .A4(new_n311_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT103), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT103), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n320_), .A2(new_n325_), .A3(new_n321_), .A4(new_n322_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT90), .ZN(new_n328_));
  NOR3_X1   g127(.A1(new_n309_), .A2(new_n310_), .A3(new_n303_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n316_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n328_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n311_), .A2(new_n317_), .A3(KEYINPUT90), .ZN(new_n332_));
  AOI22_X1  g131(.A1(new_n331_), .A2(new_n332_), .B1(new_n224_), .B2(new_n233_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n322_), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT4), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT4), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n320_), .A2(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n321_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n301_), .B1(new_n327_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT106), .ZN(new_n340_));
  INV_X1    g139(.A(new_n321_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n336_), .B1(new_n320_), .B2(new_n322_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n331_), .A2(new_n332_), .ZN(new_n343_));
  AOI21_X1  g142(.A(KEYINPUT4), .B1(new_n343_), .B2(new_n302_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n341_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n345_), .A2(new_n300_), .A3(new_n324_), .A4(new_n326_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n339_), .A2(new_n340_), .A3(new_n346_), .ZN(new_n347_));
  OAI211_X1 g146(.A(KEYINPUT106), .B(new_n301_), .C1(new_n327_), .C2(new_n338_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(G169gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G183gat), .A2(G190gat), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT23), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n355_), .B(new_n356_), .C1(G183gat), .C2(G190gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n352_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT26), .B(G190gat), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT87), .ZN(new_n360_));
  INV_X1    g159(.A(G183gat), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n360_), .B1(new_n361_), .B2(KEYINPUT25), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT25), .B(G183gat), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n359_), .B(new_n362_), .C1(new_n363_), .C2(new_n360_), .ZN(new_n364_));
  INV_X1    g163(.A(G169gat), .ZN(new_n365_));
  INV_X1    g164(.A(G176gat), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(new_n366_), .A3(KEYINPUT88), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT88), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n368_), .B1(G169gat), .B2(G176gat), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT24), .B1(new_n367_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n364_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G169gat), .A2(G176gat), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n367_), .A2(new_n369_), .A3(KEYINPUT24), .A4(new_n373_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n355_), .A2(new_n356_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n358_), .B1(new_n372_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G227gat), .A2(G233gat), .ZN(new_n378_));
  INV_X1    g177(.A(G15gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT30), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n377_), .B(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(new_n343_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G71gat), .B(G99gat), .ZN(new_n384_));
  INV_X1    g183(.A(G43gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT31), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n383_), .B(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT27), .ZN(new_n390_));
  INV_X1    g189(.A(G190gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT26), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT26), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(G190gat), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n362_), .A2(new_n392_), .A3(new_n394_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n361_), .A2(KEYINPUT25), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n361_), .A2(KEYINPUT25), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT87), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n370_), .B1(new_n395_), .B2(new_n398_), .ZN(new_n399_));
  AND2_X1   g198(.A1(new_n374_), .A2(new_n375_), .ZN(new_n400_));
  AOI22_X1  g199(.A1(new_n399_), .A2(new_n400_), .B1(new_n357_), .B2(new_n352_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT102), .B1(new_n274_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT102), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n249_), .A2(KEYINPUT21), .ZN(new_n404_));
  INV_X1    g203(.A(new_n244_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n243_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n404_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n407_), .B1(new_n256_), .B2(new_n272_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n377_), .B(new_n403_), .C1(new_n408_), .C2(new_n261_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n402_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT100), .B(KEYINPUT19), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G226gat), .A2(G233gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT20), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n363_), .A2(new_n359_), .ZN(new_n416_));
  OR3_X1    g215(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n416_), .A2(new_n374_), .A3(new_n375_), .A4(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n373_), .B(KEYINPUT101), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT22), .B(G169gat), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n357_), .B(new_n419_), .C1(new_n421_), .C2(G176gat), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n418_), .A2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n415_), .B1(new_n274_), .B2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n410_), .A2(new_n414_), .A3(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(G8gat), .B(G36gat), .Z(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT18), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G64gat), .B(G92gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n263_), .A2(new_n377_), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT20), .B1(new_n274_), .B2(new_n423_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n413_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n425_), .A2(new_n429_), .A3(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n429_), .B1(new_n425_), .B2(new_n432_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n390_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n429_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n414_), .B1(new_n410_), .B2(new_n424_), .ZN(new_n437_));
  NOR3_X1   g236(.A1(new_n430_), .A2(new_n431_), .A3(new_n413_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n436_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n425_), .A2(new_n429_), .A3(new_n432_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(KEYINPUT27), .A3(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n435_), .A2(new_n441_), .ZN(new_n442_));
  NOR4_X1   g241(.A1(new_n296_), .A2(new_n350_), .A3(new_n389_), .A4(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n289_), .ZN(new_n444_));
  NOR3_X1   g243(.A1(new_n277_), .A2(new_n280_), .A3(new_n202_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n292_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n444_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n281_), .A2(new_n293_), .A3(new_n289_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT33), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n346_), .A2(KEYINPUT104), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n425_), .A2(new_n432_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n436_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n321_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT105), .B1(new_n320_), .B2(new_n322_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n320_), .A2(KEYINPUT105), .A3(new_n322_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n341_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n455_), .B(new_n301_), .C1(new_n456_), .C2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n454_), .A2(new_n440_), .A3(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n450_), .B1(new_n346_), .B2(KEYINPUT104), .ZN(new_n461_));
  NOR3_X1   g260(.A1(new_n452_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n429_), .A2(KEYINPUT32), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n464_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n425_), .A2(new_n432_), .A3(new_n463_), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n467_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n449_), .B1(new_n462_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT107), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n447_), .A2(new_n448_), .A3(new_n435_), .A4(new_n441_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n470_), .B1(new_n471_), .B2(new_n350_), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n435_), .A2(new_n441_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n296_), .A2(new_n473_), .A3(KEYINPUT107), .A4(new_n349_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n469_), .A2(new_n472_), .A3(new_n474_), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n388_), .B(KEYINPUT91), .Z(new_n476_));
  AOI21_X1  g275(.A(new_n443_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(G1gat), .B(G8gat), .Z(new_n478_));
  INV_X1    g277(.A(G1gat), .ZN(new_n479_));
  INV_X1    g278(.A(G8gat), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT14), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT78), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT78), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n483_), .B(KEYINPUT14), .C1(new_n479_), .C2(new_n480_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G15gat), .B(G22gat), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n482_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT79), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT79), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n482_), .A2(new_n488_), .A3(new_n484_), .A4(new_n485_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n478_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n487_), .A2(new_n478_), .A3(new_n489_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G29gat), .B(G36gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G43gat), .B(G50gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT15), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n493_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT83), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n496_), .B(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G229gat), .A2(G233gat), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n502_), .B(KEYINPUT85), .Z(new_n503_));
  NAND3_X1  g302(.A1(new_n498_), .A2(new_n501_), .A3(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n496_), .B(KEYINPUT83), .ZN(new_n505_));
  INV_X1    g304(.A(new_n492_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n505_), .B1(new_n506_), .B2(new_n490_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(new_n501_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n502_), .ZN(new_n509_));
  AOI21_X1  g308(.A(KEYINPUT84), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT84), .ZN(new_n511_));
  AOI211_X1 g310(.A(new_n511_), .B(new_n502_), .C1(new_n507_), .C2(new_n501_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n504_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(G113gat), .B(G141gat), .Z(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT86), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G169gat), .B(G197gat), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n515_), .B(new_n516_), .Z(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n513_), .A2(new_n518_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n504_), .B(new_n517_), .C1(new_n510_), .C2(new_n512_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n477_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G190gat), .B(G218gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G134gat), .B(G162gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n526_), .B(KEYINPUT36), .Z(new_n527_));
  INV_X1    g326(.A(KEYINPUT35), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT75), .B(KEYINPUT34), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G232gat), .A2(G233gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G85gat), .A2(G92gat), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT64), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT9), .ZN(new_n535_));
  AND3_X1   g334(.A1(new_n533_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n534_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(G85gat), .A2(G92gat), .ZN(new_n539_));
  OAI22_X1  g338(.A1(new_n539_), .A2(KEYINPUT65), .B1(new_n533_), .B2(new_n535_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT65), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n541_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(KEYINPUT66), .B1(new_n538_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n533_), .A2(new_n535_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT64), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n533_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT66), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n548_), .A2(new_n549_), .A3(new_n542_), .A4(new_n540_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n544_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G99gat), .A2(G106gat), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT67), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n553_), .A2(KEYINPUT6), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT6), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n555_), .A2(KEYINPUT67), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n552_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(KEYINPUT67), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n553_), .A2(KEYINPUT6), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n558_), .A2(new_n559_), .A3(G99gat), .A4(G106gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n557_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(KEYINPUT10), .B(G99gat), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n562_), .A2(G106gat), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(G99gat), .ZN(new_n566_));
  INV_X1    g365(.A(G106gat), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n566_), .A2(new_n567_), .A3(KEYINPUT68), .A4(KEYINPUT7), .ZN(new_n568_));
  NAND2_X1  g367(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n569_), .B1(G99gat), .B2(G106gat), .ZN(new_n570_));
  NOR2_X1   g369(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n568_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n572_), .A2(new_n560_), .A3(new_n557_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(KEYINPUT69), .A2(KEYINPUT8), .ZN(new_n574_));
  INV_X1    g373(.A(new_n533_), .ZN(new_n575_));
  AOI211_X1 g374(.A(new_n539_), .B(new_n575_), .C1(KEYINPUT69), .C2(KEYINPUT8), .ZN(new_n576_));
  AND3_X1   g375(.A1(new_n573_), .A2(new_n574_), .A3(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n574_), .B1(new_n573_), .B2(new_n576_), .ZN(new_n578_));
  OAI22_X1  g377(.A1(new_n551_), .A2(new_n565_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(new_n497_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT76), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n573_), .A2(new_n576_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n574_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n573_), .A2(new_n574_), .A3(new_n576_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n544_), .A2(new_n550_), .ZN(new_n587_));
  AOI22_X1  g386(.A1(new_n585_), .A2(new_n586_), .B1(new_n587_), .B2(new_n564_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(new_n496_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT77), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  AOI211_X1 g390(.A(new_n528_), .B(new_n532_), .C1(new_n582_), .C2(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n532_), .A2(new_n528_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n532_), .A2(new_n528_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n582_), .A2(new_n591_), .A3(new_n594_), .A4(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n527_), .B1(new_n592_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT37), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n582_), .A2(new_n591_), .A3(new_n595_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(new_n593_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n526_), .A2(KEYINPUT36), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(new_n602_), .A3(new_n596_), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n598_), .A2(new_n599_), .A3(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n599_), .B1(new_n598_), .B2(new_n603_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(G230gat), .ZN(new_n607_));
  INV_X1    g406(.A(G233gat), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G57gat), .B(G64gat), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT11), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT71), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT71), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n610_), .A2(new_n613_), .A3(KEYINPUT11), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  OR2_X1    g414(.A1(KEYINPUT70), .A2(G71gat), .ZN(new_n616_));
  NAND2_X1  g415(.A1(KEYINPUT70), .A2(G71gat), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(G78gat), .ZN(new_n619_));
  INV_X1    g418(.A(G78gat), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n616_), .A2(new_n620_), .A3(new_n617_), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n619_), .B(new_n621_), .C1(KEYINPUT11), .C2(new_n610_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n615_), .A2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n615_), .A2(new_n622_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n609_), .B1(new_n588_), .B2(new_n625_), .ZN(new_n626_));
  NOR3_X1   g425(.A1(new_n588_), .A2(new_n625_), .A3(KEYINPUT12), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT12), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n615_), .B(new_n622_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n628_), .B1(new_n579_), .B2(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n626_), .B1(new_n627_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n609_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n588_), .B(new_n629_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n631_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(G176gat), .B(G204gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT73), .ZN(new_n636_));
  XOR2_X1   g435(.A(KEYINPUT72), .B(KEYINPUT5), .Z(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  XOR2_X1   g437(.A(G120gat), .B(G148gat), .Z(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n634_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT74), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n634_), .A2(new_n641_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n642_), .A2(new_n643_), .A3(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n634_), .A2(KEYINPUT74), .A3(new_n641_), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n645_), .A2(KEYINPUT13), .A3(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT13), .B1(new_n645_), .B2(new_n646_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(G231gat), .A2(G233gat), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n650_), .B(KEYINPUT80), .Z(new_n651_));
  XNOR2_X1  g450(.A(new_n493_), .B(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(new_n625_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  XOR2_X1   g453(.A(G183gat), .B(G211gat), .Z(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT82), .ZN(new_n656_));
  XOR2_X1   g455(.A(G127gat), .B(G155gat), .Z(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(new_n657_), .ZN(new_n658_));
  XOR2_X1   g457(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n659_));
  XNOR2_X1  g458(.A(new_n658_), .B(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n654_), .A2(KEYINPUT17), .A3(new_n660_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n660_), .B(KEYINPUT17), .Z(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(new_n653_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n606_), .A2(new_n649_), .A3(new_n664_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n523_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n666_), .A2(new_n479_), .A3(new_n350_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT38), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n475_), .A2(new_n476_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n443_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n598_), .A2(new_n603_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n649_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n664_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n675_), .A2(new_n521_), .A3(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n674_), .A2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n479_), .B1(new_n678_), .B2(new_n350_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n669_), .A2(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n680_), .B1(new_n668_), .B2(new_n667_), .ZN(G1324gat));
  NAND3_X1  g480(.A1(new_n666_), .A2(new_n480_), .A3(new_n442_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT108), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n678_), .A2(new_n442_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT39), .ZN(new_n685_));
  AND4_X1   g484(.A1(new_n683_), .A2(new_n684_), .A3(new_n685_), .A4(G8gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n480_), .B1(KEYINPUT108), .B2(KEYINPUT39), .ZN(new_n687_));
  AOI22_X1  g486(.A1(new_n684_), .A2(new_n687_), .B1(new_n683_), .B2(new_n685_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n682_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT40), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(G1325gat));
  INV_X1    g490(.A(new_n476_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n379_), .B1(new_n678_), .B2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT41), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n666_), .A2(new_n379_), .A3(new_n692_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1326gat));
  INV_X1    g495(.A(G22gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n697_), .B1(new_n678_), .B2(new_n296_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT42), .Z(new_n699_));
  NAND3_X1  g498(.A1(new_n666_), .A2(new_n697_), .A3(new_n296_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1327gat));
  INV_X1    g500(.A(new_n673_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(new_n664_), .ZN(new_n703_));
  NOR4_X1   g502(.A1(new_n477_), .A2(new_n522_), .A3(new_n649_), .A4(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(G29gat), .B1(new_n704_), .B2(new_n350_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n296_), .A2(new_n473_), .A3(new_n349_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n467_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n346_), .A2(KEYINPUT104), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT33), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(new_n451_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n708_), .B1(new_n711_), .B2(new_n460_), .ZN(new_n712_));
  AOI22_X1  g511(.A1(new_n707_), .A2(new_n470_), .B1(new_n712_), .B2(new_n449_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n692_), .B1(new_n713_), .B2(new_n474_), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n706_), .B(new_n606_), .C1(new_n714_), .C2(new_n443_), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n604_), .A2(new_n605_), .ZN(new_n716_));
  OAI21_X1  g515(.A(KEYINPUT43), .B1(new_n477_), .B2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n675_), .A2(new_n521_), .A3(new_n664_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT44), .B1(new_n718_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722_));
  AOI211_X1 g521(.A(new_n722_), .B(new_n719_), .C1(new_n715_), .C2(new_n717_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n721_), .A2(new_n723_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n350_), .A2(G29gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n705_), .B1(new_n724_), .B2(new_n725_), .ZN(G1328gat));
  INV_X1    g525(.A(KEYINPUT109), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT46), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n730_));
  INV_X1    g529(.A(G36gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n724_), .B2(new_n442_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n704_), .A2(new_n731_), .A3(new_n442_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT45), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n729_), .B(new_n730_), .C1(new_n732_), .C2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n721_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n718_), .A2(KEYINPUT44), .A3(new_n720_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n737_), .A2(new_n442_), .A3(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(G36gat), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n740_), .A2(new_n727_), .A3(new_n734_), .A4(new_n728_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n736_), .A2(new_n741_), .ZN(G1329gat));
  AOI21_X1  g541(.A(G43gat), .B1(new_n704_), .B2(new_n692_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n389_), .A2(new_n385_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n724_), .B2(new_n744_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g545(.A(G50gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n704_), .A2(new_n747_), .A3(new_n296_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n724_), .A2(KEYINPUT110), .A3(new_n296_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(G50gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT110), .B1(new_n724_), .B2(new_n296_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n748_), .B1(new_n750_), .B2(new_n751_), .ZN(G1331gat));
  NOR3_X1   g551(.A1(new_n477_), .A2(new_n521_), .A3(new_n675_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n606_), .A2(new_n664_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(G57gat), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n755_), .A2(new_n756_), .A3(new_n350_), .ZN(new_n757_));
  NOR4_X1   g556(.A1(new_n674_), .A2(new_n521_), .A3(new_n675_), .A4(new_n664_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n758_), .A2(new_n350_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n757_), .B1(new_n759_), .B2(new_n756_), .ZN(G1332gat));
  INV_X1    g559(.A(G64gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n761_), .B1(new_n758_), .B2(new_n442_), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT48), .Z(new_n763_));
  NAND3_X1  g562(.A1(new_n755_), .A2(new_n761_), .A3(new_n442_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(G1333gat));
  INV_X1    g564(.A(G71gat), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n758_), .B2(new_n692_), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n767_), .B(KEYINPUT49), .Z(new_n768_));
  NAND3_X1  g567(.A1(new_n755_), .A2(new_n766_), .A3(new_n692_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(G1334gat));
  AOI21_X1  g569(.A(new_n620_), .B1(new_n758_), .B2(new_n296_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n771_), .B(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n755_), .A2(new_n620_), .A3(new_n296_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(G1335gat));
  NAND3_X1  g574(.A1(new_n753_), .A2(new_n664_), .A3(new_n702_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(G85gat), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n777_), .A2(new_n778_), .A3(new_n350_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n675_), .A2(new_n521_), .A3(new_n676_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n718_), .A2(new_n780_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n781_), .A2(new_n349_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n779_), .B1(new_n782_), .B2(new_n778_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT112), .ZN(G1336gat));
  OAI21_X1  g583(.A(G92gat), .B1(new_n781_), .B2(new_n473_), .ZN(new_n785_));
  OR3_X1    g584(.A1(new_n776_), .A2(G92gat), .A3(new_n473_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(G1337gat));
  NOR3_X1   g586(.A1(new_n776_), .A2(new_n389_), .A3(new_n562_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n718_), .A2(new_n692_), .A3(new_n780_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(new_n789_), .B2(G99gat), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT113), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT51), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n794_), .B1(new_n790_), .B2(KEYINPUT113), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n793_), .B1(new_n792_), .B2(new_n795_), .ZN(G1338gat));
  NAND3_X1  g595(.A1(new_n777_), .A2(new_n567_), .A3(new_n296_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n718_), .A2(new_n296_), .A3(new_n780_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n798_), .A2(new_n799_), .A3(G106gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n798_), .B2(G106gat), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g602(.A1(new_n296_), .A2(new_n442_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n804_), .A2(new_n388_), .A3(new_n350_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n805_), .A2(KEYINPUT59), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n508_), .A2(new_n503_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n503_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n498_), .A2(new_n501_), .A3(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n807_), .A2(new_n518_), .A3(new_n809_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n520_), .A2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n645_), .A2(new_n646_), .A3(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT118), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n588_), .A2(new_n625_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(new_n627_), .B2(new_n630_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n609_), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT12), .B1(new_n588_), .B2(new_n625_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n579_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n821_), .A2(new_n822_), .A3(new_n626_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n821_), .B2(new_n626_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n815_), .B(new_n818_), .C1(new_n823_), .C2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n641_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n631_), .A2(KEYINPUT55), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n821_), .A2(new_n822_), .A3(new_n626_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n815_), .B1(new_n829_), .B2(new_n818_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n814_), .B1(new_n826_), .B2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n818_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT118), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n833_), .A2(KEYINPUT119), .A3(new_n641_), .A4(new_n825_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT56), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n831_), .A2(new_n834_), .A3(KEYINPUT120), .A4(new_n835_), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n521_), .A2(KEYINPUT117), .A3(new_n642_), .ZN(new_n837_));
  AOI21_X1  g636(.A(KEYINPUT117), .B1(new_n521_), .B2(new_n642_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n836_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n831_), .A2(new_n835_), .A3(new_n834_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n826_), .A2(new_n830_), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT120), .B1(new_n842_), .B2(KEYINPUT56), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n813_), .B1(new_n840_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n702_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(KEYINPUT122), .B1(new_n845_), .B2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n836_), .A2(new_n839_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n833_), .A2(KEYINPUT56), .A3(new_n641_), .A4(new_n825_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n833_), .A2(new_n641_), .A3(new_n825_), .ZN(new_n854_));
  AOI21_X1  g653(.A(KEYINPUT56), .B1(new_n854_), .B2(new_n814_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n853_), .B1(new_n855_), .B2(new_n834_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n812_), .B1(new_n850_), .B2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n857_), .A2(new_n858_), .A3(new_n847_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n849_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT58), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n835_), .B1(new_n826_), .B2(new_n830_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n851_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n811_), .A2(new_n642_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n861_), .B1(new_n863_), .B2(new_n865_), .ZN(new_n866_));
  AOI211_X1 g665(.A(KEYINPUT58), .B(new_n864_), .C1(new_n862_), .C2(new_n851_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n606_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n857_), .A2(new_n673_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n870_), .B2(new_n846_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n676_), .B1(new_n860_), .B2(new_n871_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n675_), .A2(new_n716_), .A3(new_n522_), .A4(new_n676_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(KEYINPUT54), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT116), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n873_), .A2(KEYINPUT116), .A3(KEYINPUT54), .ZN(new_n877_));
  OAI21_X1  g676(.A(KEYINPUT115), .B1(new_n873_), .B2(KEYINPUT54), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT115), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n665_), .A2(new_n879_), .A3(new_n880_), .A4(new_n522_), .ZN(new_n881_));
  AOI22_X1  g680(.A1(new_n876_), .A2(new_n877_), .B1(new_n878_), .B2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n806_), .B1(new_n872_), .B2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n868_), .A2(new_n884_), .ZN(new_n885_));
  OAI211_X1 g684(.A(KEYINPUT121), .B(new_n606_), .C1(new_n866_), .C2(new_n867_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n846_), .B1(new_n845_), .B2(new_n702_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n844_), .A2(new_n836_), .A3(new_n839_), .ZN(new_n889_));
  AOI211_X1 g688(.A(KEYINPUT122), .B(new_n848_), .C1(new_n889_), .C2(new_n812_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n858_), .B1(new_n857_), .B2(new_n847_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n887_), .B(new_n888_), .C1(new_n890_), .C2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n664_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n876_), .A2(new_n877_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n878_), .A2(new_n881_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n805_), .B1(new_n893_), .B2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n521_), .B(new_n883_), .C1(new_n897_), .C2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(G113gat), .ZN(new_n900_));
  INV_X1    g699(.A(new_n805_), .ZN(new_n901_));
  AOI22_X1  g700(.A1(new_n846_), .A2(new_n870_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n676_), .B1(new_n902_), .B2(new_n860_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n901_), .B1(new_n903_), .B2(new_n882_), .ZN(new_n904_));
  OR3_X1    g703(.A1(new_n904_), .A2(G113gat), .A3(new_n522_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n900_), .A2(new_n905_), .ZN(G1340gat));
  OAI211_X1 g705(.A(new_n649_), .B(new_n883_), .C1(new_n897_), .C2(new_n898_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(KEYINPUT123), .B(G120gat), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n907_), .A2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n908_), .A2(KEYINPUT60), .ZN(new_n912_));
  OR2_X1    g711(.A1(new_n675_), .A2(KEYINPUT60), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n908_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n911_), .B1(new_n904_), .B2(new_n915_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n897_), .A2(KEYINPUT124), .A3(new_n914_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n910_), .A2(new_n918_), .ZN(G1341gat));
  AOI21_X1  g718(.A(G127gat), .B1(new_n897_), .B2(new_n676_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n872_), .A2(new_n882_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  AOI22_X1  g721(.A1(new_n922_), .A2(new_n806_), .B1(new_n904_), .B2(KEYINPUT59), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n664_), .A2(new_n306_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(KEYINPUT125), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n920_), .B1(new_n923_), .B2(new_n925_), .ZN(G1342gat));
  AOI21_X1  g725(.A(G134gat), .B1(new_n897_), .B2(new_n702_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n606_), .A2(G134gat), .ZN(new_n928_));
  XOR2_X1   g727(.A(new_n928_), .B(KEYINPUT126), .Z(new_n929_));
  AOI21_X1  g728(.A(new_n927_), .B1(new_n923_), .B2(new_n929_), .ZN(G1343gat));
  NAND2_X1  g729(.A1(new_n893_), .A2(new_n896_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n692_), .A2(new_n349_), .A3(new_n471_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n931_), .A2(new_n521_), .A3(new_n932_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g733(.A1(new_n931_), .A2(new_n649_), .A3(new_n932_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g735(.A1(new_n931_), .A2(new_n676_), .A3(new_n932_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(KEYINPUT61), .B(G155gat), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n937_), .B(new_n938_), .ZN(G1346gat));
  INV_X1    g738(.A(G162gat), .ZN(new_n940_));
  NAND4_X1  g739(.A1(new_n931_), .A2(new_n940_), .A3(new_n702_), .A4(new_n932_), .ZN(new_n941_));
  AND3_X1   g740(.A1(new_n931_), .A2(new_n606_), .A3(new_n932_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n941_), .B1(new_n942_), .B2(new_n940_), .ZN(G1347gat));
  NAND3_X1  g742(.A1(new_n692_), .A2(new_n349_), .A3(new_n442_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n944_), .A2(new_n296_), .ZN(new_n945_));
  OAI211_X1 g744(.A(new_n521_), .B(new_n945_), .C1(new_n872_), .C2(new_n882_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(G169gat), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(new_n948_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n946_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n950_));
  OAI211_X1 g749(.A(new_n949_), .B(new_n950_), .C1(new_n421_), .C2(new_n946_), .ZN(G1348gat));
  INV_X1    g750(.A(new_n945_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n921_), .A2(new_n952_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n953_), .A2(new_n649_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n903_), .A2(new_n882_), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n955_), .A2(new_n296_), .ZN(new_n956_));
  NOR3_X1   g755(.A1(new_n675_), .A2(new_n944_), .A3(new_n366_), .ZN(new_n957_));
  AOI22_X1  g756(.A1(new_n954_), .A2(new_n366_), .B1(new_n956_), .B2(new_n957_), .ZN(G1349gat));
  NOR2_X1   g757(.A1(new_n944_), .A2(new_n664_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n956_), .A2(new_n959_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(new_n664_), .A2(new_n363_), .ZN(new_n961_));
  AOI22_X1  g760(.A1(new_n960_), .A2(new_n361_), .B1(new_n953_), .B2(new_n961_), .ZN(G1350gat));
  NAND3_X1  g761(.A1(new_n953_), .A2(new_n359_), .A3(new_n702_), .ZN(new_n963_));
  NOR3_X1   g762(.A1(new_n921_), .A2(new_n716_), .A3(new_n952_), .ZN(new_n964_));
  OAI21_X1  g763(.A(new_n963_), .B1(new_n391_), .B2(new_n964_), .ZN(G1351gat));
  NOR4_X1   g764(.A1(new_n692_), .A2(new_n350_), .A3(new_n449_), .A4(new_n473_), .ZN(new_n966_));
  INV_X1    g765(.A(new_n966_), .ZN(new_n967_));
  NOR2_X1   g766(.A1(new_n955_), .A2(new_n967_), .ZN(new_n968_));
  AOI21_X1  g767(.A(G197gat), .B1(new_n968_), .B2(new_n521_), .ZN(new_n969_));
  NOR4_X1   g768(.A1(new_n955_), .A2(new_n245_), .A3(new_n522_), .A4(new_n967_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(new_n969_), .A2(new_n970_), .ZN(G1352gat));
  NAND3_X1  g770(.A1(new_n931_), .A2(new_n649_), .A3(new_n966_), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n972_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g772(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n974_));
  INV_X1    g773(.A(new_n974_), .ZN(new_n975_));
  AOI21_X1  g774(.A(new_n664_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n976_));
  AOI21_X1  g775(.A(new_n975_), .B1(new_n968_), .B2(new_n976_), .ZN(new_n977_));
  AND4_X1   g776(.A1(new_n931_), .A2(new_n966_), .A3(new_n975_), .A4(new_n976_), .ZN(new_n978_));
  NOR2_X1   g777(.A1(new_n977_), .A2(new_n978_), .ZN(G1354gat));
  NAND3_X1  g778(.A1(new_n968_), .A2(new_n238_), .A3(new_n702_), .ZN(new_n980_));
  NOR3_X1   g779(.A1(new_n955_), .A2(new_n716_), .A3(new_n967_), .ZN(new_n981_));
  OAI21_X1  g780(.A(new_n980_), .B1(new_n238_), .B2(new_n981_), .ZN(G1355gat));
endmodule


