//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n778_,
    new_n779_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n921_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_;
  INV_X1    g000(.A(KEYINPUT101), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G225gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT96), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT4), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n209_), .A2(new_n212_), .A3(new_n213_), .A4(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  OR2_X1    g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT84), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n219_), .B1(new_n216_), .B2(KEYINPUT1), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n216_), .A2(KEYINPUT1), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT1), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n222_), .A2(KEYINPUT84), .A3(G155gat), .A4(G162gat), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n220_), .A2(new_n221_), .A3(new_n217_), .A4(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(G141gat), .B(G148gat), .Z(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n218_), .A2(new_n226_), .ZN(new_n227_));
  OR2_X1    g026(.A1(G127gat), .A2(G134gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G127gat), .A2(G134gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G113gat), .B(G120gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT82), .ZN(new_n233_));
  OR2_X1    g032(.A1(G113gat), .A2(G120gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G113gat), .A2(G120gat), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n234_), .A2(new_n228_), .A3(new_n229_), .A4(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n232_), .A2(new_n233_), .A3(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n230_), .A2(new_n231_), .A3(KEYINPUT82), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n227_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n232_), .A2(new_n236_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n218_), .A2(new_n226_), .A3(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n206_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(KEYINPUT4), .B1(new_n227_), .B2(new_n239_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n205_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT97), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n240_), .A2(new_n246_), .A3(new_n203_), .A4(new_n242_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n240_), .A2(new_n203_), .A3(new_n242_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT97), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n245_), .A2(new_n247_), .A3(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT0), .B(G57gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(G85gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(G1gat), .B(G29gat), .Z(new_n253_));
  XOR2_X1   g052(.A(new_n252_), .B(new_n253_), .Z(new_n254_));
  NAND2_X1  g053(.A1(new_n250_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n254_), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n245_), .A2(new_n256_), .A3(new_n249_), .A4(new_n247_), .ZN(new_n257_));
  AND3_X1   g056(.A1(new_n255_), .A2(KEYINPUT100), .A3(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT100), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n250_), .A2(new_n259_), .A3(new_n254_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n202_), .B1(new_n258_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n260_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n255_), .A2(KEYINPUT100), .A3(new_n257_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n262_), .A2(KEYINPUT101), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n261_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(KEYINPUT79), .A2(KEYINPUT22), .ZN(new_n267_));
  INV_X1    g066(.A(G169gat), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n267_), .B1(new_n268_), .B2(KEYINPUT80), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT80), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n270_), .A2(KEYINPUT79), .A3(KEYINPUT22), .A4(G169gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT81), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT22), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(G169gat), .ZN(new_n275_));
  AOI21_X1  g074(.A(G176gat), .B1(new_n275_), .B2(KEYINPUT80), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n272_), .A2(new_n273_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT23), .ZN(new_n278_));
  INV_X1    g077(.A(G183gat), .ZN(new_n279_));
  INV_X1    g078(.A(G190gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n278_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n280_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n281_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n277_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n273_), .B1(new_n272_), .B2(new_n276_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT24), .ZN(new_n288_));
  INV_X1    g087(.A(G176gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(new_n268_), .A3(new_n289_), .ZN(new_n290_));
  AND3_X1   g089(.A1(new_n281_), .A2(new_n283_), .A3(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT25), .B(G183gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT78), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT26), .B1(new_n280_), .B2(KEYINPUT77), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT77), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT26), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n295_), .A2(new_n296_), .A3(G190gat), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n292_), .A2(new_n293_), .A3(new_n294_), .A4(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n268_), .A2(new_n289_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n299_), .A2(KEYINPUT24), .A3(new_n285_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n291_), .A2(new_n298_), .A3(new_n300_), .ZN(new_n301_));
  OR2_X1    g100(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n295_), .A2(G190gat), .ZN(new_n304_));
  AOI22_X1  g103(.A1(new_n302_), .A2(new_n303_), .B1(new_n304_), .B2(KEYINPUT26), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n293_), .B1(new_n305_), .B2(new_n297_), .ZN(new_n306_));
  OAI22_X1  g105(.A1(new_n286_), .A2(new_n287_), .B1(new_n301_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT30), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n307_), .A2(KEYINPUT30), .ZN(new_n310_));
  OR3_X1    g109(.A1(new_n309_), .A2(G43gat), .A3(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(G43gat), .B1(new_n309_), .B2(new_n310_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G227gat), .A2(G233gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(G15gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G71gat), .B(G99gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n314_), .B(new_n315_), .Z(new_n316_));
  NAND3_X1  g115(.A1(new_n311_), .A2(new_n312_), .A3(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n316_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT83), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n319_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT83), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n321_), .A2(new_n322_), .A3(new_n317_), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n239_), .B(KEYINPUT31), .Z(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n320_), .A2(new_n323_), .A3(new_n325_), .ZN(new_n326_));
  OAI211_X1 g125(.A(KEYINPUT83), .B(new_n324_), .C1(new_n318_), .C2(new_n319_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n266_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT85), .ZN(new_n330_));
  INV_X1    g129(.A(G204gat), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n330_), .B1(new_n331_), .B2(G197gat), .ZN(new_n332_));
  INV_X1    g131(.A(G197gat), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n333_), .A2(KEYINPUT85), .A3(G204gat), .ZN(new_n334_));
  AOI22_X1  g133(.A1(new_n332_), .A2(new_n334_), .B1(G197gat), .B2(new_n331_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT21), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n333_), .A2(G204gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n331_), .A2(G197gat), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n336_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(G211gat), .B(G218gat), .Z(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n337_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n332_), .A2(new_n334_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(new_n339_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT86), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT21), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n341_), .B1(new_n335_), .B2(KEYINPUT86), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n343_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n227_), .A2(KEYINPUT29), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(G50gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(G78gat), .B(G106gat), .Z(new_n354_));
  OR2_X1    g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n353_), .A2(new_n354_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n227_), .A2(KEYINPUT29), .ZN(new_n358_));
  XOR2_X1   g157(.A(new_n358_), .B(KEYINPUT28), .Z(new_n359_));
  NAND2_X1  g158(.A1(G228gat), .A2(G233gat), .ZN(new_n360_));
  INV_X1    g159(.A(G22gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n359_), .B(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n357_), .A2(new_n363_), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n359_), .A2(new_n362_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n359_), .A2(new_n362_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n355_), .A2(new_n365_), .A3(new_n366_), .A4(new_n356_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n364_), .A2(new_n367_), .ZN(new_n368_));
  XOR2_X1   g167(.A(G8gat), .B(G36gat), .Z(new_n369_));
  XNOR2_X1  g168(.A(G64gat), .B(G92gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n371_), .B(new_n372_), .Z(new_n373_));
  INV_X1    g172(.A(KEYINPUT92), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n281_), .A2(new_n283_), .A3(new_n290_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT90), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT26), .B(G190gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n292_), .A2(new_n378_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n379_), .A2(new_n300_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n285_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT22), .B(G169gat), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n381_), .B1(new_n382_), .B2(new_n289_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n284_), .A2(KEYINPUT91), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT91), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n281_), .A2(new_n385_), .A3(new_n282_), .A4(new_n283_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  AOI22_X1  g186(.A1(new_n377_), .A2(new_n380_), .B1(new_n383_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n341_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n389_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n336_), .B1(new_n335_), .B2(KEYINPUT86), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n390_), .A2(new_n391_), .B1(new_n342_), .B2(new_n337_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n374_), .B1(new_n388_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n291_), .A2(new_n376_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n375_), .A2(KEYINPUT90), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n380_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n387_), .A2(new_n383_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(KEYINPUT92), .A3(new_n349_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n393_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT88), .ZN(new_n402_));
  AND2_X1   g201(.A1(G226gat), .A2(G233gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n305_), .A2(new_n297_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT78), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n406_), .A2(new_n291_), .A3(new_n298_), .A4(new_n300_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n287_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n408_), .A2(new_n284_), .A3(new_n277_), .A4(new_n285_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n392_), .A2(new_n407_), .A3(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(KEYINPUT89), .B1(new_n410_), .B2(KEYINPUT20), .ZN(new_n411_));
  OAI211_X1 g210(.A(KEYINPUT89), .B(KEYINPUT20), .C1(new_n307_), .C2(new_n349_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n400_), .B(new_n404_), .C1(new_n411_), .C2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n307_), .A2(new_n349_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT94), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n388_), .A2(new_n392_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n307_), .A2(new_n349_), .A3(KEYINPUT94), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n417_), .A2(KEYINPUT20), .A3(new_n418_), .A4(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n404_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n373_), .B1(new_n414_), .B2(new_n422_), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n423_), .A2(KEYINPUT102), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT27), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n425_), .B1(new_n423_), .B2(KEYINPUT102), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT20), .B1(new_n307_), .B2(new_n349_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT89), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  AOI22_X1  g228(.A1(new_n429_), .A2(new_n412_), .B1(new_n393_), .B2(new_n399_), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT93), .B1(new_n430_), .B2(new_n404_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n400_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT93), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(new_n433_), .A3(new_n421_), .ZN(new_n434_));
  OR2_X1    g233(.A1(new_n420_), .A2(new_n421_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n431_), .A2(new_n434_), .A3(new_n373_), .A4(new_n435_), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n424_), .A2(new_n426_), .A3(new_n436_), .ZN(new_n437_));
  XOR2_X1   g236(.A(KEYINPUT103), .B(KEYINPUT27), .Z(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n431_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n373_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n439_), .B1(new_n442_), .B2(new_n436_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n437_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n329_), .A2(new_n368_), .A3(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n203_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n240_), .A2(new_n242_), .A3(new_n205_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(new_n254_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT33), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n449_), .B1(new_n257_), .B2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n257_), .A2(new_n450_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT98), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n257_), .A2(KEYINPUT98), .A3(new_n450_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n451_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n442_), .A2(new_n436_), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT99), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n373_), .A2(KEYINPUT32), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n431_), .A2(new_n434_), .A3(new_n460_), .A4(new_n435_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n414_), .A2(new_n422_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n462_), .A2(KEYINPUT32), .A3(new_n373_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n461_), .A2(new_n262_), .A3(new_n463_), .A4(new_n263_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n442_), .A2(new_n456_), .A3(KEYINPUT99), .A4(new_n436_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n459_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n368_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n442_), .A2(new_n436_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(new_n438_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n368_), .B1(new_n261_), .B2(new_n264_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n424_), .A2(new_n436_), .A3(new_n426_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n469_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT104), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT104), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n444_), .A2(new_n474_), .A3(new_n470_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n467_), .A2(new_n473_), .A3(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n446_), .B1(new_n476_), .B2(new_n328_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G15gat), .B(G22gat), .ZN(new_n478_));
  INV_X1    g277(.A(G1gat), .ZN(new_n479_));
  INV_X1    g278(.A(G8gat), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT14), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G1gat), .B(G8gat), .ZN(new_n483_));
  XOR2_X1   g282(.A(new_n482_), .B(new_n483_), .Z(new_n484_));
  NAND2_X1  g283(.A1(G231gat), .A2(G233gat), .ZN(new_n485_));
  XOR2_X1   g284(.A(new_n485_), .B(KEYINPUT74), .Z(new_n486_));
  XNOR2_X1  g285(.A(new_n484_), .B(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G57gat), .B(G64gat), .ZN(new_n488_));
  OR2_X1    g287(.A1(new_n488_), .A2(KEYINPUT11), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(KEYINPUT11), .ZN(new_n490_));
  XOR2_X1   g289(.A(G71gat), .B(G78gat), .Z(new_n491_));
  NAND3_X1  g290(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n490_), .A2(new_n491_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n487_), .B(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT17), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT16), .B(G183gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(G211gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G127gat), .B(G155gat), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n498_), .B(new_n499_), .Z(new_n500_));
  NOR3_X1   g299(.A1(new_n495_), .A2(new_n496_), .A3(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(KEYINPUT17), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n501_), .B1(new_n495_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(G99gat), .ZN(new_n505_));
  INV_X1    g304(.A(G106gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  OR2_X1    g306(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n508_));
  NAND2_X1  g307(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n507_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  OAI22_X1  g309(.A1(KEYINPUT65), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT66), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G99gat), .A2(G106gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT6), .ZN(new_n515_));
  NOR2_X1   g314(.A1(G99gat), .A2(G106gat), .ZN(new_n516_));
  AND2_X1   g315(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n517_));
  NOR2_X1   g316(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n516_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT66), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n519_), .A2(new_n520_), .A3(new_n511_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n513_), .A2(new_n515_), .A3(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(G85gat), .B(G92gat), .Z(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(KEYINPUT8), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT64), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT9), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n523_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  XOR2_X1   g328(.A(KEYINPUT10), .B(G99gat), .Z(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(new_n506_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n525_), .A2(new_n526_), .A3(G85gat), .A4(G92gat), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n529_), .A2(new_n531_), .A3(new_n532_), .A4(new_n515_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n515_), .A2(new_n519_), .A3(new_n511_), .ZN(new_n534_));
  AOI21_X1  g333(.A(KEYINPUT8), .B1(new_n534_), .B2(new_n523_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n524_), .A2(new_n533_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n494_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n524_), .A2(new_n533_), .A3(new_n536_), .A4(new_n494_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n539_), .A2(KEYINPUT12), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT12), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n537_), .A2(new_n542_), .A3(new_n538_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G230gat), .A2(G233gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n539_), .A2(new_n540_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n545_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT67), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT67), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n547_), .A2(new_n551_), .A3(new_n548_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n546_), .A2(new_n550_), .A3(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G120gat), .B(G148gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(new_n331_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT5), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(new_n289_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n553_), .A2(new_n558_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n546_), .A2(new_n550_), .A3(new_n552_), .A4(new_n557_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT13), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT13), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n559_), .A2(new_n563_), .A3(new_n560_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G229gat), .A2(G233gat), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT69), .B(G43gat), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n568_), .A2(new_n352_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n352_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(G29gat), .B(G36gat), .Z(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n572_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n574_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT75), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT75), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n578_), .A2(new_n484_), .A3(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n484_), .B1(new_n578_), .B2(new_n580_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n567_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n573_), .A2(KEYINPUT15), .A3(new_n575_), .ZN(new_n584_));
  AOI21_X1  g383(.A(KEYINPUT15), .B1(new_n573_), .B2(new_n575_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n484_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n578_), .A2(new_n484_), .A3(new_n580_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(new_n589_), .A3(new_n566_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n583_), .A2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G113gat), .B(G141gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(G197gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT76), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(new_n268_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n591_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n583_), .A2(new_n590_), .A3(new_n595_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n565_), .A2(new_n599_), .ZN(new_n600_));
  NOR3_X1   g399(.A1(new_n477_), .A2(new_n504_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT8), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n519_), .A2(new_n520_), .A3(new_n511_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n520_), .B1(new_n519_), .B2(new_n511_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n602_), .B1(new_n605_), .B2(new_n515_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n535_), .B1(new_n606_), .B2(new_n523_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n607_), .A2(KEYINPUT71), .A3(new_n533_), .A4(new_n576_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(G232gat), .A2(G233gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT34), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n610_), .A2(KEYINPUT35), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT71), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n612_), .B1(new_n537_), .B2(new_n577_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n608_), .A2(new_n611_), .A3(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT72), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n608_), .A2(new_n613_), .A3(KEYINPUT72), .A4(new_n611_), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n586_), .A2(KEYINPUT70), .A3(new_n537_), .ZN(new_n618_));
  AOI21_X1  g417(.A(KEYINPUT70), .B1(new_n586_), .B2(new_n537_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n616_), .A2(new_n617_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n610_), .A2(KEYINPUT35), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT68), .Z(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n586_), .A2(new_n537_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n614_), .A2(new_n623_), .A3(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n624_), .A2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G190gat), .B(G218gat), .ZN(new_n629_));
  INV_X1    g428(.A(G134gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(G162gat), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT36), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n632_), .A2(new_n633_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n628_), .A2(new_n634_), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT73), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n626_), .B1(new_n621_), .B2(new_n623_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n639_), .A2(new_n633_), .A3(new_n632_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n637_), .A2(new_n638_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT37), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n637_), .A2(new_n638_), .A3(KEYINPUT37), .A4(new_n640_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n601_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT38), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n266_), .A2(new_n479_), .ZN(new_n649_));
  OR3_X1    g448(.A1(new_n647_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n648_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n640_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n634_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n639_), .A2(new_n653_), .A3(new_n635_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n601_), .A2(new_n656_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n657_), .A2(new_n266_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n650_), .B(new_n651_), .C1(new_n479_), .C2(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT105), .ZN(G1324gat));
  INV_X1    g459(.A(new_n647_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n444_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n661_), .A2(new_n480_), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT39), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n657_), .A2(new_n662_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n664_), .B1(new_n665_), .B2(G8gat), .ZN(new_n666_));
  AOI211_X1 g465(.A(KEYINPUT39), .B(new_n480_), .C1(new_n657_), .C2(new_n662_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n663_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT40), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n668_), .B(new_n669_), .ZN(G1325gat));
  OR3_X1    g469(.A1(new_n647_), .A2(G15gat), .A3(new_n328_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n328_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n657_), .A2(new_n672_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n673_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(KEYINPUT41), .B1(new_n673_), .B2(G15gat), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n671_), .B1(new_n674_), .B2(new_n675_), .ZN(G1326gat));
  INV_X1    g475(.A(new_n368_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n661_), .A2(new_n361_), .A3(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT42), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n657_), .A2(new_n677_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n680_), .B2(G22gat), .ZN(new_n681_));
  AOI211_X1 g480(.A(KEYINPUT42), .B(new_n361_), .C1(new_n657_), .C2(new_n677_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n678_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT106), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n683_), .B(new_n684_), .ZN(G1327gat));
  NOR2_X1   g484(.A1(new_n600_), .A2(new_n503_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n477_), .A2(new_n656_), .A3(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(G29gat), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n688_), .A2(new_n689_), .A3(new_n266_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n476_), .A2(new_n328_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(new_n445_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n691_), .B1(new_n693_), .B2(new_n645_), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n477_), .A2(KEYINPUT43), .A3(new_n646_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n686_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(KEYINPUT107), .A3(KEYINPUT44), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n474_), .B1(new_n444_), .B2(new_n470_), .ZN(new_n699_));
  AND4_X1   g498(.A1(new_n474_), .A2(new_n469_), .A3(new_n470_), .A4(new_n471_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n672_), .B1(new_n701_), .B2(new_n467_), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n691_), .B(new_n645_), .C1(new_n702_), .C2(new_n446_), .ZN(new_n703_));
  OAI21_X1  g502(.A(KEYINPUT43), .B1(new_n477_), .B2(new_n646_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n687_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n698_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n265_), .B1(new_n697_), .B2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n690_), .B1(new_n708_), .B2(new_n689_), .ZN(G1328gat));
  INV_X1    g508(.A(G36gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n688_), .A2(new_n710_), .A3(new_n662_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT45), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n444_), .B1(new_n697_), .B2(new_n707_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(new_n710_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT46), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  OAI211_X1 g515(.A(KEYINPUT46), .B(new_n712_), .C1(new_n713_), .C2(new_n710_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1329gat));
  XNOR2_X1  g517(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT44), .B1(new_n696_), .B2(KEYINPUT107), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n705_), .A2(new_n706_), .A3(new_n698_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n672_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(G43gat), .ZN(new_n723_));
  INV_X1    g522(.A(G43gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n688_), .A2(new_n724_), .A3(new_n672_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n719_), .B1(new_n723_), .B2(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n328_), .B1(new_n697_), .B2(new_n707_), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n725_), .B(new_n719_), .C1(new_n727_), .C2(new_n724_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n726_), .A2(new_n729_), .ZN(G1330gat));
  NAND3_X1  g529(.A1(new_n688_), .A2(new_n352_), .A3(new_n677_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n368_), .B1(new_n697_), .B2(new_n707_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n732_), .B2(new_n352_), .ZN(G1331gat));
  NOR4_X1   g532(.A1(new_n477_), .A2(new_n504_), .A3(new_n599_), .A4(new_n565_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n734_), .A2(new_n656_), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n735_), .A2(G57gat), .A3(new_n266_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n646_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n737_), .B(new_n738_), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n739_), .A2(KEYINPUT110), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(KEYINPUT110), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n740_), .A2(new_n266_), .A3(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(G57gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n736_), .B1(new_n742_), .B2(new_n743_), .ZN(G1332gat));
  NOR2_X1   g543(.A1(new_n444_), .A2(G64gat), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT111), .Z(new_n746_));
  NAND2_X1  g545(.A1(new_n739_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n735_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G64gat), .B1(new_n748_), .B2(new_n444_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n749_), .A2(KEYINPUT48), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(KEYINPUT48), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n747_), .B1(new_n750_), .B2(new_n751_), .ZN(G1333gat));
  INV_X1    g551(.A(G71gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n739_), .A2(new_n753_), .A3(new_n672_), .ZN(new_n754_));
  OAI21_X1  g553(.A(G71gat), .B1(new_n748_), .B2(new_n328_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n755_), .A2(KEYINPUT49), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(KEYINPUT49), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n754_), .B1(new_n756_), .B2(new_n757_), .ZN(G1334gat));
  INV_X1    g557(.A(G78gat), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n739_), .A2(new_n759_), .A3(new_n677_), .ZN(new_n760_));
  OAI21_X1  g559(.A(G78gat), .B1(new_n748_), .B2(new_n368_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n761_), .A2(KEYINPUT50), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(KEYINPUT50), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n760_), .B1(new_n762_), .B2(new_n763_), .ZN(G1335gat));
  NOR3_X1   g563(.A1(new_n565_), .A2(new_n503_), .A3(new_n599_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n693_), .A2(new_n655_), .A3(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT112), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n693_), .A2(KEYINPUT112), .A3(new_n655_), .A4(new_n765_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(G85gat), .B1(new_n770_), .B2(new_n266_), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n694_), .A2(new_n695_), .A3(KEYINPUT113), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n773_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n774_));
  OR2_X1    g573(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n775_), .A2(G85gat), .A3(new_n765_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n771_), .B1(new_n776_), .B2(new_n266_), .ZN(G1336gat));
  AOI21_X1  g576(.A(G92gat), .B1(new_n770_), .B2(new_n662_), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n775_), .A2(new_n662_), .A3(new_n765_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(G92gat), .ZN(G1337gat));
  INV_X1    g579(.A(new_n530_), .ZN(new_n781_));
  AOI211_X1 g580(.A(new_n781_), .B(new_n328_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n672_), .B(new_n765_), .C1(new_n772_), .C2(new_n774_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n783_), .B2(G99gat), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT51), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n783_), .A2(G99gat), .ZN(new_n787_));
  INV_X1    g586(.A(new_n782_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n785_), .A3(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n784_), .B1(KEYINPUT114), .B2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n786_), .B1(new_n791_), .B2(new_n793_), .ZN(G1338gat));
  AOI21_X1  g593(.A(G106gat), .B1(new_n768_), .B2(new_n769_), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n795_), .A2(KEYINPUT116), .A3(new_n677_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT116), .B1(new_n795_), .B2(new_n677_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n677_), .B(new_n765_), .C1(new_n694_), .C2(new_n695_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n798_), .A2(new_n799_), .A3(G106gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n798_), .B2(G106gat), .ZN(new_n801_));
  OAI22_X1  g600(.A1(new_n796_), .A2(new_n797_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g602(.A1(new_n662_), .A2(new_n265_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n672_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT56), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n541_), .A2(new_n548_), .A3(new_n543_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n546_), .A2(KEYINPUT55), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n544_), .A2(new_n813_), .A3(new_n545_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n811_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n809_), .B1(new_n815_), .B2(new_n557_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n813_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n818_));
  AOI211_X1 g617(.A(KEYINPUT55), .B(new_n548_), .C1(new_n541_), .C2(new_n543_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n810_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n820_), .A2(KEYINPUT56), .A3(new_n558_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n816_), .A2(new_n817_), .A3(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n560_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT56), .B1(new_n820_), .B2(new_n558_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n823_), .B1(new_n824_), .B2(KEYINPUT117), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n822_), .A2(new_n825_), .A3(new_n599_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n566_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n588_), .A2(new_n589_), .A3(new_n567_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n827_), .A2(new_n828_), .A3(new_n596_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n598_), .A2(new_n829_), .ZN(new_n830_));
  AOI211_X1 g629(.A(KEYINPUT118), .B(new_n830_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n832_));
  INV_X1    g631(.A(new_n830_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(new_n561_), .B2(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n831_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n826_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n808_), .B1(new_n836_), .B2(new_n656_), .ZN(new_n837_));
  AOI211_X1 g636(.A(new_n655_), .B(new_n807_), .C1(new_n826_), .C2(new_n835_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n816_), .A2(new_n821_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n840_), .A2(new_n560_), .A3(new_n833_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n840_), .A2(KEYINPUT58), .A3(new_n560_), .A4(new_n833_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n645_), .A2(new_n843_), .A3(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n503_), .B1(new_n839_), .B2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n599_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n643_), .A2(new_n503_), .A3(new_n644_), .A4(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n848_), .B(new_n849_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n368_), .B(new_n806_), .C1(new_n846_), .C2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(G113gat), .B1(new_n852_), .B2(new_n599_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n599_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n851_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n836_), .A2(new_n656_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n807_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n836_), .A2(new_n656_), .A3(new_n808_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n858_), .A2(new_n859_), .A3(new_n845_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n504_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n850_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n863_), .A2(KEYINPUT59), .A3(new_n368_), .A4(new_n806_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n854_), .B1(new_n856_), .B2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n853_), .B1(new_n865_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g665(.A(G120gat), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n867_), .B1(new_n565_), .B2(KEYINPUT60), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n852_), .B(new_n868_), .C1(KEYINPUT60), .C2(new_n867_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n565_), .B1(new_n856_), .B2(new_n864_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n870_), .B2(new_n867_), .ZN(G1341gat));
  AOI21_X1  g670(.A(G127gat), .B1(new_n852_), .B2(new_n503_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(KEYINPUT120), .A2(G127gat), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n873_), .B1(new_n856_), .B2(new_n864_), .ZN(new_n874_));
  OAI21_X1  g673(.A(G127gat), .B1(new_n504_), .B2(KEYINPUT120), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n872_), .B1(new_n874_), .B2(new_n875_), .ZN(G1342gat));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n677_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n878_));
  AOI21_X1  g677(.A(KEYINPUT59), .B1(new_n878_), .B2(new_n806_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n850_), .B1(new_n860_), .B2(new_n504_), .ZN(new_n880_));
  NOR4_X1   g679(.A1(new_n880_), .A2(new_n855_), .A3(new_n677_), .A4(new_n805_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n645_), .B1(new_n879_), .B2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(G134gat), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n852_), .A2(new_n630_), .A3(new_n655_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n877_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n646_), .B1(new_n856_), .B2(new_n864_), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n877_), .B(new_n884_), .C1(new_n886_), .C2(new_n630_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n885_), .A2(new_n888_), .ZN(G1343gat));
  NAND3_X1  g688(.A1(new_n804_), .A2(new_n328_), .A3(new_n677_), .ZN(new_n890_));
  XOR2_X1   g689(.A(new_n890_), .B(KEYINPUT122), .Z(new_n891_));
  NAND2_X1  g690(.A1(new_n863_), .A2(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n854_), .ZN(new_n893_));
  XOR2_X1   g692(.A(KEYINPUT123), .B(G141gat), .Z(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1344gat));
  NOR2_X1   g694(.A1(new_n892_), .A2(new_n565_), .ZN(new_n896_));
  XOR2_X1   g695(.A(new_n896_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g696(.A1(new_n892_), .A2(new_n504_), .ZN(new_n898_));
  XOR2_X1   g697(.A(KEYINPUT61), .B(G155gat), .Z(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(G1346gat));
  INV_X1    g699(.A(new_n892_), .ZN(new_n901_));
  AOI21_X1  g700(.A(G162gat), .B1(new_n901_), .B2(new_n655_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n645_), .A2(G162gat), .ZN(new_n903_));
  XOR2_X1   g702(.A(new_n903_), .B(KEYINPUT124), .Z(new_n904_));
  AOI21_X1  g703(.A(new_n902_), .B1(new_n901_), .B2(new_n904_), .ZN(G1347gat));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n878_), .A2(new_n662_), .A3(new_n329_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n854_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n906_), .B1(new_n908_), .B2(new_n268_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n382_), .ZN(new_n910_));
  OAI211_X1 g709(.A(KEYINPUT62), .B(G169gat), .C1(new_n907_), .C2(new_n854_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n909_), .A2(new_n910_), .A3(new_n911_), .ZN(G1348gat));
  NOR2_X1   g711(.A1(new_n907_), .A2(new_n565_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(new_n289_), .ZN(G1349gat));
  NOR2_X1   g713(.A1(new_n907_), .A2(new_n504_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n292_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n916_), .B1(new_n279_), .B2(new_n915_), .ZN(G1350gat));
  OAI21_X1  g716(.A(G190gat), .B1(new_n907_), .B2(new_n646_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n655_), .A2(new_n378_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n907_), .B2(new_n919_), .ZN(G1351gat));
  NAND4_X1  g719(.A1(new_n863_), .A2(new_n328_), .A3(new_n470_), .A4(new_n662_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n921_), .A2(new_n854_), .ZN(new_n922_));
  XOR2_X1   g721(.A(KEYINPUT125), .B(G197gat), .Z(new_n923_));
  XNOR2_X1  g722(.A(new_n922_), .B(new_n923_), .ZN(G1352gat));
  NOR2_X1   g723(.A1(new_n921_), .A2(new_n565_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n925_), .B(new_n926_), .ZN(G1353gat));
  NOR2_X1   g726(.A1(new_n921_), .A2(new_n504_), .ZN(new_n928_));
  NOR3_X1   g727(.A1(new_n928_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n929_));
  XOR2_X1   g728(.A(KEYINPUT63), .B(G211gat), .Z(new_n930_));
  AOI21_X1  g729(.A(new_n929_), .B1(new_n928_), .B2(new_n930_), .ZN(G1354gat));
  NOR2_X1   g730(.A1(new_n921_), .A2(new_n656_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n932_), .A2(G218gat), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n921_), .A2(new_n646_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n933_), .B1(G218gat), .B2(new_n934_), .ZN(G1355gat));
endmodule


