//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 0 0 1 1 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n883_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n919_, new_n920_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n941_;
  INV_X1    g000(.A(KEYINPUT20), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT26), .B(G190gat), .Z(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT77), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT78), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT77), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT26), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n206_), .B1(new_n207_), .B2(G190gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT25), .B(G183gat), .ZN(new_n209_));
  NAND4_X1  g008(.A1(new_n204_), .A2(new_n205_), .A3(new_n208_), .A4(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT26), .B(G190gat), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n208_), .B(new_n209_), .C1(new_n211_), .C2(new_n206_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT78), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G169gat), .B(G176gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT24), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G183gat), .ZN(new_n218_));
  INV_X1    g017(.A(G190gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT23), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G183gat), .A3(G190gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(new_n216_), .ZN(new_n225_));
  AND3_X1   g024(.A1(new_n217_), .A2(new_n223_), .A3(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n222_), .A2(KEYINPUT79), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(new_n220_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n218_), .A2(new_n219_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(G169gat), .ZN(new_n232_));
  AOI22_X1  g031(.A1(new_n214_), .A2(new_n226_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(G197gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(G204gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT87), .ZN(new_n236_));
  INV_X1    g035(.A(G204gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(G197gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT87), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n239_), .A2(new_n234_), .A3(G204gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n236_), .A2(new_n238_), .A3(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT89), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G211gat), .B(G218gat), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT21), .B1(new_n244_), .B2(KEYINPUT88), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n245_), .B1(KEYINPUT88), .B2(new_n244_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n241_), .A2(KEYINPUT21), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n235_), .A2(new_n238_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT21), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n249_), .A2(new_n244_), .ZN(new_n250_));
  AOI22_X1  g049(.A1(new_n243_), .A2(new_n246_), .B1(new_n247_), .B2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n202_), .B1(new_n233_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT92), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n209_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT25), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n255_), .A2(G183gat), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n218_), .A2(KEYINPUT25), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT92), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n254_), .A2(new_n258_), .A3(new_n211_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT93), .B(KEYINPUT24), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n215_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT94), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT94), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n259_), .A2(new_n264_), .A3(new_n261_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n260_), .A2(new_n224_), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n228_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n223_), .A2(new_n229_), .ZN(new_n269_));
  AOI22_X1  g068(.A1(new_n266_), .A2(new_n268_), .B1(new_n232_), .B2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n252_), .B1(new_n270_), .B2(new_n251_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G226gat), .A2(G233gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT19), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n273_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n270_), .A2(new_n251_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n214_), .A2(new_n226_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n230_), .A2(new_n232_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n243_), .A2(new_n246_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n247_), .A2(new_n250_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n202_), .B1(new_n279_), .B2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n275_), .B1(new_n276_), .B2(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n274_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G8gat), .B(G36gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT18), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G64gat), .B(G92gat), .ZN(new_n288_));
  XOR2_X1   g087(.A(new_n287_), .B(new_n288_), .Z(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT27), .B1(new_n285_), .B2(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT20), .B1(new_n279_), .B2(new_n282_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n265_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n264_), .B1(new_n259_), .B2(new_n261_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n268_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n269_), .A2(new_n232_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n251_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n273_), .B1(new_n291_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT95), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n276_), .A2(new_n275_), .A3(new_n283_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT95), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n300_), .B(new_n273_), .C1(new_n291_), .C2(new_n296_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n298_), .A2(new_n299_), .A3(new_n301_), .A4(new_n289_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n290_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n289_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n301_), .A2(new_n299_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n300_), .B1(new_n271_), .B2(new_n273_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n305_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n302_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT27), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT101), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT101), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n309_), .A2(new_n313_), .A3(new_n310_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n304_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(G22gat), .B(G50gat), .Z(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(G155gat), .ZN(new_n321_));
  INV_X1    g120(.A(G162gat), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n321_), .A2(new_n322_), .A3(KEYINPUT81), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT81), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n324_), .B1(G155gat), .B2(G162gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n323_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n327_), .A2(KEYINPUT84), .ZN(new_n328_));
  OR3_X1    g127(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT2), .ZN(new_n330_));
  INV_X1    g129(.A(G141gat), .ZN(new_n331_));
  INV_X1    g130(.A(G148gat), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n330_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n329_), .A2(new_n333_), .A3(new_n334_), .A4(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n327_), .A2(KEYINPUT84), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n328_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n326_), .A2(KEYINPUT1), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n323_), .A2(new_n339_), .A3(new_n325_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT82), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n326_), .A2(KEYINPUT1), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n323_), .A2(new_n339_), .A3(new_n325_), .A4(KEYINPUT82), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  XOR2_X1   g144(.A(G141gat), .B(G148gat), .Z(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(KEYINPUT83), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT83), .B1(new_n345_), .B2(new_n346_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n338_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT85), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n338_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n345_), .A2(new_n346_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT83), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n353_), .B1(new_n356_), .B2(new_n347_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT85), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n352_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT29), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n320_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  AOI211_X1 g160(.A(KEYINPUT29), .B(new_n319_), .C1(new_n352_), .C2(new_n358_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n318_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n357_), .A2(KEYINPUT85), .ZN(new_n364_));
  AOI211_X1 g163(.A(new_n351_), .B(new_n353_), .C1(new_n356_), .C2(new_n347_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n360_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(new_n319_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n359_), .A2(new_n360_), .A3(new_n320_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n367_), .A2(new_n317_), .A3(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G78gat), .B(G106gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT90), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n363_), .A2(new_n369_), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT91), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n251_), .B1(G228gat), .B2(G233gat), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n376_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n282_), .B1(new_n357_), .B2(new_n360_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n378_), .A2(G228gat), .A3(G233gat), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n375_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n377_), .A2(new_n375_), .A3(new_n379_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n372_), .B1(new_n363_), .B2(new_n369_), .ZN(new_n384_));
  NOR3_X1   g183(.A1(new_n374_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n382_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n386_), .A2(new_n380_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n363_), .A2(new_n369_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n371_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n387_), .B1(new_n389_), .B2(new_n373_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n385_), .A2(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(G1gat), .B(G29gat), .Z(new_n392_));
  XNOR2_X1  g191(.A(G57gat), .B(G85gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  XOR2_X1   g193(.A(KEYINPUT97), .B(KEYINPUT0), .Z(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G127gat), .B(G134gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G113gat), .B(G120gat), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n398_), .B(new_n399_), .Z(new_n400_));
  NAND3_X1  g199(.A1(new_n352_), .A2(new_n358_), .A3(new_n400_), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n350_), .A2(new_n400_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(KEYINPUT4), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G225gat), .A2(G233gat), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  XOR2_X1   g204(.A(KEYINPUT96), .B(KEYINPUT4), .Z(new_n406_));
  NAND4_X1  g205(.A1(new_n352_), .A2(new_n358_), .A3(new_n400_), .A4(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n403_), .A2(new_n405_), .A3(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n401_), .A2(new_n402_), .A3(new_n404_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n397_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT99), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n403_), .A2(new_n405_), .A3(new_n407_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n409_), .A2(new_n397_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n411_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n413_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(KEYINPUT99), .A3(new_n408_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n410_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G227gat), .A2(G233gat), .ZN(new_n418_));
  INV_X1    g217(.A(G71gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(G99gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n233_), .B(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(new_n400_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G15gat), .B(G43gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT80), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT30), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT31), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n424_), .B(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n417_), .A2(new_n429_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n316_), .A2(new_n391_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT100), .ZN(new_n432_));
  NOR3_X1   g231(.A1(new_n412_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT99), .B1(new_n415_), .B2(new_n408_), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n408_), .A2(new_n409_), .ZN(new_n435_));
  OAI22_X1  g234(.A1(new_n433_), .A2(new_n434_), .B1(new_n435_), .B2(new_n397_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n289_), .A2(KEYINPUT32), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n285_), .A2(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n306_), .A2(new_n307_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n438_), .B1(new_n439_), .B2(new_n437_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT33), .ZN(new_n441_));
  NOR3_X1   g240(.A1(new_n412_), .A2(new_n441_), .A3(new_n413_), .ZN(new_n442_));
  AOI21_X1  g241(.A(KEYINPUT33), .B1(new_n415_), .B2(new_n408_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n401_), .A2(KEYINPUT98), .A3(new_n402_), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT98), .B1(new_n401_), .B2(new_n402_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n405_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n407_), .A2(new_n404_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n397_), .B1(new_n448_), .B2(new_n403_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n309_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n436_), .A2(new_n440_), .B1(new_n444_), .B2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n432_), .B1(new_n451_), .B2(new_n391_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n309_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n441_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n449_), .A2(new_n447_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n415_), .A2(KEYINPUT33), .A3(new_n408_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n453_), .A2(new_n454_), .A3(new_n455_), .A4(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n440_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n457_), .B1(new_n417_), .B2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n383_), .B1(new_n374_), .B2(new_n384_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n389_), .A2(new_n387_), .A3(new_n373_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n459_), .A2(KEYINPUT100), .A3(new_n462_), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n460_), .A2(new_n417_), .A3(new_n461_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(new_n315_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n452_), .A2(new_n463_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n429_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n431_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G29gat), .B(G36gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G43gat), .B(G50gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT15), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G1gat), .B(G8gat), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n473_), .A2(KEYINPUT73), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(KEYINPUT73), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G15gat), .B(G22gat), .ZN(new_n477_));
  INV_X1    g276(.A(G1gat), .ZN(new_n478_));
  INV_X1    g277(.A(G8gat), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT14), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n476_), .B(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n472_), .A2(new_n482_), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n483_), .A2(KEYINPUT74), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G229gat), .A2(G233gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT75), .ZN(new_n486_));
  INV_X1    g285(.A(new_n471_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n482_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n483_), .A2(KEYINPUT74), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n484_), .A2(new_n486_), .A3(new_n488_), .A4(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT76), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n489_), .A2(new_n488_), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n493_), .A2(new_n484_), .A3(KEYINPUT76), .A4(new_n486_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n482_), .B(new_n487_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n495_), .A2(G229gat), .A3(G233gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n492_), .A2(new_n494_), .A3(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G113gat), .B(G141gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G169gat), .B(G197gat), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n498_), .B(new_n499_), .Z(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n497_), .A2(new_n501_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n492_), .A2(new_n494_), .A3(new_n496_), .A4(new_n500_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n468_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G232gat), .A2(G233gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT34), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT70), .B(KEYINPUT35), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(G106gat), .ZN(new_n512_));
  AND2_X1   g311(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n513_));
  NOR2_X1   g312(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n514_));
  NOR3_X1   g313(.A1(new_n513_), .A2(new_n514_), .A3(KEYINPUT64), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT64), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT10), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(new_n421_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n516_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n512_), .B1(new_n515_), .B2(new_n520_), .ZN(new_n521_));
  AND2_X1   g320(.A1(G85gat), .A2(G92gat), .ZN(new_n522_));
  NOR2_X1   g321(.A1(G85gat), .A2(G92gat), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT9), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(G92gat), .ZN(new_n525_));
  INV_X1    g324(.A(G85gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT65), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT65), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(G85gat), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n525_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n524_), .B1(new_n530_), .B2(KEYINPUT9), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G99gat), .A2(G106gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT6), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT6), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n534_), .A2(G99gat), .A3(G106gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n521_), .A2(new_n531_), .A3(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT7), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n539_), .A2(new_n421_), .A3(new_n512_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n536_), .A2(new_n538_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT8), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n522_), .A2(new_n523_), .A3(KEYINPUT66), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n542_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n537_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n511_), .B1(new_n546_), .B2(new_n487_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n547_), .B1(new_n472_), .B2(new_n546_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n509_), .A2(new_n510_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(G190gat), .B(G218gat), .Z(new_n551_));
  XNOR2_X1  g350(.A(G134gat), .B(G162gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT36), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n555_), .B(KEYINPUT71), .Z(new_n556_));
  NAND2_X1  g355(.A1(new_n550_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT37), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n553_), .B(KEYINPUT36), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n550_), .A2(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n558_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n550_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT72), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n560_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n565_), .B1(new_n564_), .B2(new_n563_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(new_n557_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT37), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n562_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G231gat), .A2(G233gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n482_), .B(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n573_), .A2(new_n574_), .A3(G78gat), .ZN(new_n575_));
  INV_X1    g374(.A(G64gat), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(G57gat), .ZN(new_n577_));
  INV_X1    g376(.A(G57gat), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(G64gat), .ZN(new_n579_));
  AOI21_X1  g378(.A(KEYINPUT11), .B1(new_n577_), .B2(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n575_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n577_), .A2(new_n579_), .A3(KEYINPUT11), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT68), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G57gat), .B(G64gat), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT68), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(new_n585_), .A3(KEYINPUT11), .ZN(new_n586_));
  OAI21_X1  g385(.A(G78gat), .B1(new_n573_), .B2(new_n574_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n581_), .A2(new_n583_), .A3(new_n586_), .A4(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n583_), .A2(new_n586_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n574_), .ZN(new_n590_));
  INV_X1    g389(.A(G78gat), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n590_), .A2(new_n591_), .A3(new_n572_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n592_), .B(new_n587_), .C1(KEYINPUT11), .C2(new_n584_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n589_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n588_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n571_), .B(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(G127gat), .B(G155gat), .Z(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT16), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G183gat), .B(G211gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT17), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n601_), .A2(new_n602_), .ZN(new_n604_));
  OR3_X1    g403(.A1(new_n597_), .A2(new_n603_), .A3(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n597_), .A2(new_n603_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n569_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT12), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n533_), .A2(new_n535_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n540_), .A2(new_n538_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n543_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(KEYINPUT8), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n615_));
  OAI21_X1  g414(.A(KEYINPUT64), .B1(new_n513_), .B2(new_n514_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n518_), .A2(new_n516_), .A3(new_n519_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n611_), .B1(new_n618_), .B2(new_n512_), .ZN(new_n619_));
  AOI22_X1  g418(.A1(new_n614_), .A2(new_n615_), .B1(new_n619_), .B2(new_n531_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n610_), .B1(new_n620_), .B2(new_n595_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n588_), .A2(new_n594_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n622_), .A2(new_n546_), .A3(KEYINPUT12), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n614_), .A2(new_n615_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n595_), .A2(new_n625_), .A3(new_n537_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(G230gat), .A2(G233gat), .ZN(new_n627_));
  AOI21_X1  g426(.A(KEYINPUT69), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT69), .ZN(new_n629_));
  INV_X1    g428(.A(new_n627_), .ZN(new_n630_));
  AOI211_X1 g429(.A(new_n629_), .B(new_n630_), .C1(new_n620_), .C2(new_n595_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n624_), .B1(new_n628_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n626_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n620_), .A2(new_n595_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n630_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n632_), .A2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(G120gat), .B(G148gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT5), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G176gat), .B(G204gat), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n638_), .B(new_n639_), .Z(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n636_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n636_), .A2(new_n641_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT13), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n642_), .A2(KEYINPUT13), .A3(new_n643_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n609_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n506_), .A2(new_n649_), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n650_), .A2(G1gat), .A3(new_n417_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n651_), .A2(KEYINPUT38), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT104), .ZN(new_n653_));
  INV_X1    g452(.A(new_n567_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n468_), .A2(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n648_), .A2(new_n505_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(new_n608_), .A3(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G1gat), .B1(new_n657_), .B2(new_n417_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT103), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n651_), .A2(KEYINPUT38), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT102), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n660_), .B(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n653_), .A2(new_n659_), .A3(new_n662_), .ZN(G1324gat));
  NOR3_X1   g462(.A1(new_n650_), .A2(G8gat), .A3(new_n315_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G8gat), .B1(new_n657_), .B2(new_n315_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT39), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT39), .ZN(new_n667_));
  OAI211_X1 g466(.A(new_n667_), .B(G8gat), .C1(new_n657_), .C2(new_n315_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n664_), .B1(new_n666_), .B2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n669_), .B(new_n671_), .ZN(G1325gat));
  OR3_X1    g471(.A1(new_n650_), .A2(G15gat), .A3(new_n467_), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n657_), .A2(new_n467_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n674_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(KEYINPUT41), .B1(new_n674_), .B2(G15gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n673_), .B1(new_n675_), .B2(new_n676_), .ZN(G1326gat));
  XNOR2_X1  g476(.A(new_n462_), .B(KEYINPUT106), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  OR3_X1    g478(.A1(new_n650_), .A2(G22gat), .A3(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G22gat), .B1(new_n657_), .B2(new_n679_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n681_), .A2(KEYINPUT42), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(KEYINPUT42), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n680_), .B1(new_n682_), .B2(new_n683_), .ZN(G1327gat));
  OAI21_X1  g483(.A(KEYINPUT43), .B1(new_n468_), .B2(new_n569_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n686_));
  INV_X1    g485(.A(new_n569_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n459_), .A2(new_n462_), .ZN(new_n688_));
  AOI22_X1  g487(.A1(new_n688_), .A2(new_n432_), .B1(new_n464_), .B2(new_n315_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n429_), .B1(new_n689_), .B2(new_n463_), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n686_), .B(new_n687_), .C1(new_n690_), .C2(new_n431_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n685_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n656_), .A2(new_n607_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(KEYINPUT44), .B1(new_n692_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696_));
  AOI211_X1 g495(.A(new_n696_), .B(new_n693_), .C1(new_n685_), .C2(new_n691_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n695_), .A2(new_n697_), .A3(new_n417_), .ZN(new_n698_));
  INV_X1    g497(.A(G29gat), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n567_), .A2(new_n608_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n701_), .A2(new_n648_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n506_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n436_), .A2(new_n699_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT107), .ZN(new_n705_));
  OAI22_X1  g504(.A1(new_n698_), .A2(new_n699_), .B1(new_n703_), .B2(new_n705_), .ZN(G1328gat));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707_));
  INV_X1    g506(.A(G36gat), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n695_), .A2(new_n697_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n709_), .B2(new_n316_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n315_), .A2(G36gat), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  OR3_X1    g511(.A1(new_n703_), .A2(KEYINPUT45), .A3(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(KEYINPUT45), .B1(new_n703_), .B2(new_n712_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n707_), .B1(new_n710_), .B2(new_n716_), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n695_), .A2(new_n697_), .A3(new_n315_), .ZN(new_n718_));
  OAI211_X1 g517(.A(KEYINPUT46), .B(new_n715_), .C1(new_n718_), .C2(new_n708_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(G1329gat));
  NAND2_X1  g519(.A1(new_n429_), .A2(G43gat), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n695_), .A2(new_n697_), .A3(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n703_), .ZN(new_n723_));
  AOI21_X1  g522(.A(G43gat), .B1(new_n723_), .B2(new_n429_), .ZN(new_n724_));
  OR3_X1    g523(.A1(new_n722_), .A2(KEYINPUT47), .A3(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(KEYINPUT47), .B1(new_n722_), .B2(new_n724_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1330gat));
  AOI21_X1  g526(.A(G50gat), .B1(new_n723_), .B2(new_n678_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n391_), .A2(G50gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n709_), .B2(new_n729_), .ZN(G1331gat));
  INV_X1    g529(.A(new_n648_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n609_), .A2(new_n731_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT108), .Z(new_n733_));
  NOR3_X1   g532(.A1(new_n733_), .A2(new_n468_), .A3(new_n504_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(new_n578_), .A3(new_n436_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n731_), .A2(new_n504_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n655_), .A2(new_n608_), .A3(new_n736_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n737_), .A2(new_n436_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n735_), .B1(new_n738_), .B2(new_n578_), .ZN(G1332gat));
  AOI21_X1  g538(.A(new_n576_), .B1(new_n737_), .B2(new_n316_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT48), .Z(new_n741_));
  NAND3_X1  g540(.A1(new_n734_), .A2(new_n576_), .A3(new_n316_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1333gat));
  AOI21_X1  g542(.A(new_n419_), .B1(new_n737_), .B2(new_n429_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT49), .Z(new_n745_));
  NAND3_X1  g544(.A1(new_n734_), .A2(new_n419_), .A3(new_n429_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1334gat));
  AOI21_X1  g546(.A(new_n591_), .B1(new_n737_), .B2(new_n678_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT50), .Z(new_n749_));
  NAND3_X1  g548(.A1(new_n734_), .A2(new_n591_), .A3(new_n678_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1335gat));
  INV_X1    g550(.A(new_n468_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n752_), .A2(new_n505_), .A3(new_n648_), .A4(new_n700_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(G85gat), .B1(new_n754_), .B2(new_n436_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n736_), .A2(new_n607_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n685_), .B2(new_n691_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT109), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n417_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(G1336gat));
  NAND3_X1  g559(.A1(new_n754_), .A2(new_n525_), .A3(new_n316_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n758_), .A2(new_n316_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n761_), .B1(new_n762_), .B2(new_n525_), .ZN(G1337gat));
  NAND3_X1  g562(.A1(new_n754_), .A2(new_n429_), .A3(new_n618_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n757_), .A2(new_n429_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(new_n421_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n766_), .B(new_n767_), .Z(G1338gat));
  NAND3_X1  g567(.A1(new_n754_), .A2(new_n512_), .A3(new_n391_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n757_), .A2(new_n391_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(G106gat), .ZN(new_n772_));
  AOI211_X1 g571(.A(KEYINPUT52), .B(new_n512_), .C1(new_n757_), .C2(new_n391_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT53), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT53), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n776_), .B(new_n769_), .C1(new_n772_), .C2(new_n773_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(G1339gat));
  NAND4_X1  g577(.A1(new_n315_), .A2(new_n462_), .A3(new_n436_), .A4(new_n429_), .ZN(new_n779_));
  XOR2_X1   g578(.A(new_n779_), .B(KEYINPUT115), .Z(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n500_), .B1(new_n495_), .B2(new_n486_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n493_), .A2(new_n484_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n782_), .B1(new_n783_), .B2(new_n486_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n503_), .A2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n785_), .B1(new_n643_), .B2(new_n642_), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n502_), .A2(new_n503_), .B1(new_n636_), .B2(new_n641_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n621_), .A2(new_n623_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n630_), .B1(new_n788_), .B2(new_n633_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n627_), .B1(new_n622_), .B2(new_n546_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n629_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n626_), .A2(KEYINPUT69), .A3(new_n627_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n788_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(KEYINPUT111), .B(KEYINPUT55), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n789_), .B1(new_n793_), .B2(new_n795_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n624_), .B(KEYINPUT55), .C1(new_n628_), .C2(new_n631_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(KEYINPUT112), .B1(new_n796_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n632_), .A2(new_n794_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT112), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n800_), .A2(new_n801_), .A3(new_n797_), .A4(new_n789_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n799_), .A2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT56), .B1(new_n803_), .B2(new_n640_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT56), .ZN(new_n805_));
  AOI211_X1 g604(.A(new_n805_), .B(new_n641_), .C1(new_n799_), .C2(new_n802_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n787_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n786_), .B1(new_n807_), .B2(KEYINPUT113), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n809_), .B(new_n787_), .C1(new_n804_), .C2(new_n806_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n654_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n785_), .B1(new_n636_), .B2(new_n641_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n812_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT58), .ZN(new_n814_));
  OR2_X1    g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n569_), .B1(new_n814_), .B2(new_n813_), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n811_), .A2(KEYINPUT57), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n807_), .A2(KEYINPUT113), .ZN(new_n818_));
  INV_X1    g617(.A(new_n786_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n810_), .A3(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n567_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT57), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n821_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(KEYINPUT114), .B1(new_n811_), .B2(KEYINPUT57), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n817_), .A2(new_n824_), .A3(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n607_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n828_), .B1(new_n649_), .B2(new_n505_), .ZN(new_n829_));
  NOR4_X1   g628(.A1(new_n609_), .A2(KEYINPUT54), .A3(new_n504_), .A4(new_n648_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n781_), .B1(new_n827_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n821_), .A2(new_n823_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n608_), .B1(new_n817_), .B2(new_n835_), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n836_), .A2(new_n831_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n781_), .A2(KEYINPUT59), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n834_), .A2(KEYINPUT59), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n504_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(G113gat), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n827_), .A2(new_n832_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT116), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n843_), .A3(new_n780_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n831_), .B1(new_n826_), .B2(new_n607_), .ZN(new_n845_));
  OAI21_X1  g644(.A(KEYINPUT116), .B1(new_n845_), .B2(new_n781_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n505_), .A2(G113gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n844_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n841_), .A2(new_n848_), .ZN(G1340gat));
  OAI21_X1  g648(.A(new_n838_), .B1(new_n831_), .B2(new_n836_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT59), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n648_), .B(new_n850_), .C1(new_n833_), .C2(new_n851_), .ZN(new_n852_));
  XOR2_X1   g651(.A(KEYINPUT117), .B(G120gat), .Z(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n854_), .ZN(new_n855_));
  OR2_X1    g654(.A1(new_n853_), .A2(KEYINPUT60), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n853_), .B1(new_n731_), .B2(KEYINPUT60), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n844_), .A2(new_n846_), .A3(new_n856_), .A4(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n855_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(KEYINPUT118), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n855_), .A2(new_n861_), .A3(new_n858_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(G1341gat));
  INV_X1    g662(.A(G127gat), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n607_), .A2(new_n864_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(KEYINPUT119), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n844_), .A2(new_n608_), .A3(new_n846_), .ZN(new_n867_));
  AOI22_X1  g666(.A1(new_n839_), .A2(new_n866_), .B1(new_n867_), .B2(new_n864_), .ZN(G1342gat));
  OAI211_X1 g667(.A(new_n687_), .B(new_n850_), .C1(new_n833_), .C2(new_n851_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(G134gat), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n567_), .A2(G134gat), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n844_), .A2(new_n846_), .A3(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT120), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n870_), .A2(KEYINPUT120), .A3(new_n872_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1343gat));
  NOR4_X1   g676(.A1(new_n316_), .A2(new_n462_), .A3(new_n417_), .A4(new_n429_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n842_), .A2(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(new_n505_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(KEYINPUT121), .B(G141gat), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n880_), .B(new_n881_), .ZN(G1344gat));
  NOR2_X1   g681(.A1(new_n879_), .A2(new_n731_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(new_n332_), .ZN(G1345gat));
  INV_X1    g683(.A(new_n879_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n885_), .A2(new_n886_), .A3(new_n608_), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT122), .B1(new_n879_), .B2(new_n607_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT61), .B(G155gat), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n887_), .A2(new_n888_), .A3(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1346gat));
  OAI21_X1  g691(.A(G162gat), .B1(new_n879_), .B2(new_n569_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n654_), .A2(new_n322_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n879_), .B2(new_n894_), .ZN(G1347gat));
  NOR3_X1   g694(.A1(new_n678_), .A2(new_n315_), .A3(new_n430_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n837_), .A2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n504_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n900_), .A2(KEYINPUT62), .ZN(new_n901_));
  INV_X1    g700(.A(G169gat), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n902_), .B1(new_n900_), .B2(KEYINPUT62), .ZN(new_n903_));
  AND3_X1   g702(.A1(new_n899_), .A2(new_n901_), .A3(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n901_), .B1(new_n899_), .B2(new_n903_), .ZN(new_n905_));
  XOR2_X1   g704(.A(KEYINPUT22), .B(G169gat), .Z(new_n906_));
  OAI22_X1  g705(.A1(new_n904_), .A2(new_n905_), .B1(new_n899_), .B2(new_n906_), .ZN(G1348gat));
  AOI21_X1  g706(.A(G176gat), .B1(new_n898_), .B2(new_n648_), .ZN(new_n908_));
  AOI21_X1  g707(.A(KEYINPUT124), .B1(new_n842_), .B2(new_n462_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT124), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n845_), .A2(new_n910_), .A3(new_n391_), .ZN(new_n911_));
  OR2_X1    g710(.A1(new_n315_), .A2(new_n430_), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n909_), .A2(new_n911_), .A3(new_n912_), .ZN(new_n913_));
  AND2_X1   g712(.A1(new_n648_), .A2(G176gat), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n908_), .B1(new_n913_), .B2(new_n914_), .ZN(G1349gat));
  AOI211_X1 g714(.A(new_n607_), .B(new_n897_), .C1(new_n258_), .C2(new_n254_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n913_), .A2(new_n608_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(new_n218_), .ZN(G1350gat));
  OAI21_X1  g717(.A(G190gat), .B1(new_n897_), .B2(new_n569_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n654_), .A2(new_n211_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n897_), .B2(new_n920_), .ZN(G1351gat));
  NAND3_X1  g720(.A1(new_n464_), .A2(new_n316_), .A3(new_n467_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n845_), .A2(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n504_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g724(.A(KEYINPUT125), .ZN(new_n926_));
  OAI211_X1 g725(.A(new_n923_), .B(new_n648_), .C1(new_n926_), .C2(new_n237_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n237_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n927_), .B(new_n928_), .ZN(G1353gat));
  NOR3_X1   g728(.A1(new_n845_), .A2(new_n607_), .A3(new_n922_), .ZN(new_n930_));
  AND2_X1   g729(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n931_));
  NOR2_X1   g730(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n930_), .B1(new_n931_), .B2(new_n932_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n933_), .B1(new_n930_), .B2(new_n932_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(KEYINPUT126), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT126), .ZN(new_n936_));
  OAI211_X1 g735(.A(new_n933_), .B(new_n936_), .C1(new_n930_), .C2(new_n932_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n935_), .A2(new_n937_), .ZN(G1354gat));
  AOI21_X1  g737(.A(G218gat), .B1(new_n923_), .B2(new_n654_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n687_), .A2(G218gat), .ZN(new_n940_));
  XOR2_X1   g739(.A(new_n940_), .B(KEYINPUT127), .Z(new_n941_));
  AOI21_X1  g740(.A(new_n939_), .B1(new_n923_), .B2(new_n941_), .ZN(G1355gat));
endmodule


