//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 0 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n879_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n915_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_;
  XOR2_X1   g000(.A(G85gat), .B(G92gat), .Z(new_n202_));
  NOR2_X1   g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT65), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT66), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT7), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT66), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT65), .B1(new_n207_), .B2(new_n206_), .ZN(new_n208_));
  AOI22_X1  g007(.A1(new_n205_), .A2(new_n206_), .B1(new_n208_), .B2(new_n203_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  XOR2_X1   g009(.A(new_n210_), .B(KEYINPUT6), .Z(new_n211_));
  OAI21_X1  g010(.A(new_n202_), .B1(new_n209_), .B2(new_n211_), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n212_), .A2(KEYINPUT67), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(KEYINPUT67), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(KEYINPUT8), .A3(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT8), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n211_), .B(KEYINPUT64), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n216_), .B(new_n202_), .C1(new_n217_), .C2(new_n209_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n215_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n202_), .A2(KEYINPUT9), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  XOR2_X1   g020(.A(KEYINPUT10), .B(G99gat), .Z(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  OAI221_X1 g022(.A(new_n220_), .B1(KEYINPUT9), .B2(new_n221_), .C1(new_n223_), .C2(G106gat), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n217_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n219_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT68), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n226_), .B(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G29gat), .B(G36gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G43gat), .B(G50gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n228_), .A2(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n225_), .A2(KEYINPUT70), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n225_), .A2(KEYINPUT70), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(new_n219_), .A3(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(KEYINPUT73), .B(KEYINPUT15), .Z(new_n236_));
  XNOR2_X1  g035(.A(new_n231_), .B(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT35), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G232gat), .A2(G233gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT34), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  AOI22_X1  g040(.A1(new_n235_), .A2(new_n237_), .B1(new_n238_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n232_), .A2(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n241_), .A2(new_n238_), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n244_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G190gat), .B(G218gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G134gat), .B(G162gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(new_n250_), .B(KEYINPUT36), .Z(new_n251_));
  NAND2_X1  g050(.A1(new_n247_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT75), .ZN(new_n253_));
  INV_X1    g052(.A(new_n251_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n254_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT75), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT37), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n250_), .A2(KEYINPUT36), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n245_), .A2(new_n246_), .A3(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n253_), .A2(new_n257_), .A3(new_n258_), .A4(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT37), .B1(new_n260_), .B2(new_n255_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT74), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  OAI211_X1 g064(.A(KEYINPUT74), .B(KEYINPUT37), .C1(new_n260_), .C2(new_n255_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n262_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT69), .B(G71gat), .ZN(new_n268_));
  INV_X1    g067(.A(G78gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G57gat), .B(G64gat), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n271_), .A2(KEYINPUT11), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n271_), .B(KEYINPUT11), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(new_n270_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n226_), .A2(new_n227_), .ZN(new_n278_));
  AOI21_X1  g077(.A(KEYINPUT68), .B1(new_n219_), .B2(new_n225_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n277_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n235_), .A2(KEYINPUT12), .A3(new_n276_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G230gat), .A2(G233gat), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT12), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n284_), .B1(new_n228_), .B2(new_n277_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n282_), .A2(new_n283_), .A3(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n283_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n228_), .A2(new_n277_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n280_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n289_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n282_), .A2(new_n285_), .A3(KEYINPUT71), .A4(new_n283_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n288_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  XOR2_X1   g093(.A(G120gat), .B(G148gat), .Z(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G176gat), .B(G204gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n294_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n299_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n288_), .A2(new_n292_), .A3(new_n293_), .A4(new_n301_), .ZN(new_n302_));
  AND3_X1   g101(.A1(new_n300_), .A2(KEYINPUT13), .A3(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(KEYINPUT13), .B1(new_n300_), .B2(new_n302_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(G127gat), .B(G155gat), .Z(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT16), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G183gat), .B(G211gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT17), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT76), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G15gat), .B(G22gat), .ZN(new_n312_));
  INV_X1    g111(.A(G1gat), .ZN(new_n313_));
  INV_X1    g112(.A(G8gat), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT14), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n312_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G1gat), .B(G8gat), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n316_), .B(new_n317_), .Z(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n311_), .B(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G231gat), .A2(G233gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n322_), .A2(new_n277_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n309_), .A2(new_n310_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n277_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n323_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n326_), .B(KEYINPUT77), .Z(new_n327_));
  NAND3_X1  g126(.A1(new_n267_), .A2(new_n305_), .A3(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT78), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n237_), .A2(new_n319_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n231_), .B(KEYINPUT79), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(new_n318_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G229gat), .A2(G233gat), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n330_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n331_), .B(new_n319_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n334_), .B1(new_n335_), .B2(new_n333_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT80), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G113gat), .B(G141gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G169gat), .B(G197gat), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n338_), .B(new_n339_), .Z(new_n340_));
  XNOR2_X1  g139(.A(new_n337_), .B(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G155gat), .A2(G162gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345_));
  NOR3_X1   g144(.A1(new_n344_), .A2(new_n345_), .A3(KEYINPUT1), .ZN(new_n346_));
  INV_X1    g145(.A(G141gat), .ZN(new_n347_));
  INV_X1    g146(.A(G148gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G141gat), .A2(G148gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n349_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT90), .B1(new_n346_), .B2(new_n352_), .ZN(new_n353_));
  AND3_X1   g152(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n354_));
  AND2_X1   g153(.A1(G141gat), .A2(G148gat), .ZN(new_n355_));
  NOR2_X1   g154(.A1(G141gat), .A2(G148gat), .ZN(new_n356_));
  NOR3_X1   g155(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT90), .ZN(new_n358_));
  INV_X1    g157(.A(new_n345_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT1), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n359_), .A2(new_n360_), .A3(new_n343_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n357_), .A2(new_n358_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT91), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT3), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT3), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n356_), .A2(new_n363_), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT2), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n351_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n365_), .A2(new_n367_), .A3(new_n369_), .A4(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n344_), .A2(new_n345_), .ZN(new_n372_));
  AOI22_X1  g171(.A1(new_n353_), .A2(new_n362_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT29), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT28), .ZN(new_n376_));
  OR2_X1    g175(.A1(G197gat), .A2(G204gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G197gat), .A2(G204gat), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(KEYINPUT21), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT21), .ZN(new_n380_));
  AND2_X1   g179(.A1(G197gat), .A2(G204gat), .ZN(new_n381_));
  NOR2_X1   g180(.A1(G197gat), .A2(G204gat), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n380_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G211gat), .B(G218gat), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n379_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(G218gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(G211gat), .ZN(new_n387_));
  INV_X1    g186(.A(G211gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(G218gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n390_), .A2(KEYINPUT21), .A3(new_n377_), .A4(new_n378_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n385_), .A2(KEYINPUT93), .A3(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(KEYINPUT93), .B1(new_n385_), .B2(new_n391_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(G233gat), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n395_), .A2(KEYINPUT92), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n395_), .A2(KEYINPUT92), .ZN(new_n397_));
  OAI21_X1  g196(.A(G228gat), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n394_), .B(new_n398_), .C1(new_n374_), .C2(new_n373_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n385_), .A2(new_n391_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n400_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n398_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(KEYINPUT94), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(KEYINPUT94), .B1(new_n401_), .B2(new_n402_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n399_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G78gat), .B(G106gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT95), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n406_), .A2(new_n409_), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n399_), .B(new_n408_), .C1(new_n404_), .C2(new_n405_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n376_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G22gat), .B(G50gat), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n410_), .A2(new_n376_), .A3(new_n411_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n414_), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n410_), .A2(new_n376_), .A3(new_n411_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n417_), .B1(new_n418_), .B2(new_n412_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n416_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G227gat), .A2(G233gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT85), .ZN(new_n422_));
  INV_X1    g221(.A(G71gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(G99gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G15gat), .B(G43gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT86), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n425_), .B(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT87), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT81), .ZN(new_n430_));
  INV_X1    g229(.A(G169gat), .ZN(new_n431_));
  INV_X1    g230(.A(G176gat), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT24), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(G183gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT25), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT25), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(G183gat), .ZN(new_n441_));
  INV_X1    g240(.A(G190gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT26), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT26), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(G190gat), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n439_), .A2(new_n441_), .A3(new_n443_), .A4(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n436_), .B1(G169gat), .B2(G176gat), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(new_n434_), .A3(new_n433_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n437_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G183gat), .A2(G190gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT23), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT82), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n450_), .A2(KEYINPUT82), .A3(KEYINPUT23), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n450_), .A2(KEYINPUT83), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT83), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n457_), .A2(G183gat), .A3(G190gat), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT23), .B1(new_n456_), .B2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n455_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT84), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n461_), .B1(new_n450_), .B2(KEYINPUT23), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT23), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n463_), .A2(KEYINPUT84), .A3(G183gat), .A4(G190gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n456_), .A2(new_n458_), .A3(KEYINPUT23), .ZN(new_n466_));
  AOI22_X1  g265(.A1(new_n465_), .A2(new_n466_), .B1(new_n438_), .B2(new_n442_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(G169gat), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  OAI22_X1  g269(.A1(new_n449_), .A2(new_n460_), .B1(new_n467_), .B2(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(new_n471_), .B(KEYINPUT30), .Z(new_n472_));
  OAI21_X1  g271(.A(new_n428_), .B1(new_n429_), .B2(new_n472_), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n473_), .A2(KEYINPUT31), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(KEYINPUT31), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n472_), .A2(new_n429_), .ZN(new_n477_));
  XOR2_X1   g276(.A(G127gat), .B(G134gat), .Z(new_n478_));
  XOR2_X1   g277(.A(G113gat), .B(G120gat), .Z(new_n479_));
  INV_X1    g278(.A(KEYINPUT89), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G127gat), .B(G134gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G113gat), .B(G120gat), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT89), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(new_n483_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n485_), .A2(KEYINPUT88), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT88), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n487_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n481_), .B(new_n484_), .C1(new_n486_), .C2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n477_), .B(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n476_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n474_), .A2(new_n475_), .A3(new_n490_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NOR3_X1   g293(.A1(KEYINPUT91), .A2(G141gat), .A3(G148gat), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n369_), .B(new_n370_), .C1(new_n495_), .C2(new_n366_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n367_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n372_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NOR3_X1   g297(.A1(new_n346_), .A2(new_n352_), .A3(KEYINPUT90), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n358_), .B1(new_n357_), .B2(new_n361_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n498_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n481_), .A2(new_n484_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n485_), .B(KEYINPUT88), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n501_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G225gat), .A2(G233gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n478_), .A2(new_n479_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n485_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n498_), .B(new_n507_), .C1(new_n499_), .C2(new_n500_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n504_), .A2(new_n505_), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n504_), .A2(KEYINPUT4), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n508_), .B(KEYINPUT4), .C1(new_n489_), .C2(new_n373_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT100), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n504_), .A2(KEYINPUT100), .A3(KEYINPUT4), .A4(new_n508_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n511_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n505_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n510_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(G1gat), .B(G29gat), .Z(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT101), .B(G85gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT0), .B(G57gat), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n521_), .B(new_n522_), .Z(new_n523_));
  OR2_X1    g322(.A1(new_n518_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n518_), .A2(new_n523_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n494_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT103), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G226gat), .A2(G233gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT19), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n438_), .A2(new_n442_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n531_), .B1(new_n455_), .B2(new_n459_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT97), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  OAI211_X1 g333(.A(KEYINPUT97), .B(new_n531_), .C1(new_n455_), .C2(new_n459_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n470_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n448_), .A2(new_n446_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n465_), .A2(new_n466_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n436_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n537_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n400_), .B1(new_n536_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT98), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  OAI211_X1 g342(.A(KEYINPUT98), .B(new_n400_), .C1(new_n536_), .C2(new_n540_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT96), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n546_), .B(KEYINPUT20), .C1(new_n394_), .C2(new_n471_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n456_), .A2(new_n458_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n453_), .B(new_n454_), .C1(new_n549_), .C2(KEYINPUT23), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n550_), .A2(new_n537_), .A3(new_n437_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n538_), .A2(new_n531_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(new_n469_), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n551_), .B(new_n553_), .C1(new_n392_), .C2(new_n393_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n546_), .B1(new_n554_), .B2(KEYINPUT20), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n548_), .A2(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n530_), .B1(new_n545_), .B2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G8gat), .B(G36gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT18), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G64gat), .B(G92gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n559_), .B(new_n560_), .Z(new_n561_));
  NOR3_X1   g360(.A1(new_n536_), .A2(new_n400_), .A3(new_n540_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n394_), .A2(new_n471_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT20), .ZN(new_n564_));
  NOR3_X1   g363(.A1(new_n562_), .A2(new_n564_), .A3(new_n530_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n557_), .A2(new_n561_), .A3(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT20), .B1(new_n394_), .B2(new_n471_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT96), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(new_n547_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n530_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n570_), .A2(new_n571_), .A3(new_n543_), .A4(new_n544_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n530_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n561_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n567_), .B(KEYINPUT27), .C1(new_n574_), .C2(KEYINPUT102), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n574_), .A2(KEYINPUT102), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n528_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n574_), .A2(KEYINPUT102), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n574_), .A2(KEYINPUT102), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT27), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n543_), .B(new_n544_), .C1(new_n555_), .C2(new_n548_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n565_), .B1(new_n581_), .B2(new_n530_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n580_), .B1(new_n582_), .B2(new_n561_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n578_), .A2(KEYINPUT103), .A3(new_n579_), .A4(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n577_), .A2(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(KEYINPUT99), .B1(new_n582_), .B2(new_n561_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n557_), .A2(new_n566_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n561_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n586_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n587_), .A2(KEYINPUT99), .A3(new_n588_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n590_), .A2(new_n580_), .A3(new_n591_), .ZN(new_n592_));
  AND4_X1   g391(.A1(new_n420_), .A2(new_n527_), .A3(new_n585_), .A4(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n494_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n526_), .B1(new_n416_), .B2(new_n419_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n585_), .A2(new_n592_), .A3(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n516_), .A2(new_n505_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n523_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n504_), .A2(new_n517_), .A3(new_n508_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n597_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT33), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n516_), .A2(new_n517_), .ZN(new_n602_));
  AND4_X1   g401(.A1(new_n601_), .A2(new_n602_), .A3(new_n523_), .A4(new_n509_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n601_), .B1(new_n518_), .B2(new_n523_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n600_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n605_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT32), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n582_), .B1(new_n607_), .B2(new_n588_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n572_), .A2(new_n573_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n609_), .A2(KEYINPUT32), .A3(new_n561_), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n526_), .A2(new_n608_), .A3(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n420_), .B1(new_n606_), .B2(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n594_), .B1(new_n596_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT104), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n593_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n577_), .A2(new_n584_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n595_), .A2(new_n592_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n612_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(new_n494_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT104), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n342_), .B1(new_n615_), .B2(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n329_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n622_), .A2(new_n313_), .A3(new_n526_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT105), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT38), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n625_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n615_), .A2(new_n620_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n253_), .A2(new_n261_), .A3(new_n257_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n327_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n628_), .A2(new_n632_), .A3(new_n341_), .A4(new_n305_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT106), .Z(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n526_), .ZN(new_n636_));
  OAI21_X1  g435(.A(G1gat), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n626_), .A2(new_n627_), .A3(new_n637_), .ZN(G1324gat));
  AND2_X1   g437(.A1(new_n585_), .A2(new_n592_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n622_), .A2(new_n314_), .A3(new_n640_), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n633_), .A2(new_n639_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT39), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n642_), .A2(new_n643_), .A3(G8gat), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n643_), .B1(new_n642_), .B2(G8gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n641_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT108), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT108), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n641_), .B(new_n648_), .C1(new_n644_), .C2(new_n645_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(G1325gat));
  INV_X1    g451(.A(G15gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(new_n634_), .B2(new_n594_), .ZN(new_n654_));
  XOR2_X1   g453(.A(KEYINPUT109), .B(KEYINPUT41), .Z(new_n655_));
  OR2_X1    g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n655_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n622_), .A2(new_n653_), .A3(new_n594_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n656_), .A2(new_n657_), .A3(new_n658_), .ZN(G1326gat));
  INV_X1    g458(.A(G22gat), .ZN(new_n660_));
  INV_X1    g459(.A(new_n420_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n634_), .B2(new_n661_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT42), .Z(new_n663_));
  NAND3_X1  g462(.A1(new_n622_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1327gat));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n262_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n628_), .A2(new_n667_), .A3(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT110), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n618_), .A2(new_n614_), .A3(new_n494_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n593_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n613_), .A2(new_n614_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n671_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n615_), .A2(new_n620_), .A3(KEYINPUT110), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n676_), .A2(new_n667_), .A3(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT43), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT111), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n678_), .A2(KEYINPUT111), .A3(KEYINPUT43), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n670_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n305_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n684_), .A2(new_n342_), .A3(new_n327_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n666_), .B1(new_n683_), .B2(new_n686_), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n678_), .A2(KEYINPUT111), .A3(KEYINPUT43), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT111), .B1(new_n678_), .B2(KEYINPUT43), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n669_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n690_), .A2(KEYINPUT44), .A3(new_n685_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n687_), .A2(G29gat), .A3(new_n526_), .A4(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(G29gat), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n629_), .A2(new_n327_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n621_), .A2(new_n305_), .A3(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n693_), .B1(new_n695_), .B2(new_n636_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n692_), .A2(new_n696_), .ZN(G1328gat));
  NAND3_X1  g496(.A1(new_n687_), .A2(new_n640_), .A3(new_n691_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(G36gat), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n695_), .A2(G36gat), .A3(new_n639_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT45), .Z(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT46), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n699_), .A2(KEYINPUT46), .A3(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1329gat));
  NAND4_X1  g505(.A1(new_n687_), .A2(G43gat), .A3(new_n594_), .A4(new_n691_), .ZN(new_n707_));
  INV_X1    g506(.A(G43gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n708_), .B1(new_n695_), .B2(new_n494_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT112), .Z(new_n710_));
  NAND2_X1  g509(.A1(new_n707_), .A2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g511(.A1(new_n687_), .A2(G50gat), .A3(new_n661_), .A4(new_n691_), .ZN(new_n713_));
  INV_X1    g512(.A(G50gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n714_), .B1(new_n695_), .B2(new_n420_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1331gat));
  NOR2_X1   g515(.A1(new_n305_), .A2(new_n341_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n717_), .A2(new_n628_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n718_), .A2(new_n632_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n719_), .A2(G57gat), .A3(new_n526_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT113), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n720_), .A2(new_n721_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n718_), .A2(new_n327_), .A3(new_n267_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(G57gat), .B1(new_n725_), .B2(new_n526_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n722_), .A2(new_n723_), .A3(new_n726_), .ZN(G1332gat));
  INV_X1    g526(.A(G64gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n719_), .B2(new_n640_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT48), .Z(new_n730_));
  NAND3_X1  g529(.A1(new_n725_), .A2(new_n728_), .A3(new_n640_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1333gat));
  AOI21_X1  g531(.A(new_n423_), .B1(new_n719_), .B2(new_n594_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT49), .Z(new_n734_));
  NAND3_X1  g533(.A1(new_n725_), .A2(new_n423_), .A3(new_n594_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1334gat));
  AOI21_X1  g535(.A(new_n269_), .B1(new_n719_), .B2(new_n661_), .ZN(new_n737_));
  XOR2_X1   g536(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n738_));
  XNOR2_X1  g537(.A(new_n737_), .B(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n725_), .A2(new_n269_), .A3(new_n661_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1335gat));
  INV_X1    g540(.A(G85gat), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n718_), .A2(new_n694_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n742_), .B1(new_n743_), .B2(new_n636_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT115), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n717_), .A2(new_n631_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n683_), .A2(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n636_), .A2(new_n742_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n745_), .B1(new_n747_), .B2(new_n748_), .ZN(G1336gat));
  INV_X1    g548(.A(new_n743_), .ZN(new_n750_));
  INV_X1    g549(.A(G92gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(new_n751_), .A3(new_n640_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n683_), .A2(new_n639_), .A3(new_n746_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n752_), .B1(new_n753_), .B2(new_n751_), .ZN(G1337gat));
  INV_X1    g553(.A(KEYINPUT117), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n755_), .A2(KEYINPUT51), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n750_), .A2(new_n594_), .A3(new_n222_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT116), .ZN(new_n758_));
  INV_X1    g557(.A(new_n746_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n690_), .A2(new_n594_), .A3(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(G99gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n756_), .B1(new_n758_), .B2(new_n761_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n755_), .A2(KEYINPUT51), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n762_), .B(new_n763_), .ZN(G1338gat));
  OR3_X1    g563(.A1(new_n743_), .A2(G106gat), .A3(new_n420_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n690_), .A2(new_n661_), .A3(new_n759_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n766_), .A2(new_n767_), .A3(G106gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n766_), .B2(G106gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n765_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT53), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n772_), .B(new_n765_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1339gat));
  INV_X1    g573(.A(new_n333_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n335_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n330_), .A2(new_n332_), .A3(new_n775_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n340_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n336_), .A2(new_n340_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n781_), .B1(new_n300_), .B2(new_n302_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT119), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n782_), .B(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n302_), .A2(new_n341_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n288_), .A2(new_n786_), .A3(new_n293_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n278_), .A2(new_n279_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT12), .B1(new_n788_), .B2(new_n276_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n280_), .A2(new_n281_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n289_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT118), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT118), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n793_), .B(new_n289_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n792_), .B(new_n794_), .C1(new_n786_), .C2(new_n286_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n299_), .B1(new_n787_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT56), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n288_), .A2(new_n786_), .A3(new_n293_), .ZN(new_n799_));
  OR2_X1    g598(.A1(new_n286_), .A2(new_n786_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n799_), .A2(new_n794_), .A3(new_n800_), .A4(new_n792_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n801_), .A2(KEYINPUT56), .A3(new_n299_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n785_), .B1(new_n798_), .B2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n629_), .B1(new_n784_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n805_));
  INV_X1    g604(.A(new_n781_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n302_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n796_), .A2(new_n797_), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT56), .B1(new_n801_), .B2(new_n299_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n808_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT58), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n267_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  AOI211_X1 g612(.A(new_n812_), .B(new_n807_), .C1(new_n798_), .C2(new_n802_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  AOI22_X1  g614(.A1(new_n804_), .A2(new_n805_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n785_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n300_), .A2(new_n302_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n783_), .B1(new_n819_), .B2(new_n806_), .ZN(new_n820_));
  AOI211_X1 g619(.A(KEYINPUT119), .B(new_n781_), .C1(new_n300_), .C2(new_n302_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n630_), .B1(new_n818_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT57), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n327_), .B1(new_n816_), .B2(new_n824_), .ZN(new_n825_));
  OR3_X1    g624(.A1(new_n328_), .A2(KEYINPUT54), .A3(new_n341_), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT54), .B1(new_n328_), .B2(new_n341_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n825_), .A2(new_n829_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n640_), .A2(new_n661_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(new_n594_), .A3(new_n526_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(G113gat), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n834_), .A3(new_n341_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n807_), .B1(new_n798_), .B2(new_n802_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n667_), .B1(new_n836_), .B2(KEYINPUT58), .ZN(new_n837_));
  OAI22_X1  g636(.A1(new_n823_), .A2(KEYINPUT57), .B1(new_n837_), .B2(new_n814_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n804_), .A2(new_n805_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n631_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n828_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n832_), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT59), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n845_));
  AOI211_X1 g644(.A(new_n845_), .B(new_n832_), .C1(new_n840_), .C2(new_n828_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n342_), .B1(new_n844_), .B2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n835_), .B1(new_n848_), .B2(new_n834_), .ZN(G1340gat));
  AOI21_X1  g648(.A(new_n305_), .B1(new_n844_), .B2(new_n847_), .ZN(new_n850_));
  INV_X1    g649(.A(G120gat), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT60), .ZN(new_n853_));
  AOI21_X1  g652(.A(G120gat), .B1(new_n684_), .B2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n854_), .B1(new_n853_), .B2(G120gat), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n833_), .A2(new_n852_), .A3(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n852_), .B1(new_n833_), .B2(new_n855_), .ZN(new_n857_));
  OAI22_X1  g656(.A1(new_n850_), .A2(new_n851_), .B1(new_n856_), .B2(new_n857_), .ZN(G1341gat));
  INV_X1    g657(.A(G127gat), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n631_), .A2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n843_), .B2(new_n846_), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n327_), .B(new_n842_), .C1(new_n825_), .C2(new_n829_), .ZN(new_n862_));
  AND3_X1   g661(.A1(new_n862_), .A2(KEYINPUT121), .A3(new_n859_), .ZN(new_n863_));
  AOI21_X1  g662(.A(KEYINPUT121), .B1(new_n862_), .B2(new_n859_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n861_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT122), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT122), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n861_), .B(new_n867_), .C1(new_n863_), .C2(new_n864_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(G1342gat));
  INV_X1    g668(.A(G134gat), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n833_), .A2(new_n870_), .A3(new_n630_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n267_), .B1(new_n844_), .B2(new_n847_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(new_n870_), .ZN(G1343gat));
  NAND4_X1  g672(.A1(new_n639_), .A2(new_n494_), .A3(new_n661_), .A4(new_n526_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n830_), .A2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n341_), .ZN(new_n876_));
  XOR2_X1   g675(.A(KEYINPUT123), .B(G141gat), .Z(new_n877_));
  XNOR2_X1  g676(.A(new_n876_), .B(new_n877_), .ZN(G1344gat));
  NAND2_X1  g677(.A1(new_n875_), .A2(new_n684_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g679(.A1(new_n875_), .A2(new_n327_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(KEYINPUT61), .B(G155gat), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n881_), .B(new_n882_), .ZN(G1346gat));
  INV_X1    g682(.A(G162gat), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n875_), .A2(new_n884_), .A3(new_n630_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n830_), .A2(new_n267_), .A3(new_n874_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n886_), .B2(new_n884_), .ZN(G1347gat));
  NOR2_X1   g686(.A1(new_n830_), .A2(new_n661_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n639_), .A2(new_n494_), .A3(new_n526_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT22), .B(G169gat), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n891_), .A2(new_n341_), .A3(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n889_), .A2(new_n341_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(KEYINPUT124), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n888_), .A2(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n894_), .B1(new_n897_), .B2(G169gat), .ZN(new_n898_));
  AOI211_X1 g697(.A(KEYINPUT62), .B(new_n431_), .C1(new_n888_), .C2(new_n896_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n893_), .B1(new_n898_), .B2(new_n899_), .ZN(G1348gat));
  AOI21_X1  g699(.A(G176gat), .B1(new_n891_), .B2(new_n684_), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n890_), .A2(new_n432_), .A3(new_n305_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1349gat));
  NAND2_X1  g702(.A1(new_n439_), .A2(new_n441_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n891_), .A2(new_n904_), .A3(new_n327_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n438_), .B1(new_n890_), .B2(new_n631_), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1350gat));
  NAND4_X1  g706(.A1(new_n891_), .A2(new_n443_), .A3(new_n445_), .A4(new_n630_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n888_), .A2(new_n667_), .A3(new_n889_), .ZN(new_n909_));
  AND3_X1   g708(.A1(new_n909_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n910_));
  AOI21_X1  g709(.A(KEYINPUT125), .B1(new_n909_), .B2(G190gat), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n908_), .B1(new_n910_), .B2(new_n911_), .ZN(G1351gat));
  NAND3_X1  g711(.A1(new_n640_), .A2(new_n494_), .A3(new_n595_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n830_), .A2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(new_n341_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g715(.A(KEYINPUT127), .ZN(new_n917_));
  INV_X1    g716(.A(new_n913_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n841_), .A2(new_n684_), .A3(new_n918_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n917_), .B1(new_n919_), .B2(G204gat), .ZN(new_n920_));
  OR2_X1    g719(.A1(new_n919_), .A2(KEYINPUT126), .ZN(new_n921_));
  INV_X1    g720(.A(G204gat), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n922_), .B1(new_n919_), .B2(KEYINPUT126), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n920_), .B1(new_n921_), .B2(new_n923_), .ZN(new_n924_));
  AND2_X1   g723(.A1(new_n921_), .A2(new_n923_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n924_), .B1(KEYINPUT127), .B2(new_n925_), .ZN(G1353gat));
  NAND2_X1  g725(.A1(new_n914_), .A2(new_n327_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n928_));
  AND2_X1   g727(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n927_), .A2(new_n928_), .A3(new_n929_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n930_), .B1(new_n927_), .B2(new_n928_), .ZN(G1354gat));
  NAND3_X1  g730(.A1(new_n914_), .A2(new_n386_), .A3(new_n630_), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n830_), .A2(new_n267_), .A3(new_n913_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n933_), .B2(new_n386_), .ZN(G1355gat));
endmodule


