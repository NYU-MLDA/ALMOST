//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 0 0 0 0 0 0 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n892_, new_n893_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G1gat), .B(G29gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G85gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT0), .B(G57gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  AND2_X1   g006(.A1(KEYINPUT88), .A2(KEYINPUT2), .ZN(new_n208_));
  NOR2_X1   g007(.A1(KEYINPUT88), .A2(KEYINPUT2), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n207_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT89), .ZN(new_n211_));
  AND3_X1   g010(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n212_));
  INV_X1    g011(.A(G141gat), .ZN(new_n213_));
  INV_X1    g012(.A(G148gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT87), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n213_), .B(new_n214_), .C1(new_n215_), .C2(KEYINPUT3), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n217_), .B(KEYINPUT87), .C1(G141gat), .C2(G148gat), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n212_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT89), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n220_), .B(new_n207_), .C1(new_n208_), .C2(new_n209_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n211_), .A2(new_n219_), .A3(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(G155gat), .B(G162gat), .Z(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n213_), .A2(new_n214_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(new_n207_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G155gat), .A2(G162gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G155gat), .A2(G162gat), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n227_), .B1(KEYINPUT1), .B2(new_n228_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n228_), .A2(KEYINPUT1), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n226_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n224_), .A2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G127gat), .B(G134gat), .Z(new_n234_));
  XOR2_X1   g033(.A(G113gat), .B(G120gat), .Z(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n233_), .A2(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n231_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(new_n236_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(KEYINPUT4), .A3(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G225gat), .A2(G233gat), .ZN(new_n242_));
  XOR2_X1   g041(.A(new_n242_), .B(KEYINPUT96), .Z(new_n243_));
  INV_X1    g042(.A(KEYINPUT98), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n236_), .B1(new_n224_), .B2(new_n232_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT97), .B(KEYINPUT4), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n244_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n248_));
  NOR4_X1   g047(.A1(new_n239_), .A2(KEYINPUT98), .A3(new_n236_), .A4(new_n246_), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n241_), .B(new_n243_), .C1(new_n248_), .C2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n243_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n238_), .A2(new_n240_), .A3(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n206_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n206_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n239_), .B(new_n237_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n251_), .B1(new_n255_), .B2(KEYINPUT4), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT98), .B1(new_n238_), .B2(new_n246_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n249_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n254_), .B1(new_n256_), .B2(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n253_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT28), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT29), .ZN(new_n263_));
  AND4_X1   g062(.A1(new_n262_), .A2(new_n224_), .A3(new_n263_), .A4(new_n232_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n262_), .B1(new_n239_), .B2(new_n263_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G22gat), .B(G50gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NOR3_X1   g066(.A1(new_n264_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n224_), .A2(new_n263_), .A3(new_n232_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT28), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n239_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n266_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n268_), .A2(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(G211gat), .B(G218gat), .Z(new_n274_));
  INV_X1    g073(.A(KEYINPUT21), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G197gat), .B(G204gat), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n274_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(KEYINPUT91), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT91), .ZN(new_n279_));
  INV_X1    g078(.A(G197gat), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(new_n280_), .A3(G204gat), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n278_), .A2(KEYINPUT21), .A3(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n277_), .A2(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n276_), .A2(new_n275_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(new_n274_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n286_), .B1(new_n239_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(KEYINPUT90), .A2(G233gat), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(KEYINPUT90), .A2(G233gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(G228gat), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n288_), .A2(new_n293_), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n286_), .B(new_n292_), .C1(new_n239_), .C2(new_n263_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(G78gat), .B(G106gat), .Z(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n297_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n294_), .A2(new_n295_), .A3(new_n299_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n273_), .A2(new_n298_), .A3(KEYINPUT93), .A4(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT93), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n302_), .B1(new_n268_), .B2(new_n272_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n267_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n270_), .A2(new_n271_), .A3(new_n266_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n305_), .A2(new_n306_), .A3(KEYINPUT93), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n294_), .A2(new_n295_), .A3(new_n299_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n299_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n307_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n261_), .B(new_n301_), .C1(new_n304_), .C2(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(G8gat), .B(G36gat), .Z(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G64gat), .B(G92gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G226gat), .A2(G233gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT19), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT20), .ZN(new_n321_));
  INV_X1    g120(.A(G169gat), .ZN(new_n322_));
  INV_X1    g121(.A(G176gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n324_), .A2(KEYINPUT24), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G183gat), .A2(G190gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT23), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT83), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT83), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n326_), .A2(new_n329_), .A3(KEYINPUT23), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(G183gat), .A3(G190gat), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n325_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT25), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(G183gat), .ZN(new_n336_));
  INV_X1    g135(.A(G183gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT25), .ZN(new_n338_));
  INV_X1    g137(.A(G190gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT26), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT26), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(G190gat), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n336_), .A2(new_n338_), .A3(new_n340_), .A4(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G169gat), .A2(G176gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n324_), .A2(KEYINPUT24), .A3(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT94), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT94), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n343_), .A2(new_n348_), .A3(new_n345_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n334_), .A2(new_n347_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT81), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n326_), .A2(new_n351_), .A3(KEYINPUT23), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n351_), .B1(new_n326_), .B2(KEYINPUT23), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n333_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(G183gat), .A2(G190gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT22), .B(G169gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(new_n323_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n359_), .A2(new_n344_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n350_), .A2(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n321_), .B1(new_n362_), .B2(new_n286_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT82), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n364_), .B1(new_n358_), .B2(new_n323_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n322_), .A2(KEYINPUT22), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT22), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(G169gat), .ZN(new_n368_));
  AND4_X1   g167(.A1(new_n364_), .A2(new_n366_), .A3(new_n368_), .A4(new_n323_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n333_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n370_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n371_));
  OAI221_X1 g170(.A(new_n344_), .B1(new_n365_), .B2(new_n369_), .C1(new_n371_), .C2(new_n355_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n336_), .A2(KEYINPUT80), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT26), .B(G190gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT25), .B(G183gat), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n373_), .B(new_n374_), .C1(new_n375_), .C2(KEYINPUT80), .ZN(new_n376_));
  INV_X1    g175(.A(new_n325_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n376_), .A2(new_n354_), .A3(new_n345_), .A4(new_n377_), .ZN(new_n378_));
  AOI22_X1  g177(.A1(new_n277_), .A2(new_n282_), .B1(new_n274_), .B2(new_n284_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n372_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n320_), .B1(new_n363_), .B2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n344_), .B1(new_n365_), .B2(new_n369_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n355_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n378_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n286_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n350_), .A2(new_n379_), .A3(new_n361_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n385_), .A2(new_n386_), .A3(KEYINPUT20), .A4(new_n320_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n317_), .B1(new_n381_), .B2(new_n388_), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n343_), .A2(new_n348_), .A3(new_n345_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n348_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  AOI22_X1  g191(.A1(new_n392_), .A2(new_n334_), .B1(new_n357_), .B2(new_n360_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n380_), .B(KEYINPUT20), .C1(new_n393_), .C2(new_n379_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n319_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n395_), .A2(new_n316_), .A3(new_n387_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n389_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT27), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n385_), .A2(new_n386_), .A3(KEYINPUT20), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n319_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n362_), .A2(new_n286_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n402_), .A2(KEYINPUT20), .A3(new_n320_), .A4(new_n380_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(new_n317_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n405_), .A2(KEYINPUT27), .A3(new_n396_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n399_), .A2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT104), .B1(new_n311_), .B2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n381_), .A2(new_n388_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n398_), .B1(new_n409_), .B2(new_n316_), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n405_), .A2(new_n410_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n301_), .B1(new_n310_), .B2(new_n304_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT104), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n411_), .A2(new_n413_), .A3(new_n414_), .A4(new_n261_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n408_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n316_), .A2(KEYINPUT32), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n418_), .B1(new_n401_), .B2(new_n403_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT102), .ZN(new_n420_));
  INV_X1    g219(.A(new_n206_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n421_), .B1(new_n255_), .B2(new_n251_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n250_), .A2(new_n422_), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n250_), .A2(new_n252_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n423_), .B1(new_n424_), .B2(new_n206_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n395_), .A2(new_n387_), .A3(new_n418_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n420_), .A2(KEYINPUT103), .A3(new_n425_), .A4(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT103), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n419_), .A2(KEYINPUT102), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT102), .ZN(new_n430_));
  AOI211_X1 g229(.A(new_n430_), .B(new_n418_), .C1(new_n401_), .C2(new_n403_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n426_), .B1(new_n253_), .B2(new_n260_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n428_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n427_), .A2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n250_), .A2(KEYINPUT33), .A3(new_n422_), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n436_), .A2(new_n396_), .A3(new_n389_), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n241_), .B(new_n251_), .C1(new_n248_), .C2(new_n249_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n206_), .B1(new_n255_), .B2(new_n243_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT100), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT100), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n438_), .A2(new_n442_), .A3(new_n439_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n437_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT33), .ZN(new_n446_));
  AOI21_X1  g245(.A(KEYINPUT99), .B1(new_n423_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT99), .ZN(new_n448_));
  AOI211_X1 g247(.A(new_n448_), .B(KEYINPUT33), .C1(new_n250_), .C2(new_n422_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT101), .B1(new_n445_), .B2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n448_), .B1(new_n260_), .B2(KEYINPUT33), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n423_), .A2(KEYINPUT99), .A3(new_n446_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT101), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n454_), .A2(new_n455_), .A3(new_n444_), .A4(new_n437_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n435_), .B1(new_n451_), .B2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n417_), .B1(new_n457_), .B2(new_n413_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n236_), .B(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n460_), .B(KEYINPUT86), .Z(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G71gat), .B(G99gat), .ZN(new_n463_));
  INV_X1    g262(.A(G43gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G227gat), .A2(G233gat), .ZN(new_n466_));
  INV_X1    g265(.A(G15gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n465_), .B(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n384_), .B(KEYINPUT30), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT84), .ZN(new_n471_));
  OR2_X1    g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n471_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n469_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n469_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n462_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n470_), .B(KEYINPUT84), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n475_), .B(new_n461_), .C1(new_n478_), .C2(new_n469_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n480_), .A2(new_n425_), .ZN(new_n481_));
  AOI21_X1  g280(.A(KEYINPUT105), .B1(new_n411_), .B2(new_n412_), .ZN(new_n482_));
  AND4_X1   g281(.A1(KEYINPUT105), .A2(new_n412_), .A3(new_n399_), .A4(new_n406_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n481_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT106), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT106), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n486_), .B(new_n481_), .C1(new_n482_), .C2(new_n483_), .ZN(new_n487_));
  AOI22_X1  g286(.A1(new_n458_), .A2(new_n480_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G190gat), .B(G218gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G134gat), .B(G162gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n491_), .A2(KEYINPUT36), .ZN(new_n492_));
  XOR2_X1   g291(.A(KEYINPUT10), .B(G99gat), .Z(new_n493_));
  INV_X1    g292(.A(G106gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT65), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT66), .B(G85gat), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT9), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n497_), .A2(new_n498_), .A3(G92gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G99gat), .A2(G106gat), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT6), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(G85gat), .B(G92gat), .Z(new_n503_));
  AOI21_X1  g302(.A(new_n502_), .B1(KEYINPUT9), .B2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n496_), .A2(new_n499_), .A3(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(G99gat), .A2(G106gat), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT7), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n503_), .B1(new_n508_), .B2(new_n502_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT8), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n505_), .A2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G29gat), .B(G36gat), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n512_), .A2(KEYINPUT72), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n512_), .A2(KEYINPUT72), .ZN(new_n514_));
  XOR2_X1   g313(.A(G43gat), .B(G50gat), .Z(new_n515_));
  OR3_X1    g314(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n515_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n511_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT74), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G232gat), .A2(G233gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n524_), .A2(KEYINPUT35), .ZN(new_n525_));
  XOR2_X1   g324(.A(KEYINPUT73), .B(KEYINPUT15), .Z(new_n526_));
  XNOR2_X1  g325(.A(new_n518_), .B(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n525_), .B1(new_n527_), .B2(new_n511_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n520_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT76), .ZN(new_n530_));
  AOI21_X1  g329(.A(KEYINPUT75), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n520_), .A2(new_n528_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT75), .ZN(new_n533_));
  OAI211_X1 g332(.A(KEYINPUT35), .B(new_n524_), .C1(new_n532_), .C2(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n531_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n524_), .A2(KEYINPUT35), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n533_), .B(new_n536_), .C1(new_n532_), .C2(KEYINPUT76), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n492_), .B1(new_n535_), .B2(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n536_), .B1(new_n529_), .B2(KEYINPUT75), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n533_), .B1(new_n532_), .B2(KEYINPUT76), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n491_), .B(KEYINPUT36), .Z(new_n543_));
  NAND3_X1  g342(.A1(new_n542_), .A2(new_n537_), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n539_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G57gat), .B(G64gat), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT67), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT11), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT68), .ZN(new_n551_));
  XOR2_X1   g350(.A(G71gat), .B(G78gat), .Z(new_n552_));
  OAI21_X1  g351(.A(new_n552_), .B1(new_n549_), .B2(KEYINPUT11), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n551_), .A2(new_n553_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G15gat), .B(G22gat), .ZN(new_n557_));
  INV_X1    g356(.A(G8gat), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G1gat), .B(G8gat), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n560_), .B(new_n561_), .Z(new_n562_));
  NAND2_X1  g361(.A1(G231gat), .A2(G233gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n556_), .B(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G127gat), .B(G155gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(G183gat), .B(G211gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT69), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n571_), .A2(KEYINPUT17), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n565_), .A2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n573_), .B1(KEYINPUT17), .B2(new_n570_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n575_), .B1(new_n565_), .B2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n571_), .A2(KEYINPUT12), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n511_), .A2(new_n579_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n511_), .A2(KEYINPUT12), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n556_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n554_), .A2(new_n511_), .A3(new_n555_), .A4(new_n579_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G230gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT64), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n584_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n556_), .A2(new_n510_), .A3(new_n505_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n554_), .A2(new_n511_), .A3(new_n555_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n589_), .A2(new_n586_), .A3(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n588_), .A2(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(G120gat), .B(G148gat), .Z(new_n593_));
  XNOR2_X1  g392(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G176gat), .B(G204gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n592_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n588_), .A2(new_n591_), .A3(new_n597_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT13), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT13), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n599_), .A2(new_n603_), .A3(new_n600_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G113gat), .B(G141gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G169gat), .B(G197gat), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n606_), .B(new_n607_), .Z(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n562_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT78), .ZN(new_n611_));
  INV_X1    g410(.A(new_n562_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(new_n518_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G229gat), .A2(G233gat), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n527_), .A2(new_n612_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n617_), .A2(new_n611_), .A3(new_n615_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n609_), .B1(new_n616_), .B2(new_n619_), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n618_), .B(new_n608_), .C1(new_n614_), .C2(new_n615_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n620_), .A2(KEYINPUT79), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT79), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n623_), .B(new_n609_), .C1(new_n616_), .C2(new_n619_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n605_), .A2(new_n626_), .ZN(new_n627_));
  NOR4_X1   g426(.A1(new_n488_), .A2(new_n546_), .A3(new_n577_), .A4(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT107), .Z(new_n629_));
  AOI21_X1  g428(.A(new_n202_), .B1(new_n629_), .B2(new_n425_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT108), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n488_), .A2(new_n625_), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n542_), .A2(new_n537_), .A3(new_n543_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n492_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n634_), .B1(new_n542_), .B2(new_n537_), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT37), .B1(new_n633_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT37), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n539_), .A2(new_n637_), .A3(new_n544_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n577_), .B1(new_n602_), .B2(new_n604_), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n632_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n641_), .A2(new_n202_), .A3(new_n425_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT38), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n631_), .A2(new_n643_), .ZN(G1324gat));
  NAND3_X1  g443(.A1(new_n641_), .A2(new_n558_), .A3(new_n407_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n628_), .A2(new_n407_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(KEYINPUT109), .B(KEYINPUT39), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n646_), .A2(G8gat), .A3(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n647_), .B1(new_n646_), .B2(G8gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n645_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n650_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g450(.A(new_n480_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n467_), .B1(new_n629_), .B2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT41), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n641_), .A2(new_n467_), .A3(new_n652_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1326gat));
  INV_X1    g455(.A(G22gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n657_), .B1(new_n629_), .B2(new_n413_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT42), .Z(new_n659_));
  NAND3_X1  g458(.A1(new_n641_), .A2(new_n657_), .A3(new_n413_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1327gat));
  INV_X1    g460(.A(new_n577_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n545_), .A2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT112), .ZN(new_n664_));
  INV_X1    g463(.A(new_n605_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(new_n632_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(G29gat), .B1(new_n668_), .B2(new_n425_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT43), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n670_), .A2(KEYINPUT110), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n485_), .A2(new_n487_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n451_), .A2(new_n456_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n427_), .A2(new_n434_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n416_), .B1(new_n675_), .B2(new_n412_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n672_), .B1(new_n676_), .B2(new_n652_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n633_), .A2(new_n635_), .A3(KEYINPUT37), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n637_), .B1(new_n539_), .B2(new_n544_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n677_), .A2(new_n680_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n670_), .A2(KEYINPUT110), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n671_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT111), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n684_), .B(new_n672_), .C1(new_n676_), .C2(new_n652_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n670_), .A2(KEYINPUT111), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n685_), .B(new_n680_), .C1(new_n488_), .C2(new_n686_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n627_), .A2(new_n662_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n683_), .A2(new_n687_), .A3(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n683_), .A2(KEYINPUT44), .A3(new_n687_), .A4(new_n688_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n425_), .A2(G29gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n669_), .B1(new_n693_), .B2(new_n694_), .ZN(G1328gat));
  OR2_X1    g494(.A1(new_n411_), .A2(G36gat), .ZN(new_n696_));
  OR3_X1    g495(.A1(new_n667_), .A2(KEYINPUT45), .A3(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT45), .B1(new_n667_), .B2(new_n696_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n691_), .A2(new_n407_), .A3(new_n692_), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n700_), .A2(KEYINPUT113), .A3(G36gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(KEYINPUT113), .B1(new_n700_), .B2(G36gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n699_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT46), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n699_), .B(KEYINPUT46), .C1(new_n701_), .C2(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1329gat));
  NAND3_X1  g506(.A1(new_n693_), .A2(G43gat), .A3(new_n652_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n464_), .B1(new_n667_), .B2(new_n480_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g510(.A(G50gat), .B1(new_n668_), .B2(new_n413_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n413_), .A2(G50gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n693_), .B2(new_n713_), .ZN(G1331gat));
  NOR2_X1   g513(.A1(new_n488_), .A2(new_n546_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n665_), .A2(new_n662_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n716_), .A2(new_n626_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n715_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G57gat), .B1(new_n719_), .B2(new_n261_), .ZN(new_n720_));
  NOR4_X1   g519(.A1(new_n488_), .A2(new_n680_), .A3(new_n716_), .A4(new_n626_), .ZN(new_n721_));
  INV_X1    g520(.A(G57gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n722_), .A3(new_n425_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n720_), .A2(new_n723_), .ZN(G1332gat));
  INV_X1    g523(.A(G64gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n718_), .B2(new_n407_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT48), .Z(new_n727_));
  NAND3_X1  g526(.A1(new_n721_), .A2(new_n725_), .A3(new_n407_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1333gat));
  INV_X1    g528(.A(G71gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n730_), .B1(new_n718_), .B2(new_n652_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(KEYINPUT114), .B(KEYINPUT49), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n731_), .B(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n721_), .A2(new_n730_), .A3(new_n652_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1334gat));
  INV_X1    g534(.A(G78gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n736_), .B1(new_n718_), .B2(new_n413_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n737_), .B(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n721_), .A2(new_n736_), .A3(new_n413_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1335gat));
  INV_X1    g540(.A(G85gat), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n664_), .A2(new_n605_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n488_), .A2(new_n626_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n742_), .B1(new_n745_), .B2(new_n261_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT116), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n425_), .A2(new_n497_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n682_), .B1(new_n488_), .B2(new_n639_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n671_), .ZN(new_n750_));
  NOR3_X1   g549(.A1(new_n605_), .A2(new_n662_), .A3(new_n626_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n687_), .A2(new_n749_), .A3(new_n750_), .A4(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT117), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT117), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n683_), .A2(new_n754_), .A3(new_n687_), .A4(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT118), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n753_), .A2(KEYINPUT118), .A3(new_n755_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n748_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n747_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT119), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT119), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n763_), .B1(new_n747_), .B2(new_n760_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(G1336gat));
  INV_X1    g564(.A(new_n745_), .ZN(new_n766_));
  INV_X1    g565(.A(G92gat), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n766_), .A2(new_n767_), .A3(new_n407_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n411_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n768_), .B1(new_n769_), .B2(new_n767_), .ZN(G1337gat));
  NAND3_X1  g569(.A1(new_n766_), .A2(new_n493_), .A3(new_n652_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT120), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n756_), .A2(new_n652_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n773_), .B2(G99gat), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n480_), .B1(new_n753_), .B2(new_n755_), .ZN(new_n775_));
  INV_X1    g574(.A(G99gat), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n775_), .A2(KEYINPUT120), .A3(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n771_), .B1(new_n774_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT51), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n780_), .B(new_n771_), .C1(new_n774_), .C2(new_n777_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1338gat));
  NAND3_X1  g581(.A1(new_n766_), .A2(new_n494_), .A3(new_n413_), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n752_), .A2(new_n412_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n784_), .A2(new_n785_), .A3(G106gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n784_), .B2(G106gat), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n783_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g588(.A1(new_n622_), .A2(new_n600_), .A3(new_n624_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n582_), .A2(new_n586_), .A3(new_n583_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n588_), .A2(KEYINPUT55), .A3(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n586_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n597_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n792_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT56), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n792_), .A2(KEYINPUT56), .A3(new_n795_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n790_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n615_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n617_), .A2(new_n611_), .A3(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n609_), .B(new_n802_), .C1(new_n614_), .C2(new_n801_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n621_), .A2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n545_), .B1(new_n800_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n600_), .A2(new_n621_), .A3(new_n803_), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n792_), .A2(KEYINPUT56), .A3(new_n795_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT56), .B1(new_n792_), .B2(new_n795_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n809_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT58), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n809_), .B(KEYINPUT58), .C1(new_n810_), .C2(new_n811_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n814_), .A2(new_n636_), .A3(new_n638_), .A4(new_n815_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n545_), .B(KEYINPUT57), .C1(new_n800_), .C2(new_n805_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n808_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n577_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n640_), .B(new_n625_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT54), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n639_), .A2(new_n822_), .A3(new_n625_), .A4(new_n640_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n480_), .B1(new_n819_), .B2(new_n824_), .ZN(new_n825_));
  OR2_X1    g624(.A1(new_n482_), .A2(new_n483_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n425_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n825_), .A2(KEYINPUT59), .A3(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT59), .B1(new_n825_), .B2(new_n828_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(G113gat), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n832_), .A2(new_n833_), .A3(new_n625_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n819_), .A2(new_n824_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n835_), .A2(new_n652_), .A3(new_n828_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n833_), .B1(new_n836_), .B2(new_n625_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(KEYINPUT121), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n834_), .A2(new_n838_), .ZN(G1340gat));
  INV_X1    g638(.A(new_n836_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n605_), .A2(G120gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(KEYINPUT60), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n836_), .A2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n605_), .B1(new_n844_), .B2(new_n829_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n842_), .B1(new_n845_), .B2(KEYINPUT122), .ZN(new_n846_));
  OAI211_X1 g645(.A(KEYINPUT122), .B(new_n665_), .C1(new_n830_), .C2(new_n831_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(G120gat), .B1(new_n846_), .B2(new_n848_), .ZN(new_n849_));
  OR2_X1    g648(.A1(new_n842_), .A2(KEYINPUT60), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1341gat));
  INV_X1    g650(.A(G127gat), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n840_), .A2(new_n852_), .A3(new_n662_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n577_), .B1(new_n844_), .B2(new_n829_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n854_), .B2(new_n852_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT123), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1342gat));
  OAI21_X1  g656(.A(G134gat), .B1(new_n832_), .B2(new_n639_), .ZN(new_n858_));
  OR3_X1    g657(.A1(new_n836_), .A2(G134gat), .A3(new_n545_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(G1343gat));
  NAND2_X1  g659(.A1(new_n480_), .A2(new_n413_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n861_), .A2(new_n261_), .A3(new_n407_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n835_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n626_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT124), .B(G141gat), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1344gat));
  NAND2_X1  g665(.A1(new_n863_), .A2(new_n665_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g667(.A1(new_n863_), .A2(new_n662_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(KEYINPUT125), .ZN(new_n870_));
  XOR2_X1   g669(.A(KEYINPUT61), .B(G155gat), .Z(new_n871_));
  XNOR2_X1  g670(.A(new_n870_), .B(new_n871_), .ZN(G1346gat));
  INV_X1    g671(.A(G162gat), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n863_), .A2(new_n873_), .A3(new_n546_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n863_), .A2(new_n680_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(new_n873_), .ZN(G1347gat));
  INV_X1    g675(.A(KEYINPUT126), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n835_), .A2(new_n652_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n407_), .A2(new_n261_), .A3(new_n412_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n626_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n877_), .B1(new_n881_), .B2(G169gat), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n881_), .A2(new_n877_), .A3(G169gat), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n883_), .A2(KEYINPUT62), .A3(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT62), .ZN(new_n886_));
  INV_X1    g685(.A(new_n881_), .ZN(new_n887_));
  AOI22_X1  g686(.A1(new_n882_), .A2(new_n886_), .B1(new_n358_), .B2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n885_), .A2(new_n888_), .ZN(G1348gat));
  NAND2_X1  g688(.A1(new_n880_), .A2(new_n665_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g690(.A1(new_n880_), .A2(new_n662_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n375_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n893_), .B1(new_n337_), .B2(new_n892_), .ZN(G1350gat));
  OR2_X1    g693(.A1(new_n878_), .A2(new_n879_), .ZN(new_n895_));
  OAI21_X1  g694(.A(G190gat), .B1(new_n895_), .B2(new_n639_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n546_), .A2(new_n374_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(KEYINPUT127), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n896_), .B1(new_n895_), .B2(new_n898_), .ZN(G1351gat));
  NOR3_X1   g698(.A1(new_n861_), .A2(new_n425_), .A3(new_n411_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n835_), .A2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n626_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n665_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g704(.A1(new_n901_), .A2(new_n662_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n907_));
  AND2_X1   g706(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n906_), .A2(new_n907_), .A3(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n909_), .B1(new_n906_), .B2(new_n907_), .ZN(G1354gat));
  INV_X1    g709(.A(G218gat), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n901_), .A2(new_n911_), .A3(new_n546_), .ZN(new_n912_));
  AND2_X1   g711(.A1(new_n901_), .A2(new_n680_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n911_), .ZN(G1355gat));
endmodule


