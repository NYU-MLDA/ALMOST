//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 0 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n780_, new_n781_, new_n782_, new_n783_, new_n785_,
    new_n786_, new_n787_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n906_, new_n907_, new_n908_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n948_, new_n949_, new_n950_, new_n952_, new_n953_, new_n955_,
    new_n956_, new_n958_, new_n959_, new_n960_, new_n961_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n975_, new_n976_;
  XOR2_X1   g000(.A(G1gat), .B(G8gat), .Z(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  AND2_X1   g002(.A1(G15gat), .A2(G22gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G15gat), .A2(G22gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT14), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n207_), .B1(G1gat), .B2(G8gat), .ZN(new_n208_));
  NOR3_X1   g007(.A1(new_n206_), .A2(new_n208_), .A3(KEYINPUT75), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT75), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G15gat), .B(G22gat), .ZN(new_n211_));
  INV_X1    g010(.A(G1gat), .ZN(new_n212_));
  INV_X1    g011(.A(G8gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT14), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n210_), .B1(new_n211_), .B2(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n203_), .B1(new_n209_), .B2(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT75), .B1(new_n206_), .B2(new_n208_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n211_), .A2(new_n210_), .A3(new_n214_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(new_n202_), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(G36gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(G29gat), .ZN(new_n221_));
  INV_X1    g020(.A(G29gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(G36gat), .ZN(new_n223_));
  INV_X1    g022(.A(G50gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(G43gat), .ZN(new_n225_));
  INV_X1    g024(.A(G43gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(G50gat), .ZN(new_n227_));
  AND4_X1   g026(.A1(new_n221_), .A2(new_n223_), .A3(new_n225_), .A4(new_n227_), .ZN(new_n228_));
  AOI22_X1  g027(.A1(new_n221_), .A2(new_n223_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n216_), .A2(new_n219_), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT77), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n231_), .A2(new_n232_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n216_), .A2(new_n219_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n230_), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT76), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT76), .ZN(new_n238_));
  AOI211_X1 g037(.A(new_n238_), .B(new_n230_), .C1(new_n216_), .C2(new_n219_), .ZN(new_n239_));
  OAI22_X1  g038(.A1(new_n233_), .A2(new_n234_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G229gat), .A2(G233gat), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n230_), .A2(KEYINPUT15), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n230_), .A2(KEYINPUT15), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n244_), .A2(new_n245_), .A3(new_n219_), .A4(new_n216_), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n241_), .B(new_n246_), .C1(new_n237_), .C2(new_n239_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT78), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n219_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n202_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n236_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(new_n238_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n235_), .A2(KEYINPUT76), .A3(new_n236_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n255_), .A2(KEYINPUT78), .A3(new_n241_), .A4(new_n246_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n243_), .A2(new_n249_), .A3(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G169gat), .B(G197gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(G141gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT79), .B(G113gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n257_), .A2(new_n262_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n243_), .A2(new_n249_), .A3(new_n256_), .A4(new_n261_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT80), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  XOR2_X1   g066(.A(G155gat), .B(G162gat), .Z(new_n268_));
  OR2_X1    g067(.A1(G141gat), .A2(G148gat), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT2), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G141gat), .A2(G148gat), .ZN(new_n271_));
  AOI22_X1  g070(.A1(new_n269_), .A2(KEYINPUT3), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  OR3_X1    g071(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT89), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n268_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT1), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n268_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n279_), .A2(new_n269_), .A3(new_n271_), .A4(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n277_), .A2(new_n281_), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n282_), .A2(KEYINPUT29), .ZN(new_n283_));
  XOR2_X1   g082(.A(G22gat), .B(G50gat), .Z(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT28), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n283_), .B(new_n285_), .Z(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  OR2_X1    g086(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(G204gat), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT92), .ZN(new_n291_));
  INV_X1    g090(.A(G204gat), .ZN(new_n292_));
  AOI22_X1  g091(.A1(new_n290_), .A2(new_n291_), .B1(G197gat), .B2(new_n292_), .ZN(new_n293_));
  XOR2_X1   g092(.A(KEYINPUT90), .B(G197gat), .Z(new_n294_));
  NAND3_X1  g093(.A1(new_n294_), .A2(KEYINPUT92), .A3(G204gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT93), .B(KEYINPUT21), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n293_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT94), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT94), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n293_), .A2(new_n295_), .A3(new_n299_), .A4(new_n296_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  OR3_X1    g100(.A1(new_n292_), .A2(KEYINPUT91), .A3(G197gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT91), .B1(new_n292_), .B2(G197gat), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n302_), .B(new_n303_), .C1(new_n294_), .C2(G204gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT21), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G211gat), .B(G218gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n301_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n293_), .A2(new_n295_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n306_), .ZN(new_n311_));
  AND3_X1   g110(.A1(new_n310_), .A2(KEYINPUT21), .A3(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n309_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G228gat), .A2(G233gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n282_), .A2(KEYINPUT29), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n312_), .B1(new_n301_), .B2(new_n308_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n316_), .ZN(new_n319_));
  OAI211_X1 g118(.A(G228gat), .B(G233gat), .C1(new_n318_), .C2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G78gat), .B(G106gat), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n317_), .A2(new_n320_), .A3(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n322_), .B1(new_n317_), .B2(new_n320_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n287_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n317_), .A2(new_n320_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(new_n321_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n317_), .A2(new_n320_), .A3(new_n322_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n327_), .A2(new_n286_), .A3(new_n328_), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n325_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT30), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT22), .B(G169gat), .ZN(new_n332_));
  INV_X1    g131(.A(G176gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G169gat), .A2(G176gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  AND2_X1   g136(.A1(G183gat), .A2(G190gat), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT23), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n340_), .B1(new_n338_), .B2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(G183gat), .A2(G190gat), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n337_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  OR3_X1    g143(.A1(new_n341_), .A2(KEYINPUT84), .A3(new_n338_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n338_), .A2(new_n339_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT84), .B1(new_n341_), .B2(new_n338_), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n345_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(G169gat), .A2(G176gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT82), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(KEYINPUT24), .A3(new_n335_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT25), .B(G183gat), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT26), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT81), .B1(new_n354_), .B2(G190gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT26), .B(G190gat), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n353_), .B(new_n355_), .C1(new_n356_), .C2(KEYINPUT81), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n349_), .B(KEYINPUT82), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT24), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n352_), .A2(new_n357_), .A3(new_n360_), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n344_), .B(KEYINPUT85), .C1(new_n348_), .C2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n345_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n364_), .A2(new_n357_), .A3(new_n352_), .A4(new_n360_), .ZN(new_n365_));
  AOI21_X1  g164(.A(KEYINPUT85), .B1(new_n365_), .B2(new_n344_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n331_), .B1(new_n363_), .B2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n344_), .B1(new_n348_), .B2(new_n361_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT85), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(KEYINPUT30), .A3(new_n362_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G15gat), .B(G43gat), .ZN(new_n372_));
  AND3_X1   g171(.A1(new_n367_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n372_), .B1(new_n367_), .B2(new_n371_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G227gat), .A2(G233gat), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n375_), .B(KEYINPUT86), .Z(new_n376_));
  NOR3_X1   g175(.A1(new_n373_), .A2(new_n374_), .A3(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n376_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n372_), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n363_), .A2(new_n366_), .A3(new_n331_), .ZN(new_n380_));
  AOI21_X1  g179(.A(KEYINPUT30), .B1(new_n370_), .B2(new_n362_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n379_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n367_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n378_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G127gat), .B(G134gat), .ZN(new_n385_));
  XOR2_X1   g184(.A(G113gat), .B(G120gat), .Z(new_n386_));
  INV_X1    g185(.A(KEYINPUT87), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G113gat), .B(G120gat), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n389_), .A2(KEYINPUT87), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n385_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT88), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n386_), .A2(new_n387_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n389_), .A2(KEYINPUT87), .ZN(new_n394_));
  INV_X1    g193(.A(new_n385_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n393_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n391_), .A2(new_n392_), .A3(new_n396_), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n393_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT88), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT31), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G71gat), .B(G99gat), .ZN(new_n402_));
  XOR2_X1   g201(.A(new_n401_), .B(new_n402_), .Z(new_n403_));
  NOR3_X1   g202(.A1(new_n377_), .A2(new_n384_), .A3(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n401_), .B(new_n402_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n376_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n382_), .A2(new_n383_), .A3(new_n378_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n405_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n330_), .B1(new_n404_), .B2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n403_), .B1(new_n377_), .B2(new_n384_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n325_), .A2(new_n329_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n406_), .A2(new_n405_), .A3(new_n407_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n410_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n409_), .A2(new_n413_), .ZN(new_n414_));
  XOR2_X1   g213(.A(KEYINPUT97), .B(KEYINPUT18), .Z(new_n415_));
  XNOR2_X1  g214(.A(G8gat), .B(G36gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G64gat), .B(G92gat), .ZN(new_n418_));
  XOR2_X1   g217(.A(new_n417_), .B(new_n418_), .Z(new_n419_));
  NAND2_X1  g218(.A1(G226gat), .A2(G233gat), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n420_), .B(KEYINPUT95), .Z(new_n421_));
  XOR2_X1   g220(.A(new_n421_), .B(KEYINPUT19), .Z(new_n422_));
  INV_X1    g221(.A(KEYINPUT20), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n370_), .A2(new_n362_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n423_), .B1(new_n424_), .B2(new_n314_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n342_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n356_), .A2(new_n353_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n349_), .A2(new_n359_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n426_), .A2(new_n352_), .A3(new_n427_), .A4(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n343_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n336_), .B1(new_n364_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n318_), .A2(new_n429_), .A3(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n422_), .B1(new_n425_), .B2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n429_), .B1(new_n431_), .B2(KEYINPUT96), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT96), .ZN(new_n436_));
  AOI211_X1 g235(.A(new_n436_), .B(new_n336_), .C1(new_n364_), .C2(new_n430_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n307_), .B1(new_n298_), .B2(new_n300_), .ZN(new_n438_));
  OAI22_X1  g237(.A1(new_n435_), .A2(new_n437_), .B1(new_n438_), .B2(new_n312_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n318_), .A2(new_n370_), .A3(new_n362_), .ZN(new_n440_));
  AND4_X1   g239(.A1(KEYINPUT20), .A2(new_n439_), .A3(new_n440_), .A4(new_n422_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n419_), .B1(new_n434_), .B2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n439_), .A2(new_n440_), .A3(KEYINPUT20), .ZN(new_n443_));
  INV_X1    g242(.A(new_n422_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n435_), .A2(new_n437_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n444_), .B1(new_n446_), .B2(new_n318_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n425_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n419_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n445_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n442_), .A2(KEYINPUT27), .A3(new_n450_), .ZN(new_n451_));
  OR2_X1    g250(.A1(new_n451_), .A2(KEYINPUT100), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT27), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n445_), .A2(new_n448_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n419_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n450_), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n453_), .A2(new_n456_), .B1(new_n451_), .B2(KEYINPUT100), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G225gat), .A2(G233gat), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n400_), .A2(new_n282_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n395_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n398_), .A2(new_n461_), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n462_), .A2(new_n282_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n460_), .A2(new_n463_), .A3(KEYINPUT4), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT98), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT4), .ZN(new_n466_));
  AND4_X1   g265(.A1(new_n465_), .A2(new_n400_), .A3(new_n466_), .A4(new_n282_), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n397_), .A2(new_n399_), .B1(new_n277_), .B2(new_n281_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n465_), .B1(new_n468_), .B2(new_n466_), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n459_), .B(new_n464_), .C1(new_n467_), .C2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT99), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n460_), .A2(new_n463_), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n470_), .A2(new_n471_), .B1(new_n458_), .B2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n400_), .A2(new_n466_), .A3(new_n282_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT98), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n468_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n477_), .A2(KEYINPUT99), .A3(new_n459_), .A4(new_n464_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n473_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G1gat), .B(G29gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT0), .ZN(new_n481_));
  INV_X1    g280(.A(G57gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(G85gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n479_), .A2(new_n485_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n467_), .A2(new_n469_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n464_), .A2(new_n459_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n471_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n472_), .A2(new_n458_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n489_), .A2(new_n484_), .A3(new_n478_), .A4(new_n490_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n486_), .A2(new_n491_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n414_), .A2(new_n452_), .A3(new_n457_), .A4(new_n492_), .ZN(new_n493_));
  NOR3_X1   g292(.A1(new_n404_), .A2(new_n411_), .A3(new_n408_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT33), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n491_), .A2(new_n495_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n473_), .A2(KEYINPUT33), .A3(new_n484_), .A4(new_n478_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n484_), .B1(new_n472_), .B2(new_n459_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n464_), .A2(new_n458_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n499_), .B1(new_n500_), .B2(new_n487_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n455_), .A2(new_n450_), .A3(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n498_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n449_), .A2(KEYINPUT32), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n445_), .A2(new_n448_), .A3(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n434_), .A2(new_n441_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n505_), .B1(new_n506_), .B2(new_n504_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n507_), .B1(new_n486_), .B2(new_n491_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n494_), .B1(new_n503_), .B2(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n267_), .B1(new_n493_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT12), .ZN(new_n511_));
  XOR2_X1   g310(.A(G85gat), .B(G92gat), .Z(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NOR3_X1   g314(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n517_));
  NOR3_X1   g316(.A1(new_n515_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT66), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(KEYINPUT66), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n513_), .B1(new_n518_), .B2(new_n523_), .ZN(new_n524_));
  AND2_X1   g323(.A1(KEYINPUT68), .A2(KEYINPUT8), .ZN(new_n525_));
  OR2_X1    g324(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n526_));
  INV_X1    g325(.A(G106gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n526_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT64), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n515_), .A2(new_n517_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n526_), .A2(KEYINPUT64), .A3(new_n527_), .A4(new_n528_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G85gat), .A2(G92gat), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT9), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT65), .B(G92gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(G85gat), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n537_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  OAI22_X1  g340(.A1(new_n524_), .A2(new_n525_), .B1(new_n534_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT67), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n543_), .B1(new_n512_), .B2(new_n525_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n521_), .A2(new_n522_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G99gat), .A2(G106gat), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT6), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(G99gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(new_n527_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n548_), .B(new_n514_), .C1(new_n550_), .C2(KEYINPUT7), .ZN(new_n551_));
  OAI21_X1  g350(.A(KEYINPUT67), .B1(new_n545_), .B2(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n544_), .B1(new_n552_), .B2(KEYINPUT8), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n542_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT69), .ZN(new_n555_));
  INV_X1    g354(.A(G64gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(G57gat), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n482_), .A2(G64gat), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n557_), .A2(new_n558_), .A3(KEYINPUT11), .ZN(new_n559_));
  AOI21_X1  g358(.A(KEYINPUT11), .B1(new_n557_), .B2(new_n558_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G71gat), .B(G78gat), .ZN(new_n561_));
  NOR3_X1   g360(.A1(new_n559_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G57gat), .B(G64gat), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n563_), .A2(new_n561_), .A3(KEYINPUT11), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n555_), .B1(new_n562_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n560_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n563_), .A2(KEYINPUT11), .ZN(new_n568_));
  INV_X1    g367(.A(new_n561_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n567_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(KEYINPUT69), .A3(new_n564_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n566_), .A2(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n511_), .B1(new_n554_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(G230gat), .ZN(new_n574_));
  INV_X1    g373(.A(G233gat), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n576_), .B1(new_n554_), .B2(new_n572_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n562_), .A2(new_n565_), .ZN(new_n578_));
  OAI211_X1 g377(.A(KEYINPUT12), .B(new_n578_), .C1(new_n542_), .C2(new_n553_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n573_), .A2(new_n577_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n576_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n544_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n543_), .B1(new_n518_), .B2(new_n523_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT8), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n583_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n541_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n512_), .B1(new_n545_), .B2(new_n551_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n525_), .ZN(new_n590_));
  AOI22_X1  g389(.A1(new_n587_), .A2(new_n588_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n572_), .B1(new_n586_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n554_), .A2(new_n572_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n582_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n581_), .A2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G120gat), .B(G148gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(new_n292_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT5), .B(G176gat), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n598_), .B(new_n599_), .Z(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT70), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n596_), .B(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT13), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G127gat), .B(G155gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT16), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(G183gat), .ZN(new_n607_));
  INV_X1    g406(.A(G211gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT17), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n235_), .B(new_n612_), .Z(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n611_), .B1(new_n572_), .B2(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n615_), .B1(new_n572_), .B2(new_n614_), .ZN(new_n616_));
  AOI211_X1 g415(.A(new_n610_), .B(new_n609_), .C1(new_n614_), .C2(new_n578_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n617_), .B1(new_n578_), .B2(new_n614_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G232gat), .A2(G233gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT71), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT34), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT35), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n623_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n591_), .A2(new_n586_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n625_), .B1(new_n626_), .B2(new_n230_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n244_), .A2(new_n245_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n554_), .A2(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n624_), .B1(new_n627_), .B2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G190gat), .B(G218gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G134gat), .B(G162gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n633_), .A2(KEYINPUT36), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n626_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n624_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n554_), .A2(new_n236_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n635_), .A2(new_n636_), .A3(new_n625_), .A4(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n630_), .A2(new_n634_), .A3(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT72), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n630_), .A2(new_n638_), .A3(KEYINPUT72), .A4(new_n634_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n630_), .A2(new_n638_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n633_), .B(KEYINPUT36), .Z(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  XOR2_X1   g445(.A(KEYINPUT73), .B(KEYINPUT37), .Z(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n643_), .A2(new_n646_), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT74), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n643_), .A2(new_n646_), .ZN(new_n651_));
  AOI22_X1  g450(.A1(new_n649_), .A2(new_n650_), .B1(new_n651_), .B2(KEYINPUT37), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n643_), .A2(KEYINPUT74), .A3(new_n646_), .A4(new_n648_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  AND4_X1   g453(.A1(new_n510_), .A2(new_n604_), .A3(new_n619_), .A4(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n492_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(new_n212_), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT38), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n619_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n651_), .ZN(new_n661_));
  AOI211_X1 g460(.A(new_n660_), .B(new_n661_), .C1(new_n493_), .C2(new_n509_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n604_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n265_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n662_), .A2(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(G1gat), .B1(new_n666_), .B2(new_n492_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n657_), .A2(new_n658_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n659_), .A2(new_n667_), .A3(new_n668_), .ZN(G1324gat));
  NAND2_X1  g468(.A1(new_n457_), .A2(new_n452_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n655_), .A2(new_n213_), .A3(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n670_), .ZN(new_n672_));
  OAI21_X1  g471(.A(G8gat), .B1(new_n666_), .B2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT101), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT39), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT101), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n676_), .B(G8gat), .C1(new_n666_), .C2(new_n672_), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n674_), .A2(new_n675_), .A3(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n675_), .B1(new_n674_), .B2(new_n677_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n671_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT40), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  OAI211_X1 g481(.A(KEYINPUT40), .B(new_n671_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1325gat));
  NOR2_X1   g483(.A1(new_n404_), .A2(new_n408_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G15gat), .B1(new_n666_), .B2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT102), .B(KEYINPUT41), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n687_), .ZN(new_n689_));
  INV_X1    g488(.A(G15gat), .ZN(new_n690_));
  INV_X1    g489(.A(new_n685_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n655_), .A2(new_n690_), .A3(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n688_), .A2(new_n689_), .A3(new_n692_), .ZN(G1326gat));
  OAI21_X1  g492(.A(G22gat), .B1(new_n666_), .B2(new_n330_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT42), .ZN(new_n695_));
  INV_X1    g494(.A(G22gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n655_), .A2(new_n696_), .A3(new_n411_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(G1327gat));
  AND4_X1   g497(.A1(new_n510_), .A2(new_n604_), .A3(new_n660_), .A4(new_n661_), .ZN(new_n699_));
  AOI21_X1  g498(.A(G29gat), .B1(new_n699_), .B2(new_n656_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n652_), .A2(new_n702_), .A3(new_n653_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n493_), .B2(new_n509_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT103), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n649_), .A2(new_n650_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n651_), .A2(KEYINPUT37), .ZN(new_n708_));
  AND4_X1   g507(.A1(new_n705_), .A2(new_n707_), .A3(new_n653_), .A4(new_n708_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n706_), .A2(new_n709_), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n410_), .A2(new_n412_), .A3(new_n411_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n411_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n492_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n509_), .B1(new_n713_), .B2(new_n670_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n710_), .A2(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n704_), .B1(new_n715_), .B2(KEYINPUT43), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n665_), .A2(new_n660_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n701_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n717_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n702_), .B1(new_n710_), .B2(new_n714_), .ZN(new_n720_));
  OAI211_X1 g519(.A(KEYINPUT44), .B(new_n719_), .C1(new_n720_), .C2(new_n704_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n718_), .A2(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n492_), .A2(new_n222_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n700_), .B1(new_n722_), .B2(new_n723_), .ZN(G1328gat));
  NAND3_X1  g523(.A1(new_n699_), .A2(new_n220_), .A3(new_n670_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT45), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n718_), .A2(new_n670_), .A3(new_n721_), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n727_), .A2(KEYINPUT104), .A3(G36gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT104), .B1(new_n727_), .B2(G36gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n726_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n731_), .B(new_n726_), .C1(new_n728_), .C2(new_n729_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1329gat));
  NOR2_X1   g534(.A1(new_n685_), .A2(new_n226_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n718_), .A2(new_n721_), .A3(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT106), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT106), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n718_), .A2(new_n739_), .A3(new_n721_), .A4(new_n736_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n699_), .A2(new_n691_), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n738_), .B(new_n740_), .C1(G43gat), .C2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g542(.A(G50gat), .B1(new_n699_), .B2(new_n411_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n330_), .A2(new_n224_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n722_), .B2(new_n745_), .ZN(G1331gat));
  NOR2_X1   g545(.A1(new_n604_), .A2(new_n265_), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n747_), .A2(new_n619_), .A3(new_n654_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(new_n714_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n750_), .A2(new_n482_), .A3(new_n656_), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n662_), .A2(new_n267_), .A3(new_n663_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n752_), .A2(new_n656_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n751_), .B1(new_n753_), .B2(new_n482_), .ZN(G1332gat));
  AOI21_X1  g553(.A(new_n556_), .B1(new_n752_), .B2(new_n670_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT48), .Z(new_n756_));
  NAND2_X1  g555(.A1(new_n670_), .A2(new_n556_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT107), .Z(new_n758_));
  OAI21_X1  g557(.A(new_n756_), .B1(new_n749_), .B2(new_n758_), .ZN(G1333gat));
  INV_X1    g558(.A(G71gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n752_), .B2(new_n691_), .ZN(new_n761_));
  XOR2_X1   g560(.A(new_n761_), .B(KEYINPUT49), .Z(new_n762_));
  NAND3_X1  g561(.A1(new_n750_), .A2(new_n760_), .A3(new_n691_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1334gat));
  INV_X1    g563(.A(G78gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n752_), .B2(new_n411_), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT50), .Z(new_n767_));
  NAND3_X1  g566(.A1(new_n750_), .A2(new_n765_), .A3(new_n411_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(G1335gat));
  INV_X1    g568(.A(new_n716_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n747_), .A2(new_n660_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT109), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(G85gat), .B1(new_n773_), .B2(new_n492_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n714_), .A2(new_n660_), .A3(new_n661_), .A4(new_n747_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT108), .ZN(new_n776_));
  INV_X1    g575(.A(G85gat), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(new_n777_), .A3(new_n656_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n774_), .A2(new_n778_), .ZN(G1336gat));
  AOI21_X1  g578(.A(G92gat), .B1(new_n776_), .B2(new_n670_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n773_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n670_), .A2(new_n538_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT110), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n780_), .B1(new_n781_), .B2(new_n783_), .ZN(G1337gat));
  NAND4_X1  g583(.A1(new_n776_), .A2(new_n691_), .A3(new_n526_), .A4(new_n528_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n773_), .A2(new_n685_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n785_), .B1(new_n786_), .B2(new_n549_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g587(.A1(new_n776_), .A2(new_n527_), .A3(new_n411_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n770_), .A2(new_n411_), .A3(new_n772_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n790_), .A2(new_n791_), .A3(G106gat), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n790_), .B2(G106gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n789_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n580_), .A2(new_n796_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n594_), .B(new_n579_), .C1(new_n592_), .C2(KEYINPUT12), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n576_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n573_), .A2(new_n577_), .A3(KEYINPUT55), .A4(new_n579_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n797_), .A2(new_n799_), .A3(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT113), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT56), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n600_), .A2(new_n803_), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n801_), .A2(new_n802_), .A3(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT56), .B1(new_n801_), .B2(new_n601_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n802_), .B1(new_n801_), .B2(new_n804_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n805_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n596_), .A2(new_n600_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n265_), .A2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT114), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n812_));
  INV_X1    g611(.A(new_n810_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n807_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n801_), .A2(new_n601_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n803_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n816_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n812_), .B(new_n813_), .C1(new_n817_), .C2(new_n805_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n240_), .A2(new_n241_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n255_), .A2(new_n242_), .A3(new_n246_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n262_), .A3(new_n821_), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n264_), .A2(new_n819_), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n819_), .B1(new_n264_), .B2(new_n822_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n603_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n811_), .A2(new_n818_), .A3(new_n825_), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n826_), .A2(KEYINPUT57), .A3(new_n651_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT57), .B1(new_n826_), .B2(new_n651_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n654_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n801_), .A2(new_n804_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT116), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT116), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n801_), .A2(new_n833_), .A3(new_n804_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n816_), .A2(new_n832_), .A3(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n824_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n264_), .A2(new_n819_), .A3(new_n822_), .ZN(new_n837_));
  AOI22_X1  g636(.A1(new_n836_), .A2(new_n837_), .B1(new_n596_), .B2(new_n600_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n835_), .A2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT58), .B1(new_n839_), .B2(KEYINPUT117), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842_));
  AOI211_X1 g641(.A(new_n841_), .B(new_n842_), .C1(new_n835_), .C2(new_n838_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n830_), .B1(new_n840_), .B2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n829_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n660_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n654_), .A2(new_n267_), .A3(new_n604_), .A4(new_n619_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  XOR2_X1   g647(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(KEYINPUT112), .A3(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT112), .ZN(new_n851_));
  INV_X1    g650(.A(new_n849_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n847_), .B2(new_n852_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n850_), .B(new_n853_), .C1(new_n848_), .C2(new_n849_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n846_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n656_), .A2(new_n712_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n670_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n855_), .A2(new_n856_), .A3(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n266_), .A2(G113gat), .ZN(new_n860_));
  XOR2_X1   g659(.A(new_n860_), .B(KEYINPUT120), .Z(new_n861_));
  INV_X1    g660(.A(new_n858_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n844_), .A2(KEYINPUT118), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n826_), .A2(new_n651_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n826_), .A2(KEYINPUT57), .A3(new_n651_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n809_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n833_), .B1(new_n801_), .B2(new_n804_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n806_), .A2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n868_), .B1(new_n870_), .B2(new_n834_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n842_), .B1(new_n871_), .B2(new_n841_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n839_), .A2(KEYINPUT117), .A3(KEYINPUT58), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n874_), .A2(new_n875_), .A3(new_n830_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n863_), .A2(new_n866_), .A3(new_n867_), .A4(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT119), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n875_), .B1(new_n874_), .B2(new_n830_), .ZN(new_n879_));
  AOI211_X1 g678(.A(KEYINPUT118), .B(new_n654_), .C1(new_n872_), .C2(new_n873_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n881_), .A2(new_n882_), .A3(new_n829_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n878_), .A2(new_n883_), .A3(new_n660_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n862_), .B1(new_n884_), .B2(new_n854_), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n859_), .B(new_n861_), .C1(new_n885_), .C2(new_n856_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(G113gat), .B1(new_n885_), .B2(new_n265_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1340gat));
  OAI211_X1 g688(.A(new_n663_), .B(new_n859_), .C1(new_n885_), .C2(new_n856_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(G120gat), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT60), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n892_), .B1(new_n604_), .B2(G120gat), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n885_), .B(new_n893_), .C1(new_n892_), .C2(G120gat), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n891_), .A2(new_n894_), .ZN(G1341gat));
  OAI211_X1 g694(.A(new_n619_), .B(new_n859_), .C1(new_n885_), .C2(new_n856_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(G127gat), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n884_), .A2(new_n854_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n858_), .ZN(new_n899_));
  OR3_X1    g698(.A1(new_n899_), .A2(G127gat), .A3(new_n660_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n897_), .A2(new_n900_), .ZN(G1342gat));
  OAI211_X1 g700(.A(new_n830_), .B(new_n859_), .C1(new_n885_), .C2(new_n856_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(G134gat), .ZN(new_n903_));
  OR3_X1    g702(.A1(new_n899_), .A2(G134gat), .A3(new_n651_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1343gat));
  NOR3_X1   g704(.A1(new_n670_), .A2(new_n492_), .A3(new_n413_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n898_), .A2(new_n265_), .A3(new_n906_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(KEYINPUT121), .B(G141gat), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n907_), .B(new_n908_), .ZN(G1344gat));
  NAND3_X1  g708(.A1(new_n898_), .A2(new_n663_), .A3(new_n906_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(KEYINPUT122), .B(G148gat), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n910_), .B(new_n911_), .ZN(G1345gat));
  NAND3_X1  g711(.A1(new_n898_), .A2(new_n619_), .A3(new_n906_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(KEYINPUT61), .B(G155gat), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n913_), .B(new_n914_), .ZN(G1346gat));
  AND4_X1   g714(.A1(G162gat), .A2(new_n898_), .A3(new_n710_), .A4(new_n906_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n906_), .ZN(new_n917_));
  AOI211_X1 g716(.A(new_n651_), .B(new_n917_), .C1(new_n884_), .C2(new_n854_), .ZN(new_n918_));
  OAI21_X1  g717(.A(KEYINPUT123), .B1(new_n918_), .B2(G162gat), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n898_), .A2(new_n661_), .A3(new_n906_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n921_));
  INV_X1    g720(.A(G162gat), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n920_), .A2(new_n921_), .A3(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n916_), .B1(new_n919_), .B2(new_n923_), .ZN(G1347gat));
  XOR2_X1   g723(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n925_));
  INV_X1    g724(.A(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n670_), .A2(new_n492_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n927_), .A2(new_n685_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n330_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n929_), .B1(new_n846_), .B2(new_n854_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n930_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n931_), .A2(new_n664_), .ZN(new_n932_));
  INV_X1    g731(.A(G169gat), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n926_), .B1(new_n932_), .B2(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n932_), .A2(new_n332_), .ZN(new_n935_));
  OAI211_X1 g734(.A(G169gat), .B(new_n925_), .C1(new_n931_), .C2(new_n664_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n934_), .A2(new_n935_), .A3(new_n936_), .ZN(G1348gat));
  NOR4_X1   g736(.A1(new_n927_), .A2(new_n333_), .A3(new_n685_), .A4(new_n604_), .ZN(new_n938_));
  AND3_X1   g737(.A1(new_n898_), .A2(new_n330_), .A3(new_n938_), .ZN(new_n939_));
  AOI21_X1  g738(.A(G176gat), .B1(new_n930_), .B2(new_n663_), .ZN(new_n940_));
  OAI21_X1  g739(.A(KEYINPUT125), .B1(new_n939_), .B2(new_n940_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n940_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n411_), .B1(new_n884_), .B2(new_n854_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(new_n938_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n942_), .A2(new_n944_), .A3(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n941_), .A2(new_n946_), .ZN(G1349gat));
  NOR3_X1   g746(.A1(new_n931_), .A2(new_n353_), .A3(new_n660_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n943_), .A2(new_n619_), .A3(new_n928_), .ZN(new_n949_));
  INV_X1    g748(.A(G183gat), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n948_), .B1(new_n949_), .B2(new_n950_), .ZN(G1350gat));
  OAI21_X1  g750(.A(G190gat), .B1(new_n931_), .B2(new_n654_), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n930_), .A2(new_n356_), .A3(new_n661_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n952_), .A2(new_n953_), .ZN(G1351gat));
  NOR2_X1   g753(.A1(new_n927_), .A2(new_n413_), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n898_), .A2(new_n265_), .A3(new_n955_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n956_), .B(G197gat), .ZN(G1352gat));
  AND2_X1   g756(.A1(new_n898_), .A2(new_n955_), .ZN(new_n958_));
  AOI21_X1  g757(.A(G204gat), .B1(new_n958_), .B2(new_n663_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n898_), .A2(new_n955_), .ZN(new_n960_));
  NOR3_X1   g759(.A1(new_n960_), .A2(new_n292_), .A3(new_n604_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n959_), .A2(new_n961_), .ZN(G1353gat));
  INV_X1    g761(.A(KEYINPUT63), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n963_), .A2(new_n608_), .A3(KEYINPUT126), .ZN(new_n964_));
  XOR2_X1   g763(.A(new_n964_), .B(KEYINPUT127), .Z(new_n965_));
  INV_X1    g764(.A(new_n965_), .ZN(new_n966_));
  AOI21_X1  g765(.A(new_n660_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n967_));
  AND3_X1   g766(.A1(new_n898_), .A2(new_n955_), .A3(new_n967_), .ZN(new_n968_));
  AOI21_X1  g767(.A(KEYINPUT126), .B1(new_n963_), .B2(new_n608_), .ZN(new_n969_));
  OAI21_X1  g768(.A(new_n966_), .B1(new_n968_), .B2(new_n969_), .ZN(new_n970_));
  INV_X1    g769(.A(new_n969_), .ZN(new_n971_));
  INV_X1    g770(.A(new_n967_), .ZN(new_n972_));
  OAI211_X1 g771(.A(new_n965_), .B(new_n971_), .C1(new_n960_), .C2(new_n972_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n970_), .A2(new_n973_), .ZN(G1354gat));
  OR3_X1    g773(.A1(new_n960_), .A2(G218gat), .A3(new_n651_), .ZN(new_n975_));
  OAI21_X1  g774(.A(G218gat), .B1(new_n960_), .B2(new_n654_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n975_), .A2(new_n976_), .ZN(G1355gat));
endmodule


