//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1 1 0 1 0 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n952_, new_n953_, new_n954_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n965_, new_n966_;
  XNOR2_X1  g000(.A(G127gat), .B(G155gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G211gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT16), .B(G183gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  AND2_X1   g004(.A1(new_n205_), .A2(KEYINPUT17), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(KEYINPUT17), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  OR2_X1    g007(.A1(KEYINPUT69), .A2(G15gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(KEYINPUT69), .A2(G15gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(G22gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G1gat), .ZN(new_n214_));
  INV_X1    g013(.A(G8gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT14), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n209_), .A2(G22gat), .A3(new_n210_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n213_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  XOR2_X1   g017(.A(G1gat), .B(G8gat), .Z(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n213_), .A2(new_n219_), .A3(new_n216_), .A4(new_n217_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G231gat), .A2(G233gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n223_), .B(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G71gat), .B(G78gat), .ZN(new_n226_));
  OR2_X1    g025(.A1(G57gat), .A2(G64gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G57gat), .A2(G64gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT11), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT11), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n227_), .A2(new_n231_), .A3(new_n228_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n226_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n226_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n234_), .B1(KEYINPUT11), .B2(new_n229_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n225_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n236_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n223_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n239_), .A2(new_n224_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n223_), .B1(G231gat), .B2(G233gat), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n238_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT71), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n237_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n243_), .B1(new_n237_), .B2(new_n242_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n208_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT72), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  OAI211_X1 g047(.A(KEYINPUT72), .B(new_n208_), .C1(new_n244_), .C2(new_n245_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT73), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n237_), .A2(new_n242_), .A3(new_n206_), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n252_), .B(KEYINPUT70), .Z(new_n253_));
  AND3_X1   g052(.A1(new_n250_), .A2(new_n251_), .A3(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n251_), .B1(new_n250_), .B2(new_n253_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(G85gat), .B(G92gat), .Z(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT9), .ZN(new_n258_));
  XOR2_X1   g057(.A(KEYINPUT10), .B(G99gat), .Z(new_n259_));
  INV_X1    g058(.A(G106gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT9), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n262_), .A2(G85gat), .A3(G92gat), .ZN(new_n263_));
  AND3_X1   g062(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n264_));
  AOI21_X1  g063(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n258_), .A2(new_n261_), .A3(new_n263_), .A4(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT8), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NOR3_X1   g069(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT64), .B1(new_n264_), .B2(new_n265_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G99gat), .A2(G106gat), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT6), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT64), .ZN(new_n277_));
  NAND3_X1  g076(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n276_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n272_), .A2(new_n273_), .A3(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n268_), .B1(new_n280_), .B2(new_n257_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n257_), .A2(new_n268_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n282_), .B1(new_n266_), .B2(new_n272_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n267_), .B1(new_n281_), .B2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT65), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT65), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n286_), .B(new_n267_), .C1(new_n281_), .C2(new_n283_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G29gat), .B(G36gat), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G43gat), .B(G50gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(G43gat), .B(G50gat), .Z(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n289_), .ZN(new_n294_));
  AND3_X1   g093(.A1(new_n292_), .A2(new_n294_), .A3(KEYINPUT15), .ZN(new_n295_));
  AOI21_X1  g094(.A(KEYINPUT15), .B1(new_n292_), .B2(new_n294_), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n288_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G232gat), .A2(G233gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT34), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT35), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n292_), .A2(new_n294_), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n304_), .B(new_n267_), .C1(new_n281_), .C2(new_n283_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n298_), .A2(new_n303_), .A3(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n301_), .A2(new_n302_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n307_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n298_), .A2(new_n309_), .A3(new_n303_), .A4(new_n305_), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G190gat), .B(G218gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G134gat), .B(G162gat), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n312_), .B(new_n313_), .Z(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT36), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n311_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n314_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT67), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n318_), .B1(new_n319_), .B2(KEYINPUT36), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n319_), .A2(KEYINPUT36), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n308_), .A2(new_n320_), .A3(new_n321_), .A4(new_n310_), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n322_), .A2(KEYINPUT68), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(KEYINPUT68), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n317_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT37), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n238_), .A2(KEYINPUT12), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n236_), .B(new_n267_), .C1(new_n281_), .C2(new_n283_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT12), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n284_), .A2(new_n238_), .ZN(new_n331_));
  AOI22_X1  g130(.A1(new_n288_), .A2(new_n328_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G230gat), .A2(G233gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n331_), .A2(new_n329_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(G230gat), .A3(G233gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  XOR2_X1   g136(.A(G176gat), .B(G204gat), .Z(new_n338_));
  XNOR2_X1  g137(.A(G120gat), .B(G148gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT66), .B(KEYINPUT5), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n337_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n342_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n334_), .A2(new_n336_), .A3(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT13), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n317_), .B(KEYINPUT37), .C1(new_n323_), .C2(new_n324_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n256_), .A2(new_n327_), .A3(new_n347_), .A4(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G226gat), .A2(G233gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT19), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT80), .ZN(new_n353_));
  NOR2_X1   g152(.A1(KEYINPUT79), .A2(G176gat), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(KEYINPUT79), .A2(G176gat), .ZN(new_n356_));
  OR2_X1    g155(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n358_));
  AOI22_X1  g157(.A1(new_n355_), .A2(new_n356_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n353_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n356_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n358_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n365_));
  OAI22_X1  g164(.A1(new_n354_), .A2(new_n363_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n366_), .A2(KEYINPUT80), .A3(new_n360_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G183gat), .A2(G190gat), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT23), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n370_), .B(new_n371_), .C1(G183gat), .C2(G190gat), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n362_), .A2(new_n367_), .A3(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT25), .B(G183gat), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT77), .ZN(new_n375_));
  INV_X1    g174(.A(G190gat), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT26), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  OR2_X1    g176(.A1(new_n376_), .A2(KEYINPUT26), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n374_), .B(new_n377_), .C1(new_n378_), .C2(new_n375_), .ZN(new_n379_));
  INV_X1    g178(.A(G169gat), .ZN(new_n380_));
  INV_X1    g179(.A(G176gat), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n380_), .A2(new_n381_), .A3(KEYINPUT78), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT78), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n383_), .B1(G169gat), .B2(G176gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT24), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n370_), .A2(new_n371_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n382_), .A2(new_n384_), .A3(KEYINPUT24), .A4(new_n360_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n379_), .A2(new_n387_), .A3(new_n389_), .A4(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n373_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT81), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT81), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n373_), .A2(new_n394_), .A3(new_n391_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G211gat), .B(G218gat), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT88), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  OR2_X1    g197(.A1(G211gat), .A2(G218gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G211gat), .A2(G218gat), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n399_), .A2(KEYINPUT88), .A3(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n398_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G197gat), .A2(G204gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT86), .B(G204gat), .ZN(new_n404_));
  OAI211_X1 g203(.A(KEYINPUT21), .B(new_n403_), .C1(new_n404_), .C2(G197gat), .ZN(new_n405_));
  INV_X1    g204(.A(G204gat), .ZN(new_n406_));
  OR3_X1    g205(.A1(new_n406_), .A2(KEYINPUT87), .A3(G197gat), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT87), .B1(new_n406_), .B2(G197gat), .ZN(new_n408_));
  INV_X1    g207(.A(G197gat), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n407_), .B(new_n408_), .C1(new_n404_), .C2(new_n409_), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n402_), .B(new_n405_), .C1(new_n410_), .C2(KEYINPUT21), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n410_), .A2(KEYINPUT21), .A3(new_n398_), .A4(new_n401_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n393_), .A2(new_n395_), .A3(new_n414_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n415_), .A2(KEYINPUT20), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT26), .B(G190gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n374_), .A2(new_n417_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n387_), .A2(new_n418_), .A3(new_n389_), .A4(new_n390_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n366_), .A2(new_n372_), .A3(new_n360_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n413_), .A2(KEYINPUT91), .A3(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(KEYINPUT91), .B1(new_n413_), .B2(new_n421_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n352_), .B1(new_n416_), .B2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n414_), .B1(new_n393_), .B2(new_n395_), .ZN(new_n427_));
  OAI211_X1 g226(.A(KEYINPUT20), .B(new_n352_), .C1(new_n413_), .C2(new_n421_), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT92), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n373_), .A2(new_n394_), .A3(new_n391_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n394_), .B1(new_n373_), .B2(new_n391_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n413_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n428_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT92), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n432_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n429_), .A2(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(G8gat), .B(G36gat), .Z(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(G92gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT18), .B(G64gat), .ZN(new_n439_));
  XOR2_X1   g238(.A(new_n438_), .B(new_n439_), .Z(new_n440_));
  NOR3_X1   g239(.A1(new_n426_), .A2(new_n436_), .A3(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT20), .B1(new_n413_), .B2(new_n421_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT97), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  OAI211_X1 g243(.A(KEYINPUT97), .B(KEYINPUT20), .C1(new_n413_), .C2(new_n421_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n432_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n351_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT98), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n416_), .A2(new_n352_), .A3(new_n425_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT98), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n446_), .A2(new_n450_), .A3(new_n351_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n448_), .A2(new_n449_), .A3(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n441_), .B1(new_n440_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT27), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n440_), .B1(new_n426_), .B2(new_n436_), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n429_), .A2(new_n435_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n440_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n415_), .A2(KEYINPUT20), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n351_), .B1(new_n458_), .B2(new_n424_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n456_), .A2(new_n457_), .A3(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(KEYINPUT27), .B1(new_n455_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n454_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(G155gat), .ZN(new_n464_));
  INV_X1    g263(.A(G162gat), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT1), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT1), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n467_), .A2(G155gat), .A3(G162gat), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n466_), .B(new_n468_), .C1(G155gat), .C2(G162gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G141gat), .A2(G148gat), .ZN(new_n470_));
  INV_X1    g269(.A(G141gat), .ZN(new_n471_));
  INV_X1    g270(.A(G148gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n469_), .A2(new_n470_), .A3(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G155gat), .B(G162gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT83), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT3), .ZN(new_n480_));
  OAI211_X1 g279(.A(new_n479_), .B(new_n480_), .C1(G141gat), .C2(G148gat), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n471_), .B(new_n472_), .C1(KEYINPUT83), .C2(KEYINPUT3), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n478_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT2), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n470_), .A2(new_n484_), .ZN(new_n485_));
  AOI211_X1 g284(.A(KEYINPUT84), .B(new_n475_), .C1(new_n483_), .C2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT84), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n481_), .A2(new_n482_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n478_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(new_n485_), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n475_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n487_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n474_), .B1(new_n486_), .B2(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(G22gat), .B(G50gat), .Z(new_n494_));
  OR3_X1    g293(.A1(new_n493_), .A2(KEYINPUT29), .A3(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n494_), .B1(new_n493_), .B2(KEYINPUT29), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n496_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(G78gat), .B(G106gat), .Z(new_n502_));
  INV_X1    g301(.A(new_n474_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n490_), .A2(new_n491_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT84), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n490_), .A2(new_n487_), .A3(new_n491_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n503_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT29), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n413_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G228gat), .A2(G233gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n413_), .B(new_n510_), .C1(new_n507_), .C2(new_n508_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n502_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n501_), .A2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n512_), .A2(new_n513_), .A3(new_n502_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT89), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n512_), .A2(new_n513_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n502_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n519_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n520_), .A2(new_n518_), .A3(new_n521_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT90), .B1(new_n525_), .B2(new_n501_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT90), .ZN(new_n527_));
  AOI211_X1 g326(.A(new_n527_), .B(new_n500_), .C1(new_n523_), .C2(new_n524_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n517_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT93), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G127gat), .B(G134gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G113gat), .B(G120gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n493_), .A2(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n530_), .B1(new_n535_), .B2(KEYINPUT4), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n533_), .B(new_n474_), .C1(new_n486_), .C2(new_n492_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n535_), .A2(KEYINPUT4), .A3(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G225gat), .A2(G233gat), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT4), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n493_), .A2(KEYINPUT93), .A3(new_n541_), .A4(new_n534_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n536_), .A2(new_n538_), .A3(new_n540_), .A4(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n535_), .A2(new_n539_), .A3(new_n537_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G1gat), .B(G29gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(G85gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT0), .B(G57gat), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n547_), .B(new_n548_), .Z(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n545_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n543_), .A2(new_n544_), .A3(new_n549_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n393_), .A2(new_n395_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G15gat), .B(G43gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT31), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n555_), .B(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G71gat), .B(G99gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT82), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(new_n533_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G227gat), .A2(G233gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT30), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n561_), .B(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n558_), .B(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n554_), .A2(new_n565_), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n463_), .A2(new_n529_), .A3(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n461_), .B1(new_n453_), .B2(KEYINPUT27), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n529_), .A2(new_n568_), .A3(new_n554_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n457_), .A2(KEYINPUT32), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n456_), .A2(new_n570_), .A3(new_n459_), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n448_), .A2(new_n449_), .A3(new_n451_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n553_), .B(new_n571_), .C1(new_n572_), .C2(new_n570_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT95), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n505_), .A2(new_n506_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n533_), .B1(new_n575_), .B2(new_n474_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n537_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n574_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n535_), .A2(KEYINPUT95), .A3(new_n537_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n578_), .A2(new_n540_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n550_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT96), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n536_), .A2(new_n538_), .A3(new_n539_), .A4(new_n542_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n580_), .A2(KEYINPUT96), .A3(new_n550_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n583_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT33), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n552_), .A2(new_n587_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n586_), .A2(new_n588_), .A3(new_n460_), .A4(new_n455_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n552_), .A2(new_n587_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT94), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n552_), .A2(KEYINPUT94), .A3(new_n587_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n573_), .B1(new_n589_), .B2(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n514_), .B1(new_n518_), .B2(new_n516_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n524_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n501_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(new_n527_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n525_), .A2(KEYINPUT90), .A3(new_n501_), .ZN(new_n600_));
  AOI22_X1  g399(.A1(new_n599_), .A2(new_n600_), .B1(new_n516_), .B2(new_n515_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n595_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n569_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n565_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n567_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n295_), .A2(new_n296_), .ZN(new_n606_));
  OAI21_X1  g405(.A(KEYINPUT75), .B1(new_n239_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT75), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n297_), .A2(new_n608_), .A3(new_n223_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n239_), .A2(new_n304_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n607_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G229gat), .A2(G233gat), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n223_), .B(new_n304_), .Z(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n613_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT74), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT74), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n615_), .A2(new_n618_), .A3(new_n613_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n614_), .A2(new_n617_), .A3(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G113gat), .B(G141gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G169gat), .B(G197gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n620_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n623_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n614_), .A2(new_n617_), .A3(new_n619_), .A4(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT76), .ZN(new_n628_));
  OAI21_X1  g427(.A(KEYINPUT99), .B1(new_n605_), .B2(new_n628_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n601_), .A2(new_n568_), .A3(new_n554_), .A4(new_n565_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n599_), .A2(new_n600_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n553_), .B1(new_n631_), .B2(new_n517_), .ZN(new_n632_));
  AOI22_X1  g431(.A1(new_n632_), .A2(new_n568_), .B1(new_n595_), .B2(new_n601_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n630_), .B1(new_n633_), .B2(new_n565_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n635_));
  INV_X1    g434(.A(new_n628_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n634_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n349_), .B1(new_n629_), .B2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n638_), .A2(new_n214_), .A3(new_n553_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n640_), .A2(KEYINPUT38), .ZN(new_n641_));
  INV_X1    g440(.A(new_n325_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n605_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n256_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n347_), .A2(new_n627_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n643_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(KEYINPUT100), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT100), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n643_), .A2(new_n649_), .A3(new_n646_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(G1gat), .B1(new_n651_), .B2(new_n554_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n640_), .A2(KEYINPUT38), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n641_), .A2(new_n652_), .A3(new_n653_), .ZN(G1324gat));
  XNOR2_X1  g453(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(KEYINPUT102), .B1(new_n647_), .B2(new_n568_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT102), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n643_), .A2(new_n658_), .A3(new_n463_), .A4(new_n646_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n657_), .A2(G8gat), .A3(new_n659_), .ZN(new_n660_));
  XOR2_X1   g459(.A(KEYINPUT103), .B(KEYINPUT39), .Z(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n657_), .A2(G8gat), .A3(new_n659_), .A4(new_n661_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n568_), .A2(G8gat), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n638_), .A2(KEYINPUT101), .A3(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(KEYINPUT101), .B1(new_n638_), .B2(new_n666_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n656_), .B1(new_n665_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n669_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n671_), .A2(new_n664_), .A3(new_n663_), .A4(new_n655_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(G1325gat));
  INV_X1    g472(.A(G15gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n638_), .A2(new_n674_), .A3(new_n565_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n648_), .A2(new_n565_), .A3(new_n650_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n676_), .A2(G15gat), .A3(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n677_), .B1(new_n676_), .B2(G15gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n675_), .B1(new_n678_), .B2(new_n679_), .ZN(G1326gat));
  NAND3_X1  g479(.A1(new_n648_), .A2(new_n529_), .A3(new_n650_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(G22gat), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT106), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT106), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n681_), .A2(new_n684_), .A3(G22gat), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT42), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n683_), .A2(KEYINPUT42), .A3(new_n685_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n638_), .A2(new_n212_), .A3(new_n529_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n688_), .A2(new_n689_), .A3(new_n690_), .ZN(G1327gat));
  INV_X1    g490(.A(new_n645_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n327_), .A2(new_n348_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n634_), .B2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n565_), .B1(new_n569_), .B2(new_n602_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n693_), .B(new_n694_), .C1(new_n696_), .C2(new_n567_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n644_), .B(new_n692_), .C1(new_n695_), .C2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n700_), .A2(KEYINPUT107), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(KEYINPUT107), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n699_), .A2(new_n701_), .A3(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n694_), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT43), .B1(new_n605_), .B2(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n256_), .B1(new_n705_), .B2(new_n697_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n706_), .A2(KEYINPUT107), .A3(new_n700_), .A4(new_n692_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n703_), .A2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n553_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT108), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n708_), .A2(new_n711_), .A3(new_n553_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n710_), .A2(G29gat), .A3(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n629_), .A2(new_n637_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n256_), .A2(new_n325_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n347_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n714_), .A2(new_n718_), .ZN(new_n719_));
  OR3_X1    g518(.A1(new_n719_), .A2(G29gat), .A3(new_n554_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n713_), .A2(new_n720_), .ZN(G1328gat));
  INV_X1    g520(.A(G36gat), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n714_), .A2(new_n722_), .A3(new_n463_), .A4(new_n718_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT45), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n568_), .B1(new_n703_), .B2(new_n707_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n725_), .B2(new_n722_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT46), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n724_), .B(KEYINPUT46), .C1(new_n725_), .C2(new_n722_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1329gat));
  NAND3_X1  g529(.A1(new_n708_), .A2(G43gat), .A3(new_n565_), .ZN(new_n731_));
  INV_X1    g530(.A(G43gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n732_), .B1(new_n719_), .B2(new_n604_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n731_), .A2(new_n733_), .A3(new_n735_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1330gat));
  NOR2_X1   g538(.A1(new_n719_), .A2(new_n601_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n708_), .A2(new_n529_), .ZN(new_n741_));
  MUX2_X1   g540(.A(new_n740_), .B(new_n741_), .S(G50gat), .Z(G1331gat));
  NAND4_X1  g541(.A1(new_n643_), .A2(new_n256_), .A3(new_n717_), .A4(new_n628_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n744_), .A2(G57gat), .A3(new_n553_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT111), .Z(new_n746_));
  INV_X1    g545(.A(new_n627_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n704_), .A2(new_n256_), .A3(new_n717_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(KEYINPUT110), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n749_), .A2(new_n605_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(KEYINPUT110), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(G57gat), .B1(new_n753_), .B2(new_n553_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n746_), .A2(new_n754_), .ZN(G1332gat));
  OAI21_X1  g554(.A(G64gat), .B1(new_n743_), .B2(new_n568_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT48), .Z(new_n757_));
  NOR3_X1   g556(.A1(new_n752_), .A2(G64gat), .A3(new_n568_), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1333gat));
  OAI21_X1  g558(.A(G71gat), .B1(new_n743_), .B2(new_n604_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT49), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n752_), .A2(G71gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n761_), .B1(new_n604_), .B2(new_n762_), .ZN(G1334gat));
  NOR2_X1   g562(.A1(new_n743_), .A2(new_n601_), .ZN(new_n764_));
  INV_X1    g563(.A(G78gat), .ZN(new_n765_));
  OR3_X1    g564(.A1(new_n764_), .A2(KEYINPUT112), .A3(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(KEYINPUT112), .B1(new_n764_), .B2(new_n765_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT50), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n753_), .A2(new_n765_), .A3(new_n529_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n766_), .A2(KEYINPUT50), .A3(new_n767_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n770_), .A2(new_n771_), .A3(new_n772_), .ZN(G1335gat));
  NOR2_X1   g572(.A1(new_n347_), .A2(new_n627_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n634_), .A2(new_n715_), .A3(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(G85gat), .B1(new_n776_), .B2(new_n553_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n706_), .A2(new_n774_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n778_), .A2(new_n553_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n777_), .B1(new_n779_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g579(.A(G92gat), .B1(new_n776_), .B2(new_n463_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n463_), .A2(G92gat), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n778_), .B2(new_n782_), .ZN(G1337gat));
  AND3_X1   g582(.A1(new_n776_), .A2(new_n565_), .A3(new_n259_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n778_), .A2(new_n565_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n785_), .B2(G99gat), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT51), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n786_), .B(new_n788_), .ZN(G1338gat));
  NAND3_X1  g588(.A1(new_n776_), .A2(new_n260_), .A3(new_n529_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n706_), .A2(new_n529_), .A3(new_n774_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n791_), .A2(new_n792_), .A3(G106gat), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n791_), .B2(G106gat), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n790_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT53), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n797_), .B(new_n790_), .C1(new_n793_), .C2(new_n794_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(G1339gat));
  NAND2_X1  g598(.A1(new_n288_), .A2(new_n328_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n330_), .A2(new_n331_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n333_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n334_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n332_), .A2(KEYINPUT55), .A3(new_n333_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n342_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT56), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(KEYINPUT114), .A3(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n344_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n810_), .B1(new_n811_), .B2(KEYINPUT56), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(KEYINPUT56), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n809_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n334_), .A2(new_n336_), .A3(new_n344_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n747_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n344_), .B1(new_n334_), .B2(new_n336_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n815_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n611_), .A2(KEYINPUT115), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n607_), .A2(new_n609_), .A3(new_n822_), .A4(new_n610_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n821_), .A2(new_n613_), .A3(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n615_), .A2(new_n612_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n824_), .A2(new_n623_), .A3(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n626_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n818_), .B1(new_n820_), .B2(new_n827_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n826_), .A2(new_n626_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n829_), .A2(new_n346_), .A3(KEYINPUT116), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n817_), .A2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n833_), .A2(KEYINPUT57), .A3(new_n325_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n831_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(new_n642_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n807_), .A2(new_n808_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n813_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(new_n345_), .A3(new_n829_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT58), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n839_), .A2(KEYINPUT58), .A3(new_n345_), .A4(new_n829_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n694_), .A3(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n834_), .A2(new_n837_), .A3(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n644_), .ZN(new_n846_));
  OR3_X1    g645(.A1(new_n349_), .A2(KEYINPUT54), .A3(new_n636_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT54), .B1(new_n349_), .B2(new_n636_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n846_), .A2(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n463_), .A2(new_n529_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n851_), .A2(new_n553_), .A3(new_n565_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n850_), .A2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(G113gat), .B1(new_n855_), .B2(new_n627_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n846_), .A2(KEYINPUT117), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n845_), .A2(new_n858_), .A3(new_n644_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n849_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n852_), .A2(KEYINPUT59), .ZN(new_n862_));
  AOI22_X1  g661(.A1(new_n861_), .A2(new_n862_), .B1(KEYINPUT59), .B2(new_n854_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n636_), .A2(G113gat), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n856_), .B1(new_n863_), .B2(new_n864_), .ZN(G1340gat));
  INV_X1    g664(.A(G120gat), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n866_), .B1(new_n347_), .B2(KEYINPUT60), .ZN(new_n867_));
  OAI21_X1  g666(.A(KEYINPUT118), .B1(new_n866_), .B2(KEYINPUT60), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n854_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n870_), .B2(new_n867_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n863_), .A2(new_n717_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n871_), .B1(new_n873_), .B2(new_n866_), .ZN(G1341gat));
  INV_X1    g673(.A(G127gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n875_), .B1(new_n854_), .B2(new_n644_), .ZN(new_n876_));
  AOI22_X1  g675(.A1(new_n845_), .A2(new_n644_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n877_));
  OAI21_X1  g676(.A(KEYINPUT59), .B1(new_n877_), .B2(new_n852_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n849_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n879_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n862_), .ZN(new_n881_));
  OAI211_X1 g680(.A(G127gat), .B(new_n878_), .C1(new_n880_), .C2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n876_), .B1(new_n882_), .B2(new_n644_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  OAI211_X1 g684(.A(KEYINPUT119), .B(new_n876_), .C1(new_n882_), .C2(new_n644_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1342gat));
  INV_X1    g686(.A(KEYINPUT120), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n694_), .B(new_n878_), .C1(new_n880_), .C2(new_n881_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(G134gat), .ZN(new_n890_));
  NOR4_X1   g689(.A1(new_n877_), .A2(G134gat), .A3(new_n325_), .A4(new_n852_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n888_), .B1(new_n890_), .B2(new_n892_), .ZN(new_n893_));
  AOI211_X1 g692(.A(KEYINPUT120), .B(new_n891_), .C1(new_n889_), .C2(G134gat), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1343gat));
  NOR3_X1   g694(.A1(new_n463_), .A2(new_n601_), .A3(new_n554_), .ZN(new_n896_));
  AND3_X1   g695(.A1(new_n850_), .A2(new_n604_), .A3(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n627_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n717_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g700(.A1(new_n897_), .A2(new_n256_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(KEYINPUT121), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT121), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n897_), .A2(new_n904_), .A3(new_n256_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n905_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT61), .B(G155gat), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n908_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n903_), .A2(new_n905_), .A3(new_n907_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1346gat));
  AND3_X1   g710(.A1(new_n897_), .A2(G162gat), .A3(new_n694_), .ZN(new_n912_));
  AOI21_X1  g711(.A(G162gat), .B1(new_n897_), .B2(new_n642_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1347gat));
  NOR3_X1   g713(.A1(new_n529_), .A2(new_n568_), .A3(new_n566_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n861_), .A2(new_n915_), .ZN(new_n916_));
  OAI21_X1  g715(.A(G169gat), .B1(new_n916_), .B2(new_n747_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n915_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n880_), .A2(new_n920_), .ZN(new_n921_));
  OAI211_X1 g720(.A(new_n921_), .B(new_n627_), .C1(new_n365_), .C2(new_n364_), .ZN(new_n922_));
  OAI211_X1 g721(.A(KEYINPUT62), .B(G169gat), .C1(new_n916_), .C2(new_n747_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n919_), .A2(new_n922_), .A3(new_n923_), .ZN(G1348gat));
  NAND2_X1  g723(.A1(new_n850_), .A2(new_n915_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n925_), .A2(new_n381_), .A3(new_n347_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n921_), .A2(new_n717_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n355_), .A2(new_n356_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n926_), .B1(new_n927_), .B2(new_n928_), .ZN(G1349gat));
  INV_X1    g728(.A(G183gat), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n930_), .B1(new_n925_), .B2(new_n644_), .ZN(new_n931_));
  OR2_X1    g730(.A1(new_n644_), .A2(new_n374_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n916_), .B2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(KEYINPUT122), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n935_));
  OAI211_X1 g734(.A(new_n935_), .B(new_n931_), .C1(new_n916_), .C2(new_n932_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n934_), .A2(new_n936_), .ZN(G1350gat));
  OAI21_X1  g736(.A(G190gat), .B1(new_n916_), .B2(new_n704_), .ZN(new_n938_));
  AND2_X1   g737(.A1(new_n642_), .A2(new_n417_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n921_), .A2(new_n939_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n938_), .A2(KEYINPUT123), .A3(new_n940_), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT123), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n376_), .B1(new_n921_), .B2(new_n694_), .ZN(new_n943_));
  AND3_X1   g742(.A1(new_n861_), .A2(new_n915_), .A3(new_n939_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n942_), .B1(new_n943_), .B2(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n941_), .A2(new_n945_), .ZN(G1351gat));
  NOR2_X1   g745(.A1(new_n877_), .A2(new_n565_), .ZN(new_n947_));
  NOR3_X1   g746(.A1(new_n601_), .A2(new_n568_), .A3(new_n553_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(new_n948_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n949_), .A2(new_n747_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(new_n409_), .ZN(G1352gat));
  INV_X1    g750(.A(new_n949_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n952_), .A2(new_n717_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n953_), .A2(G204gat), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n954_), .B1(new_n953_), .B2(new_n404_), .ZN(G1353gat));
  AOI21_X1  g754(.A(new_n644_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n956_), .B(KEYINPUT124), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n949_), .A2(new_n957_), .ZN(new_n958_));
  INV_X1    g757(.A(KEYINPUT126), .ZN(new_n959_));
  NOR2_X1   g758(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n960_), .B(KEYINPUT125), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n958_), .A2(new_n959_), .A3(new_n961_), .ZN(new_n962_));
  XNOR2_X1  g761(.A(new_n961_), .B(new_n959_), .ZN(new_n963_));
  OAI21_X1  g762(.A(new_n962_), .B1(new_n963_), .B2(new_n958_), .ZN(G1354gat));
  AOI21_X1  g763(.A(G218gat), .B1(new_n952_), .B2(new_n642_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n949_), .A2(new_n704_), .ZN(new_n966_));
  AOI21_X1  g765(.A(new_n965_), .B1(G218gat), .B2(new_n966_), .ZN(G1355gat));
endmodule


