//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n845_, new_n846_,
    new_n847_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G113gat), .B(G120gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(KEYINPUT82), .Z(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT31), .ZN(new_n206_));
  INV_X1    g005(.A(G169gat), .ZN(new_n207_));
  INV_X1    g006(.A(G176gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n207_), .A2(new_n208_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n210_), .A2(KEYINPUT24), .A3(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT78), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT23), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n211_), .A2(KEYINPUT24), .ZN(new_n218_));
  NOR3_X1   g017(.A1(new_n214_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n212_), .A2(new_n213_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT25), .B(G183gat), .ZN(new_n221_));
  INV_X1    g020(.A(G190gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT26), .B1(new_n222_), .B2(KEYINPUT77), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n222_), .A2(KEYINPUT26), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n221_), .B(new_n223_), .C1(new_n224_), .C2(KEYINPUT77), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n220_), .A2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n216_), .B1(G183gat), .B2(G190gat), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n227_), .A2(new_n210_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT22), .B1(new_n207_), .B2(KEYINPUT79), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n207_), .A2(KEYINPUT22), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n208_), .B(new_n229_), .C1(new_n230_), .C2(KEYINPUT79), .ZN(new_n231_));
  AOI22_X1  g030(.A1(new_n219_), .A2(new_n226_), .B1(new_n228_), .B2(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(G71gat), .B(G99gat), .Z(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT81), .ZN(new_n234_));
  XOR2_X1   g033(.A(G15gat), .B(G43gat), .Z(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n232_), .B(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G227gat), .A2(G233gat), .ZN(new_n238_));
  XOR2_X1   g037(.A(new_n238_), .B(KEYINPUT80), .Z(new_n239_));
  XOR2_X1   g038(.A(new_n239_), .B(KEYINPUT30), .Z(new_n240_));
  XNOR2_X1  g039(.A(new_n237_), .B(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n206_), .B1(new_n241_), .B2(KEYINPUT83), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n242_), .B1(KEYINPUT83), .B2(new_n241_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(KEYINPUT83), .A3(new_n206_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G141gat), .A2(G148gat), .ZN(new_n246_));
  OR2_X1    g045(.A1(G141gat), .A2(G148gat), .ZN(new_n247_));
  OR2_X1    g046(.A1(G155gat), .A2(G162gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G155gat), .A2(G162gat), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n248_), .B1(KEYINPUT1), .B2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT84), .B1(new_n249_), .B2(KEYINPUT1), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n249_), .A2(KEYINPUT84), .A3(KEYINPUT1), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n246_), .B(new_n247_), .C1(new_n252_), .C2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n247_), .B(KEYINPUT3), .ZN(new_n255_));
  XOR2_X1   g054(.A(new_n246_), .B(KEYINPUT2), .Z(new_n256_));
  OAI211_X1 g055(.A(new_n248_), .B(new_n249_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n254_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT29), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT28), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT85), .B(G197gat), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT86), .ZN(new_n264_));
  INV_X1    g063(.A(G204gat), .ZN(new_n265_));
  NOR3_X1   g064(.A1(new_n263_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n263_), .A2(new_n265_), .ZN(new_n268_));
  INV_X1    g067(.A(G197gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n264_), .B1(new_n269_), .B2(G204gat), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n267_), .B(KEYINPUT87), .C1(new_n268_), .C2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT87), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n268_), .A2(new_n270_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n272_), .B1(new_n273_), .B2(new_n266_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G211gat), .B(G218gat), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT21), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n271_), .A2(new_n274_), .A3(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n276_), .B1(new_n273_), .B2(new_n266_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n276_), .B1(G197gat), .B2(G204gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n280_), .B1(new_n263_), .B2(G204gat), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(new_n281_), .A3(new_n275_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n278_), .A2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n283_), .B1(new_n260_), .B2(new_n259_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n262_), .B(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G228gat), .A2(G233gat), .ZN(new_n286_));
  INV_X1    g085(.A(G78gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(G106gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G22gat), .B(G50gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n285_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n283_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(new_n232_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT20), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT26), .B(G190gat), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n217_), .B1(new_n221_), .B2(new_n297_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n298_), .B(new_n212_), .C1(KEYINPUT24), .C2(new_n211_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT22), .B(G169gat), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n209_), .B1(new_n300_), .B2(new_n208_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n227_), .A2(new_n301_), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n302_), .A2(KEYINPUT88), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(KEYINPUT88), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n299_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n296_), .B1(new_n305_), .B2(new_n283_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n295_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G226gat), .A2(G233gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT19), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n219_), .A2(new_n226_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n228_), .A2(new_n231_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n296_), .B1(new_n283_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n309_), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n314_), .B(new_n315_), .C1(new_n283_), .C2(new_n305_), .ZN(new_n316_));
  XOR2_X1   g115(.A(G8gat), .B(G36gat), .Z(new_n317_));
  XNOR2_X1  g116(.A(G64gat), .B(G92gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n319_), .B(new_n320_), .Z(new_n321_));
  NAND3_X1  g120(.A1(new_n310_), .A2(new_n316_), .A3(new_n321_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n278_), .A2(new_n282_), .A3(new_n299_), .A4(new_n302_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n315_), .B1(new_n314_), .B2(new_n323_), .ZN(new_n324_));
  OR2_X1    g123(.A1(new_n324_), .A2(KEYINPUT93), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(KEYINPUT93), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT94), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n327_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n295_), .A2(new_n306_), .A3(KEYINPUT94), .A4(new_n315_), .ZN(new_n329_));
  AOI22_X1  g128(.A1(new_n325_), .A2(new_n326_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  OAI211_X1 g129(.A(KEYINPUT27), .B(new_n322_), .C1(new_n330_), .C2(new_n321_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n204_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n258_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n254_), .A2(new_n204_), .A3(new_n257_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n333_), .A2(KEYINPUT4), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT4), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n258_), .A2(new_n336_), .A3(new_n332_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G225gat), .A2(G233gat), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G1gat), .B(G29gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(G85gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT0), .B(G57gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n333_), .A2(new_n334_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(new_n339_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n341_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n345_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n347_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n339_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n349_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n348_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n321_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n314_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n315_), .B1(new_n305_), .B2(new_n283_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n315_), .B1(new_n295_), .B2(new_n306_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n355_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT90), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n322_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT27), .ZN(new_n363_));
  OAI211_X1 g162(.A(KEYINPUT90), .B(new_n355_), .C1(new_n358_), .C2(new_n359_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n362_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  AND4_X1   g164(.A1(new_n293_), .A2(new_n331_), .A3(new_n354_), .A4(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n362_), .A2(new_n364_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n345_), .B1(new_n341_), .B2(new_n347_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT33), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT33), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n346_), .A2(new_n339_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n371_), .A2(new_n349_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n335_), .A2(new_n339_), .A3(new_n337_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n370_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n369_), .B1(new_n374_), .B2(new_n368_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n367_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n321_), .A2(KEYINPUT32), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT91), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n310_), .A2(new_n316_), .A3(new_n380_), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n381_), .A2(KEYINPUT92), .B1(new_n352_), .B2(new_n348_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT92), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n310_), .A2(new_n383_), .A3(new_n380_), .A4(new_n316_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n382_), .B(new_n384_), .C1(new_n330_), .C2(new_n378_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n293_), .B1(new_n377_), .B2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n245_), .B1(new_n366_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT95), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n331_), .A2(new_n365_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n389_), .A2(new_n293_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n245_), .A2(new_n353_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT95), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n393_), .B(new_n245_), .C1(new_n366_), .C2(new_n386_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n388_), .A2(new_n392_), .A3(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT76), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G15gat), .B(G22gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT73), .B(G8gat), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(G1gat), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT14), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n397_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G1gat), .B(G8gat), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n397_), .B(new_n404_), .C1(new_n401_), .C2(new_n402_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G29gat), .B(G36gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G43gat), .B(G50gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n408_), .A2(new_n411_), .ZN(new_n412_));
  XOR2_X1   g211(.A(new_n409_), .B(new_n410_), .Z(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT15), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT15), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n411_), .A2(new_n415_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n406_), .A2(new_n414_), .A3(new_n407_), .A4(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G229gat), .A2(G233gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT75), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n412_), .A2(new_n417_), .A3(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n406_), .A2(new_n407_), .A3(new_n413_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n418_), .B1(new_n412_), .B2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n396_), .B1(new_n420_), .B2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G113gat), .B(G141gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G169gat), .B(G197gat), .ZN(new_n425_));
  XOR2_X1   g224(.A(new_n424_), .B(new_n425_), .Z(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n423_), .A2(new_n427_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n396_), .B(new_n426_), .C1(new_n420_), .C2(new_n422_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(G230gat), .ZN(new_n432_));
  INV_X1    g231(.A(G233gat), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  AND2_X1   g233(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n435_));
  NOR2_X1   g234(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n436_));
  NOR3_X1   g235(.A1(new_n435_), .A2(new_n436_), .A3(KEYINPUT64), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT64), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT10), .ZN(new_n439_));
  INV_X1    g238(.A(G99gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n438_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n289_), .B1(new_n437_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G99gat), .A2(G106gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT6), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT6), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(G99gat), .A3(G106gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(G85gat), .ZN(new_n450_));
  INV_X1    g249(.A(G92gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G85gat), .A2(G92gat), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n452_), .A2(KEYINPUT9), .A3(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT9), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n455_), .A2(G85gat), .A3(G92gat), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n449_), .A2(new_n454_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n444_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n452_), .A2(KEYINPUT65), .A3(new_n453_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NOR3_X1   g260(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  AOI211_X1 g262(.A(KEYINPUT8), .B(new_n459_), .C1(new_n463_), .C2(new_n449_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT8), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT7), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(new_n440_), .A3(new_n289_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n447_), .B1(G99gat), .B2(G106gat), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n445_), .A2(KEYINPUT6), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n460_), .B(new_n467_), .C1(new_n468_), .C2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n459_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n465_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n458_), .B1(new_n464_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT66), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  XOR2_X1   g274(.A(G71gat), .B(G78gat), .Z(new_n476_));
  XNOR2_X1  g275(.A(G57gat), .B(G64gat), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n476_), .B1(KEYINPUT11), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT67), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n479_), .B1(new_n477_), .B2(KEYINPUT11), .ZN(new_n480_));
  INV_X1    g279(.A(G64gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(G57gat), .ZN(new_n482_));
  INV_X1    g281(.A(G57gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(G64gat), .ZN(new_n484_));
  AND4_X1   g283(.A1(new_n479_), .A2(new_n482_), .A3(new_n484_), .A4(KEYINPUT11), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n478_), .B1(new_n480_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n482_), .A2(new_n484_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT11), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT67), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n477_), .A2(new_n479_), .A3(KEYINPUT11), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n487_), .A2(new_n488_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .A4(new_n476_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n486_), .A2(new_n492_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n458_), .B(KEYINPUT66), .C1(new_n464_), .C2(new_n472_), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n475_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n493_), .B1(new_n475_), .B2(new_n494_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n434_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G120gat), .B(G148gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT5), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G176gat), .B(G204gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT68), .ZN(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT64), .B1(new_n435_), .B2(new_n436_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n441_), .A2(new_n438_), .A3(new_n442_), .ZN(new_n504_));
  AOI21_X1  g303(.A(G106gat), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n449_), .A2(new_n454_), .A3(new_n456_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n468_), .A2(new_n469_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n467_), .A2(new_n460_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n471_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT8), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n470_), .A2(new_n465_), .A3(new_n471_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n507_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n486_), .A2(new_n492_), .A3(KEYINPUT12), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n502_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n486_), .A2(new_n492_), .A3(KEYINPUT12), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n516_), .A2(new_n473_), .A3(KEYINPUT68), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n518_), .B1(new_n496_), .B2(KEYINPUT12), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n475_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n434_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n497_), .B(new_n501_), .C1(new_n519_), .C2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT70), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n520_), .A2(new_n521_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n493_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n511_), .A2(new_n512_), .ZN(new_n527_));
  AOI21_X1  g326(.A(KEYINPUT66), .B1(new_n527_), .B2(new_n458_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n494_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n526_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT12), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n525_), .A2(new_n532_), .A3(new_n518_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT70), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n533_), .A2(new_n534_), .A3(new_n497_), .A4(new_n501_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n524_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT71), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n533_), .A2(new_n497_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n501_), .B(KEYINPUT69), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n536_), .A2(new_n537_), .A3(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n537_), .B1(new_n536_), .B2(new_n540_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT13), .ZN(new_n543_));
  OR3_X1    g342(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n543_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n475_), .A2(new_n411_), .A3(new_n494_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n473_), .A2(new_n414_), .A3(new_n416_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G232gat), .A2(G233gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT34), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n548_), .B(new_n549_), .C1(KEYINPUT35), .C2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(KEYINPUT35), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G190gat), .B(G218gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT72), .ZN(new_n556_));
  XOR2_X1   g355(.A(G134gat), .B(G162gat), .Z(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT36), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n554_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n554_), .A2(new_n559_), .A3(new_n558_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n563_), .A2(KEYINPUT37), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT37), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n565_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G231gat), .A2(G233gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n493_), .B(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n569_), .B(new_n408_), .Z(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(G127gat), .B(G155gat), .Z(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT16), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G183gat), .B(G211gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT74), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT17), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n571_), .A2(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n578_), .B1(new_n577_), .B2(new_n575_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n570_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n567_), .A2(new_n582_), .ZN(new_n583_));
  AND4_X1   g382(.A1(new_n395_), .A2(new_n431_), .A3(new_n547_), .A4(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n584_), .B(KEYINPUT96), .Z(new_n585_));
  NAND3_X1  g384(.A1(new_n585_), .A2(new_n400_), .A3(new_n353_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT97), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT38), .ZN(new_n588_));
  OR3_X1    g387(.A1(new_n586_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n563_), .B(KEYINPUT98), .Z(new_n590_));
  AND2_X1   g389(.A1(new_n395_), .A2(new_n590_), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n546_), .A2(new_n430_), .A3(new_n582_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n400_), .B1(new_n593_), .B2(new_n353_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n586_), .B1(new_n588_), .B2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n587_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n589_), .A2(new_n595_), .A3(new_n596_), .ZN(G1324gat));
  NAND2_X1  g396(.A1(new_n593_), .A2(new_n389_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(G8gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT39), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n585_), .A2(new_n389_), .A3(new_n399_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT40), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n600_), .A2(KEYINPUT40), .A3(new_n601_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(G1325gat));
  INV_X1    g405(.A(new_n245_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n593_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(G15gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(KEYINPUT99), .B(KEYINPUT41), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n610_), .ZN(new_n612_));
  INV_X1    g411(.A(G15gat), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n585_), .A2(new_n613_), .A3(new_n607_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n611_), .A2(new_n612_), .A3(new_n614_), .ZN(G1326gat));
  INV_X1    g414(.A(G22gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n293_), .B(KEYINPUT100), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n616_), .B1(new_n593_), .B2(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n619_), .B(KEYINPUT42), .Z(new_n620_));
  NAND3_X1  g419(.A1(new_n585_), .A2(new_n616_), .A3(new_n618_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(G1327gat));
  AND2_X1   g421(.A1(new_n395_), .A2(new_n431_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n590_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(new_n582_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n625_), .A2(new_n546_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n623_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(G29gat), .B1(new_n628_), .B2(new_n353_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT103), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n394_), .A2(new_n392_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n331_), .A2(new_n293_), .A3(new_n354_), .A4(new_n365_), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n330_), .A2(new_n378_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n381_), .A2(KEYINPUT92), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n634_), .A2(new_n384_), .A3(new_n353_), .ZN(new_n635_));
  AOI22_X1  g434(.A1(new_n633_), .A2(new_n635_), .B1(new_n367_), .B2(new_n376_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n632_), .B1(new_n636_), .B2(new_n293_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n393_), .B1(new_n637_), .B2(new_n245_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n567_), .B1(new_n631_), .B2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT43), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT43), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n641_), .B(new_n567_), .C1(new_n631_), .C2(new_n638_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n547_), .A2(new_n431_), .A3(new_n582_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(KEYINPUT101), .ZN(new_n644_));
  INV_X1    g443(.A(new_n582_), .ZN(new_n645_));
  OR4_X1    g444(.A1(KEYINPUT101), .A2(new_n546_), .A3(new_n430_), .A4(new_n645_), .ZN(new_n646_));
  AOI22_X1  g445(.A1(new_n640_), .A2(new_n642_), .B1(new_n644_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n630_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT102), .B1(KEYINPUT103), .B2(KEYINPUT44), .ZN(new_n650_));
  OAI22_X1  g449(.A1(new_n649_), .A2(KEYINPUT44), .B1(new_n647_), .B2(new_n650_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n353_), .A2(G29gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n629_), .B1(new_n651_), .B2(new_n652_), .ZN(G1328gat));
  INV_X1    g452(.A(KEYINPUT46), .ZN(new_n654_));
  INV_X1    g453(.A(G36gat), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n623_), .A2(new_n655_), .A3(new_n389_), .A4(new_n626_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT45), .Z(new_n657_));
  NAND2_X1  g456(.A1(new_n646_), .A2(new_n644_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n642_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n641_), .B1(new_n395_), .B2(new_n567_), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n648_), .B(new_n658_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT44), .B1(new_n661_), .B2(KEYINPUT103), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n647_), .A2(new_n650_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n389_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n657_), .B1(new_n664_), .B2(G36gat), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT104), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n654_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n655_), .B1(new_n651_), .B2(new_n389_), .ZN(new_n668_));
  OAI211_X1 g467(.A(KEYINPUT104), .B(KEYINPUT46), .C1(new_n668_), .C2(new_n657_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n667_), .A2(new_n669_), .ZN(G1329gat));
  INV_X1    g469(.A(G43gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n671_), .B1(new_n651_), .B2(new_n607_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT47), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n627_), .A2(G43gat), .A3(new_n245_), .ZN(new_n674_));
  OR3_X1    g473(.A1(new_n672_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n673_), .B1(new_n672_), .B2(new_n674_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1330gat));
  AOI21_X1  g476(.A(G50gat), .B1(new_n628_), .B2(new_n618_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n293_), .A2(G50gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n678_), .B1(new_n651_), .B2(new_n679_), .ZN(G1331gat));
  NOR3_X1   g479(.A1(new_n547_), .A2(new_n431_), .A3(new_n582_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n591_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(G57gat), .B1(new_n683_), .B2(new_n354_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n395_), .A2(new_n430_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n546_), .A2(new_n583_), .A3(KEYINPUT105), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n687_));
  INV_X1    g486(.A(new_n583_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n687_), .B1(new_n547_), .B2(new_n688_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n685_), .A2(new_n686_), .A3(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n690_), .A2(new_n483_), .A3(new_n353_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n684_), .A2(new_n691_), .ZN(G1332gat));
  AOI21_X1  g491(.A(new_n481_), .B1(new_n682_), .B2(new_n389_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT48), .Z(new_n694_));
  NAND3_X1  g493(.A1(new_n690_), .A2(new_n481_), .A3(new_n389_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1333gat));
  INV_X1    g495(.A(G71gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n697_), .B1(new_n682_), .B2(new_n607_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT49), .Z(new_n699_));
  NAND3_X1  g498(.A1(new_n690_), .A2(new_n697_), .A3(new_n607_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1334gat));
  AOI21_X1  g500(.A(new_n287_), .B1(new_n682_), .B2(new_n618_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT50), .Z(new_n703_));
  NAND3_X1  g502(.A1(new_n690_), .A2(new_n287_), .A3(new_n618_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1335gat));
  NOR2_X1   g504(.A1(new_n625_), .A2(new_n547_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n685_), .A2(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n450_), .B1(new_n707_), .B2(new_n354_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT106), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n640_), .A2(new_n642_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n547_), .A2(new_n431_), .A3(new_n645_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n712_), .A2(KEYINPUT107), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(KEYINPUT107), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n354_), .A2(new_n450_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n709_), .B1(new_n715_), .B2(new_n716_), .ZN(G1336gat));
  INV_X1    g516(.A(new_n707_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n718_), .A2(new_n451_), .A3(new_n389_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n389_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n720_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n719_), .B1(new_n721_), .B2(new_n451_), .ZN(G1337gat));
  OAI211_X1 g521(.A(new_n718_), .B(new_n607_), .C1(new_n437_), .C2(new_n443_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT108), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n245_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n725_), .B2(new_n440_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT51), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT51), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n724_), .B(new_n728_), .C1(new_n440_), .C2(new_n725_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1338gat));
  NAND3_X1  g529(.A1(new_n710_), .A2(new_n293_), .A3(new_n711_), .ZN(new_n731_));
  AOI21_X1  g530(.A(KEYINPUT110), .B1(new_n731_), .B2(G106gat), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT52), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n731_), .A2(KEYINPUT110), .A3(G106gat), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n732_), .A2(new_n733_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n293_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n707_), .A2(G106gat), .A3(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT109), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n736_), .A2(new_n737_), .A3(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT53), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT53), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n736_), .A2(new_n743_), .A3(new_n737_), .A4(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1339gat));
  NAND3_X1  g544(.A1(new_n390_), .A2(new_n607_), .A3(new_n353_), .ZN(new_n746_));
  XOR2_X1   g545(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n747_));
  NAND3_X1  g546(.A1(new_n547_), .A2(new_n430_), .A3(new_n583_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT54), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT55), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n750_), .B1(new_n519_), .B2(new_n522_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n525_), .A2(new_n532_), .A3(KEYINPUT55), .A4(new_n518_), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n518_), .B(new_n520_), .C1(new_n496_), .C2(KEYINPUT12), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(new_n434_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n751_), .A2(new_n752_), .A3(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n755_), .A2(KEYINPUT56), .A3(new_n539_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT112), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n539_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT56), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT112), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n755_), .A2(new_n761_), .A3(KEYINPUT56), .A4(new_n539_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n757_), .A2(new_n760_), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n412_), .A2(new_n421_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n419_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n419_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n412_), .A2(new_n417_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n427_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n420_), .A2(new_n422_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(new_n770_), .B2(new_n427_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n536_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n763_), .B(new_n772_), .C1(new_n773_), .C2(KEYINPUT58), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n567_), .ZN(new_n775_));
  AOI211_X1 g574(.A(new_n773_), .B(KEYINPUT58), .C1(new_n763_), .C2(new_n772_), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n771_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n430_), .B1(new_n524_), .B2(new_n535_), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n755_), .A2(KEYINPUT56), .A3(new_n539_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT56), .B1(new_n755_), .B2(new_n539_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n779_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT111), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n779_), .B(new_n784_), .C1(new_n780_), .C2(new_n781_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n778_), .A2(new_n783_), .A3(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT57), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(new_n590_), .A3(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n787_), .B1(new_n786_), .B2(new_n590_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n777_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n582_), .ZN(new_n792_));
  AOI211_X1 g591(.A(new_n746_), .B(new_n747_), .C1(new_n749_), .C2(new_n792_), .ZN(new_n793_));
  XOR2_X1   g592(.A(new_n793_), .B(KEYINPUT119), .Z(new_n794_));
  NOR2_X1   g593(.A1(new_n775_), .A2(new_n776_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n786_), .A2(new_n590_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT57), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n795_), .B1(new_n797_), .B2(new_n788_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n582_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n777_), .B(new_n799_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n749_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  OAI211_X1 g604(.A(KEYINPUT115), .B(new_n749_), .C1(new_n800_), .C2(new_n802_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n746_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n805_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n808_), .A2(new_n809_), .A3(KEYINPUT59), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(new_n808_), .B2(KEYINPUT59), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n431_), .B(new_n794_), .C1(new_n810_), .C2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(G113gat), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n808_), .B(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(G113gat), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n816_), .A3(new_n431_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n813_), .A2(new_n817_), .ZN(G1340gat));
  OAI211_X1 g617(.A(new_n546_), .B(new_n794_), .C1(new_n810_), .C2(new_n811_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(G120gat), .ZN(new_n820_));
  INV_X1    g619(.A(G120gat), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n821_), .B1(new_n547_), .B2(KEYINPUT60), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n815_), .B(new_n822_), .C1(KEYINPUT60), .C2(new_n821_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n820_), .A2(new_n823_), .ZN(G1341gat));
  XNOR2_X1  g623(.A(new_n793_), .B(KEYINPUT119), .ZN(new_n825_));
  INV_X1    g624(.A(new_n811_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n808_), .A2(new_n809_), .A3(KEYINPUT59), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n825_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(G127gat), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n829_), .B1(new_n645_), .B2(KEYINPUT120), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n830_), .B1(KEYINPUT120), .B2(new_n829_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n805_), .A2(new_n806_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(new_n814_), .A3(new_n807_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n808_), .A2(KEYINPUT116), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n645_), .A3(new_n834_), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n828_), .A2(new_n831_), .B1(new_n829_), .B2(new_n835_), .ZN(G1342gat));
  OAI211_X1 g635(.A(new_n567_), .B(new_n794_), .C1(new_n810_), .C2(new_n811_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(G134gat), .ZN(new_n838_));
  INV_X1    g637(.A(G134gat), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n815_), .A2(new_n839_), .A3(new_n624_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(G1343gat));
  NOR4_X1   g640(.A1(new_n607_), .A2(new_n389_), .A3(new_n738_), .A4(new_n354_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n832_), .A2(new_n431_), .A3(new_n842_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g643(.A1(new_n832_), .A2(new_n842_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n845_), .A2(new_n547_), .ZN(new_n846_));
  XOR2_X1   g645(.A(KEYINPUT121), .B(G148gat), .Z(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(G1345gat));
  NOR2_X1   g647(.A1(new_n845_), .A2(new_n582_), .ZN(new_n849_));
  XOR2_X1   g648(.A(KEYINPUT61), .B(G155gat), .Z(new_n850_));
  XNOR2_X1  g649(.A(new_n849_), .B(new_n850_), .ZN(G1346gat));
  INV_X1    g650(.A(new_n567_), .ZN(new_n852_));
  OAI21_X1  g651(.A(G162gat), .B1(new_n845_), .B2(new_n852_), .ZN(new_n853_));
  OR2_X1    g652(.A1(new_n590_), .A2(G162gat), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n845_), .B2(new_n854_), .ZN(G1347gat));
  AND2_X1   g654(.A1(new_n749_), .A2(new_n792_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n617_), .A2(new_n389_), .A3(new_n391_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n207_), .B1(new_n858_), .B2(new_n431_), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n859_), .A2(KEYINPUT62), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n858_), .A2(new_n300_), .A3(new_n431_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n859_), .A2(KEYINPUT62), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n860_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT122), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n860_), .A2(new_n865_), .A3(new_n861_), .A4(new_n862_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n866_), .ZN(G1348gat));
  AND3_X1   g666(.A1(new_n391_), .A2(new_n738_), .A3(new_n389_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n832_), .A2(G176gat), .A3(new_n546_), .A4(new_n868_), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n869_), .A2(KEYINPUT123), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(KEYINPUT123), .ZN(new_n871_));
  AOI21_X1  g670(.A(G176gat), .B1(new_n858_), .B2(new_n546_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n870_), .A2(new_n871_), .A3(new_n872_), .ZN(G1349gat));
  INV_X1    g672(.A(new_n858_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n874_), .A2(new_n221_), .A3(new_n582_), .ZN(new_n875_));
  AND3_X1   g674(.A1(new_n832_), .A2(new_n645_), .A3(new_n868_), .ZN(new_n876_));
  OR2_X1    g675(.A1(new_n876_), .A2(KEYINPUT124), .ZN(new_n877_));
  AOI21_X1  g676(.A(G183gat), .B1(new_n876_), .B2(KEYINPUT124), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n875_), .B1(new_n877_), .B2(new_n878_), .ZN(G1350gat));
  OAI21_X1  g678(.A(G190gat), .B1(new_n874_), .B2(new_n852_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n858_), .A2(new_n297_), .A3(new_n624_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1351gat));
  NAND2_X1  g681(.A1(KEYINPUT125), .A2(G197gat), .ZN(new_n883_));
  NOR4_X1   g682(.A1(new_n720_), .A2(new_n607_), .A3(new_n738_), .A4(new_n353_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n832_), .A2(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n883_), .B1(new_n885_), .B2(new_n430_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(KEYINPUT125), .A2(G197gat), .ZN(new_n887_));
  XOR2_X1   g686(.A(new_n887_), .B(KEYINPUT126), .Z(new_n888_));
  XNOR2_X1  g687(.A(new_n886_), .B(new_n888_), .ZN(G1352gat));
  AND2_X1   g688(.A1(new_n832_), .A2(new_n884_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n546_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n265_), .A2(KEYINPUT127), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(G1353gat));
  XNOR2_X1  g692(.A(KEYINPUT63), .B(G211gat), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n890_), .A2(new_n645_), .A3(new_n894_), .ZN(new_n895_));
  OAI22_X1  g694(.A1(new_n885_), .A2(new_n582_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(G1354gat));
  OAI21_X1  g696(.A(G218gat), .B1(new_n885_), .B2(new_n852_), .ZN(new_n898_));
  OR2_X1    g697(.A1(new_n590_), .A2(G218gat), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n885_), .B2(new_n899_), .ZN(G1355gat));
endmodule


