//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 0 0 1 0 0 0 0 0 1 1 0 1 0 0 0 0 1 0 0 1 1 0 0 1 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_;
  INV_X1    g000(.A(G141gat), .ZN(new_n202_));
  INV_X1    g001(.A(G148gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  AND2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT89), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT1), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT88), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n209_), .A2(KEYINPUT1), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n206_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n204_), .A2(KEYINPUT3), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n204_), .A2(KEYINPUT3), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n205_), .A2(KEYINPUT90), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n216_), .B(new_n217_), .C1(new_n218_), .C2(KEYINPUT2), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n218_), .A2(KEYINPUT2), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n209_), .B(new_n212_), .C1(new_n219_), .C2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n215_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT91), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT91), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n215_), .A2(new_n221_), .A3(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT29), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT95), .B(G204gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(G197gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT94), .B(G197gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(G204gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT21), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n230_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT96), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(G211gat), .B(G218gat), .Z(new_n237_));
  OAI22_X1  g036(.A1(G197gat), .A2(new_n229_), .B1(new_n231_), .B2(G204gat), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n237_), .B1(new_n238_), .B2(KEYINPUT21), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n236_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n230_), .A2(new_n232_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n241_), .A2(KEYINPUT21), .A3(new_n237_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G228gat), .A2(G233gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n242_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n246_), .B1(new_n236_), .B2(new_n239_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n247_), .B1(KEYINPUT29), .B2(new_n222_), .ZN(new_n248_));
  OAI22_X1  g047(.A1(new_n228_), .A2(new_n245_), .B1(new_n248_), .B2(new_n244_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G78gat), .B(G106gat), .ZN(new_n250_));
  XOR2_X1   g049(.A(new_n249_), .B(new_n250_), .Z(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n249_), .A2(new_n250_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT97), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n215_), .A2(new_n221_), .A3(new_n224_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n224_), .B1(new_n215_), .B2(new_n221_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n227_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT93), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT93), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n226_), .A2(new_n259_), .A3(new_n227_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(G22gat), .B(G50gat), .Z(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n258_), .A2(new_n260_), .A3(new_n262_), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n264_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n265_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n254_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n252_), .A2(new_n269_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n251_), .B(new_n254_), .C1(new_n267_), .C2(new_n268_), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G226gat), .A2(G233gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n276_));
  INV_X1    g075(.A(G169gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G183gat), .A2(G190gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT23), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT84), .B(G190gat), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n280_), .B1(G183gat), .B2(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n278_), .B1(new_n282_), .B2(KEYINPUT85), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n283_), .B1(KEYINPUT85), .B2(new_n282_), .ZN(new_n284_));
  OR3_X1    g083(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n280_), .A2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(G176gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n288_), .B1(new_n277_), .B2(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n291_), .B1(new_n281_), .B2(KEYINPUT26), .ZN(new_n292_));
  INV_X1    g091(.A(G183gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT25), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT83), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n293_), .A2(KEYINPUT83), .A3(KEYINPUT25), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT25), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(G183gat), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n296_), .A2(new_n297_), .A3(new_n299_), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n286_), .B(new_n290_), .C1(new_n292_), .C2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n284_), .A2(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n243_), .A2(new_n302_), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n294_), .A2(new_n299_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT26), .B(G190gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT99), .B1(new_n306_), .B2(new_n290_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n280_), .A2(new_n285_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n306_), .A2(KEYINPUT99), .A3(new_n290_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n278_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n280_), .B1(G183gat), .B2(G190gat), .ZN(new_n312_));
  AOI22_X1  g111(.A1(new_n309_), .A2(new_n310_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT20), .B1(new_n247_), .B2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n275_), .B1(new_n303_), .B2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G8gat), .B(G36gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT18), .ZN(new_n317_));
  XOR2_X1   g116(.A(G64gat), .B(G92gat), .Z(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n243_), .A2(new_n302_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT20), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n321_), .B1(new_n247_), .B2(new_n313_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n275_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n320_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  AND3_X1   g123(.A1(new_n315_), .A2(new_n319_), .A3(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n319_), .B1(new_n315_), .B2(new_n324_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n327_), .A2(KEYINPUT27), .ZN(new_n328_));
  NOR3_X1   g127(.A1(new_n303_), .A2(new_n314_), .A3(new_n275_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n323_), .B1(new_n320_), .B2(new_n322_), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n319_), .B(KEYINPUT102), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n325_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n333_), .A2(new_n334_), .A3(KEYINPUT27), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n328_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n272_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n302_), .B(KEYINPUT30), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT87), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G71gat), .B(G99gat), .ZN(new_n341_));
  INV_X1    g140(.A(G43gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT86), .B(G15gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G227gat), .A2(G233gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n345_), .B(new_n346_), .Z(new_n347_));
  NAND2_X1  g146(.A1(new_n340_), .A2(new_n347_), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n339_), .B(KEYINPUT87), .Z(new_n349_));
  OAI21_X1  g148(.A(new_n348_), .B1(new_n349_), .B2(new_n347_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G127gat), .B(G134gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G113gat), .B(G120gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n353_), .B(KEYINPUT31), .Z(new_n354_));
  XOR2_X1   g153(.A(new_n350_), .B(new_n354_), .Z(new_n355_));
  NOR3_X1   g154(.A1(new_n255_), .A2(new_n256_), .A3(new_n353_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n353_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n222_), .A2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT4), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G225gat), .A2(G233gat), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n223_), .A2(new_n225_), .A3(new_n357_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT4), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n359_), .A2(new_n361_), .A3(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n360_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G1gat), .B(G29gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT100), .B(KEYINPUT0), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  XOR2_X1   g169(.A(G57gat), .B(G85gat), .Z(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n367_), .A2(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n372_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n355_), .A2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n338_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n358_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n362_), .A2(new_n380_), .A3(new_n361_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n363_), .B1(new_n362_), .B2(new_n380_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n382_), .B1(new_n363_), .B2(new_n362_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n372_), .B(new_n381_), .C1(new_n383_), .C2(new_n361_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n327_), .B(new_n384_), .C1(KEYINPUT33), .C2(new_n374_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n374_), .A2(KEYINPUT33), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT101), .B1(new_n385_), .B2(new_n387_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n327_), .A2(new_n384_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT101), .ZN(new_n390_));
  OR2_X1    g189(.A1(new_n374_), .A2(KEYINPUT33), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n389_), .A2(new_n390_), .A3(new_n391_), .A4(new_n386_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n315_), .A2(new_n324_), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n319_), .A2(KEYINPUT32), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n395_), .B1(new_n331_), .B2(new_n394_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n376_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n388_), .A2(new_n392_), .A3(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n272_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n376_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n337_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n355_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n379_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT69), .ZN(new_n405_));
  NOR2_X1   g204(.A1(G99gat), .A2(G106gat), .ZN(new_n406_));
  NOR2_X1   g205(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  OAI22_X1  g207(.A1(KEYINPUT67), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  AND2_X1   g209(.A1(G99gat), .A2(G106gat), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT66), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n413_), .A2(KEYINPUT6), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n415_), .A2(KEYINPUT66), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n412_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(KEYINPUT66), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n413_), .A2(KEYINPUT6), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n419_), .A3(new_n411_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n410_), .B1(new_n417_), .B2(new_n420_), .ZN(new_n421_));
  XOR2_X1   g220(.A(G85gat), .B(G92gat), .Z(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n405_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n418_), .A2(new_n419_), .A3(new_n411_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n411_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  OAI211_X1 g226(.A(KEYINPUT69), .B(new_n422_), .C1(new_n427_), .C2(new_n410_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n424_), .A2(new_n428_), .A3(KEYINPUT8), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT70), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT70), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n424_), .A2(new_n428_), .A3(new_n431_), .A4(KEYINPUT8), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT68), .ZN(new_n433_));
  AOI211_X1 g232(.A(KEYINPUT8), .B(new_n423_), .C1(new_n421_), .C2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT68), .B1(new_n427_), .B2(new_n410_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n430_), .A2(new_n432_), .A3(new_n436_), .ZN(new_n437_));
  XOR2_X1   g236(.A(KEYINPUT10), .B(G99gat), .Z(new_n438_));
  INV_X1    g237(.A(G106gat), .ZN(new_n439_));
  AOI22_X1  g238(.A1(KEYINPUT9), .A2(new_n422_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(KEYINPUT65), .B(G85gat), .ZN(new_n441_));
  INV_X1    g240(.A(G92gat), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n442_), .A2(KEYINPUT9), .ZN(new_n443_));
  OAI221_X1 g242(.A(new_n440_), .B1(new_n425_), .B2(new_n426_), .C1(new_n441_), .C2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n437_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT71), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G29gat), .B(G36gat), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n447_), .A2(KEYINPUT73), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(KEYINPUT73), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G43gat), .B(G50gat), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n450_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT71), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n437_), .A2(new_n455_), .A3(new_n444_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n446_), .A2(new_n454_), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT74), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n446_), .A2(KEYINPUT74), .A3(new_n454_), .A4(new_n456_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n454_), .B(KEYINPUT15), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n445_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n459_), .A2(new_n460_), .A3(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT35), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G190gat), .B(G218gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT76), .ZN(new_n466_));
  XOR2_X1   g265(.A(G134gat), .B(G162gat), .Z(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  AOI22_X1  g268(.A1(new_n463_), .A2(new_n464_), .B1(KEYINPUT36), .B2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G232gat), .A2(G233gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT75), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n474_), .B1(new_n463_), .B2(new_n475_), .ZN(new_n476_));
  AOI22_X1  g275(.A1(new_n457_), .A2(new_n458_), .B1(new_n445_), .B2(new_n461_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n477_), .A2(KEYINPUT75), .A3(new_n460_), .A4(new_n473_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n470_), .A2(new_n476_), .A3(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n469_), .A2(KEYINPUT36), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n480_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n470_), .A2(new_n476_), .A3(new_n482_), .A4(new_n478_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n404_), .A2(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(G57gat), .B(G64gat), .Z(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT72), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT11), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G71gat), .B(G78gat), .Z(new_n491_));
  OR2_X1    g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n488_), .A2(new_n489_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n490_), .A2(new_n493_), .A3(new_n491_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n437_), .A2(new_n455_), .A3(new_n444_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n455_), .B1(new_n437_), .B2(new_n444_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n496_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT12), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G230gat), .A2(G233gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT64), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n446_), .A2(new_n495_), .A3(new_n456_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n445_), .A2(new_n496_), .A3(KEYINPUT12), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n501_), .A2(new_n504_), .A3(new_n505_), .A4(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n499_), .A2(new_n505_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(new_n503_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G120gat), .B(G148gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT5), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G176gat), .B(G204gat), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n512_), .B(new_n513_), .Z(new_n514_));
  NAND2_X1  g313(.A1(new_n510_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n514_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n507_), .A2(new_n509_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT13), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n515_), .A2(KEYINPUT13), .A3(new_n517_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G15gat), .B(G22gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(KEYINPUT77), .B(G8gat), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n524_), .A2(G1gat), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT14), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n523_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(G1gat), .B(G8gat), .Z(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n448_), .A2(new_n449_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n450_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n533_), .A2(KEYINPUT80), .A3(new_n451_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT80), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n535_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n530_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT81), .ZN(new_n538_));
  NOR3_X1   g337(.A1(new_n452_), .A2(new_n535_), .A3(new_n453_), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT80), .B1(new_n533_), .B2(new_n451_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n529_), .B(new_n538_), .C1(new_n539_), .C2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n536_), .A2(new_n534_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n538_), .B1(new_n543_), .B2(new_n529_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n537_), .B1(new_n542_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT82), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G229gat), .A2(G233gat), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n529_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT81), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n541_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n552_), .A2(KEYINPUT82), .A3(new_n537_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n547_), .A2(new_n549_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n461_), .A2(new_n530_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n552_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(new_n548_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n554_), .A2(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G113gat), .B(G141gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(G169gat), .B(G197gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n558_), .B(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n522_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n495_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(new_n530_), .ZN(new_n568_));
  XOR2_X1   g367(.A(G127gat), .B(G155gat), .Z(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G183gat), .B(G211gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT17), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n568_), .A2(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n573_), .B(KEYINPUT17), .Z(new_n576_));
  AOI21_X1  g375(.A(new_n575_), .B1(new_n568_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n565_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n486_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT104), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n486_), .A2(KEYINPUT104), .A3(new_n579_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(G1gat), .B1(new_n585_), .B2(new_n377_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT38), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT37), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n484_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n481_), .A2(KEYINPUT37), .A3(new_n483_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n591_), .A2(new_n578_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT79), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n404_), .A2(new_n565_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT103), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n593_), .A2(KEYINPUT103), .A3(new_n594_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n377_), .A2(G1gat), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n597_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT105), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n600_), .A2(new_n601_), .A3(new_n587_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n601_), .B1(new_n600_), .B2(new_n587_), .ZN(new_n603_));
  OAI221_X1 g402(.A(new_n586_), .B1(new_n587_), .B2(new_n600_), .C1(new_n602_), .C2(new_n603_), .ZN(G1324gat));
  NOR2_X1   g403(.A1(new_n337_), .A2(new_n524_), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n597_), .A2(new_n598_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT106), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n486_), .A2(new_n579_), .A3(new_n336_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(G8gat), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n608_), .B1(new_n610_), .B2(KEYINPUT39), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT39), .ZN(new_n612_));
  AOI211_X1 g411(.A(KEYINPUT106), .B(new_n612_), .C1(new_n609_), .C2(G8gat), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT107), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n615_), .B1(new_n610_), .B2(KEYINPUT39), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n609_), .A2(KEYINPUT107), .A3(new_n612_), .A4(G8gat), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n607_), .B(KEYINPUT40), .C1(new_n614_), .C2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT40), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n618_), .A2(new_n613_), .A3(new_n611_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n620_), .B1(new_n621_), .B2(new_n606_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n619_), .A2(new_n622_), .ZN(G1325gat));
  NAND2_X1  g422(.A1(new_n584_), .A2(new_n355_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(G15gat), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT108), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT108), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n624_), .A2(new_n627_), .A3(G15gat), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT41), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n597_), .A2(new_n598_), .ZN(new_n632_));
  INV_X1    g431(.A(G15gat), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n632_), .A2(new_n633_), .A3(new_n355_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n626_), .A2(KEYINPUT41), .A3(new_n628_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n631_), .A2(new_n634_), .A3(new_n635_), .ZN(G1326gat));
  INV_X1    g435(.A(G22gat), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n272_), .B(KEYINPUT109), .Z(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n637_), .B1(new_n584_), .B2(new_n639_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT42), .Z(new_n641_));
  NAND3_X1  g440(.A1(new_n632_), .A2(new_n637_), .A3(new_n639_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1327gat));
  AOI22_X1  g442(.A1(new_n398_), .A2(new_n272_), .B1(new_n400_), .B2(new_n337_), .ZN(new_n644_));
  OAI22_X1  g443(.A1(new_n644_), .A2(new_n355_), .B1(new_n338_), .B2(new_n378_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n484_), .A2(new_n577_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(new_n564_), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT111), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n645_), .A2(KEYINPUT111), .A3(new_n564_), .A4(new_n646_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(G29gat), .B1(new_n652_), .B2(new_n376_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT43), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n645_), .A2(new_n654_), .A3(new_n591_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT110), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n591_), .A2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n589_), .A2(KEYINPUT110), .A3(new_n590_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n404_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n655_), .B1(new_n659_), .B2(new_n654_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n565_), .A2(new_n577_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n660_), .A2(KEYINPUT44), .A3(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT44), .B1(new_n660_), .B2(new_n661_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n376_), .A2(G29gat), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n653_), .B1(new_n664_), .B2(new_n665_), .ZN(G1328gat));
  NOR2_X1   g465(.A1(new_n337_), .A2(G36gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n649_), .A2(new_n650_), .A3(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(KEYINPUT112), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT112), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n649_), .A2(new_n670_), .A3(new_n650_), .A4(new_n667_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n669_), .A2(KEYINPUT45), .A3(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT45), .B1(new_n669_), .B2(new_n671_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n662_), .A2(new_n663_), .A3(new_n337_), .ZN(new_n675_));
  INV_X1    g474(.A(G36gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n674_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT46), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n674_), .B(KEYINPUT46), .C1(new_n675_), .C2(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1329gat));
  NOR4_X1   g480(.A1(new_n662_), .A2(new_n663_), .A3(new_n342_), .A4(new_n403_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT47), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n342_), .B1(new_n651_), .B2(new_n403_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n683_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n685_), .ZN(new_n687_));
  OAI21_X1  g486(.A(KEYINPUT47), .B1(new_n682_), .B2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(G1330gat));
  AOI21_X1  g488(.A(G50gat), .B1(new_n652_), .B2(new_n639_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n272_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n691_), .A2(G50gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n690_), .B1(new_n664_), .B2(new_n692_), .ZN(G1331gat));
  INV_X1    g492(.A(new_n522_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n563_), .A2(new_n577_), .ZN(new_n695_));
  NOR4_X1   g494(.A1(new_n404_), .A2(new_n485_), .A3(new_n694_), .A4(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(G57gat), .A3(new_n376_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT114), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n404_), .A2(new_n562_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n699_), .A2(KEYINPUT113), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(KEYINPUT113), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n700_), .A2(new_n701_), .A3(new_n694_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n702_), .A2(new_n593_), .A3(new_n376_), .ZN(new_n703_));
  INV_X1    g502(.A(G57gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n698_), .B1(new_n703_), .B2(new_n704_), .ZN(G1332gat));
  NAND2_X1  g504(.A1(new_n696_), .A2(new_n336_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(G64gat), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n707_), .A2(KEYINPUT48), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(KEYINPUT48), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n702_), .A2(new_n593_), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n337_), .A2(G64gat), .ZN(new_n711_));
  OAI22_X1  g510(.A1(new_n708_), .A2(new_n709_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT115), .ZN(G1333gat));
  NAND2_X1  g512(.A1(new_n696_), .A2(new_n355_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(G71gat), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n715_), .A2(KEYINPUT49), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n715_), .A2(KEYINPUT49), .ZN(new_n717_));
  OR2_X1    g516(.A1(new_n403_), .A2(G71gat), .ZN(new_n718_));
  OAI22_X1  g517(.A1(new_n716_), .A2(new_n717_), .B1(new_n710_), .B2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT116), .ZN(G1334gat));
  INV_X1    g519(.A(G78gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n721_), .B1(new_n696_), .B2(new_n639_), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT50), .Z(new_n723_));
  NAND2_X1  g522(.A1(new_n639_), .A2(new_n721_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n723_), .B1(new_n710_), .B2(new_n724_), .ZN(G1335gat));
  AND2_X1   g524(.A1(new_n702_), .A2(new_n646_), .ZN(new_n726_));
  AOI21_X1  g525(.A(G85gat), .B1(new_n726_), .B2(new_n376_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n522_), .A2(new_n578_), .A3(new_n563_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT117), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n660_), .A2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT118), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n377_), .A2(new_n441_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n727_), .B1(new_n731_), .B2(new_n732_), .ZN(G1336gat));
  AOI21_X1  g532(.A(G92gat), .B1(new_n726_), .B2(new_n336_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n337_), .A2(new_n442_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n731_), .B2(new_n735_), .ZN(G1337gat));
  NAND3_X1  g535(.A1(new_n726_), .A2(new_n438_), .A3(new_n355_), .ZN(new_n737_));
  OAI21_X1  g536(.A(G99gat), .B1(new_n730_), .B2(new_n403_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT51), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT51), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n737_), .A2(new_n741_), .A3(new_n738_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(G1338gat));
  NAND4_X1  g542(.A1(new_n702_), .A2(new_n439_), .A3(new_n691_), .A4(new_n646_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n660_), .A2(new_n691_), .A3(new_n729_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n745_), .A2(new_n746_), .A3(G106gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n745_), .B2(G106gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g549(.A(KEYINPUT123), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT55), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT120), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n503_), .B2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n446_), .A2(new_n456_), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT12), .B1(new_n755_), .B2(new_n496_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n505_), .A2(new_n506_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n754_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n754_), .B1(new_n752_), .B2(new_n503_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n501_), .A2(new_n505_), .A3(new_n506_), .A4(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n758_), .A2(new_n760_), .A3(new_n514_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT56), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n758_), .A2(new_n760_), .A3(KEYINPUT56), .A4(new_n514_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n547_), .A2(new_n553_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n548_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n556_), .A2(new_n548_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n768_), .A2(new_n561_), .ZN(new_n769_));
  AOI22_X1  g568(.A1(new_n558_), .A2(new_n561_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n770_), .A2(new_n517_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT58), .B1(new_n765_), .B2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n765_), .A2(KEYINPUT58), .A3(new_n771_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n590_), .ZN(new_n775_));
  AOI21_X1  g574(.A(KEYINPUT37), .B1(new_n481_), .B2(new_n483_), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n773_), .B(new_n774_), .C1(new_n775_), .C2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT121), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n764_), .A2(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n495_), .B1(new_n446_), .B2(new_n456_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n505_), .B(new_n506_), .C1(new_n780_), .C2(KEYINPUT12), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n516_), .B1(new_n781_), .B2(new_n754_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n782_), .A2(KEYINPUT121), .A3(KEYINPUT56), .A4(new_n760_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n779_), .A2(new_n763_), .A3(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT122), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n562_), .A2(new_n517_), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n784_), .A2(new_n785_), .A3(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n785_), .B1(new_n784_), .B2(new_n786_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n518_), .A2(new_n770_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  NOR3_X1   g589(.A1(new_n787_), .A2(new_n788_), .A3(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n484_), .A2(KEYINPUT57), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n777_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n784_), .A2(new_n786_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT122), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n784_), .A2(new_n786_), .A3(new_n785_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n796_), .A3(new_n789_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT57), .B1(new_n797_), .B2(new_n484_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n751_), .B1(new_n793_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n800_), .B1(new_n791_), .B2(new_n485_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n792_), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n765_), .A2(KEYINPUT58), .A3(new_n771_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n803_), .A2(new_n772_), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n797_), .A2(new_n802_), .B1(new_n591_), .B2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n801_), .A2(new_n805_), .A3(KEYINPUT123), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n799_), .A2(new_n578_), .A3(new_n806_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n591_), .A2(new_n522_), .A3(new_n695_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(KEYINPUT119), .A2(KEYINPUT54), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  XOR2_X1   g609(.A(KEYINPUT119), .B(KEYINPUT54), .Z(new_n811_));
  OAI21_X1  g610(.A(new_n810_), .B1(new_n808_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n807_), .A2(new_n812_), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n338_), .A2(new_n403_), .A3(new_n377_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n813_), .A2(new_n562_), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(G113gat), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n814_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n818_), .A2(KEYINPUT59), .ZN(new_n819_));
  INV_X1    g618(.A(new_n812_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n577_), .B1(new_n801_), .B2(new_n805_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n819_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n563_), .A2(new_n816_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n818_), .B1(new_n807_), .B2(new_n812_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT59), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n822_), .B(new_n823_), .C1(new_n824_), .C2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n817_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT124), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT124), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n817_), .A2(new_n826_), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(G1340gat));
  NAND2_X1  g630(.A1(new_n813_), .A2(new_n814_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT59), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n833_), .A2(new_n522_), .A3(new_n822_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(G120gat), .ZN(new_n835_));
  INV_X1    g634(.A(G120gat), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n836_), .B1(new_n694_), .B2(KEYINPUT60), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n824_), .B(new_n837_), .C1(KEYINPUT60), .C2(new_n836_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n835_), .A2(new_n838_), .ZN(G1341gat));
  NAND3_X1  g638(.A1(new_n833_), .A2(new_n577_), .A3(new_n822_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(G127gat), .ZN(new_n841_));
  OR3_X1    g640(.A1(new_n832_), .A2(G127gat), .A3(new_n578_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(G1342gat));
  AOI21_X1  g642(.A(G134gat), .B1(new_n824_), .B2(new_n485_), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n844_), .A2(KEYINPUT125), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(KEYINPUT125), .ZN(new_n846_));
  OR2_X1    g645(.A1(new_n820_), .A2(new_n821_), .ZN(new_n847_));
  AOI22_X1  g646(.A1(new_n832_), .A2(KEYINPUT59), .B1(new_n847_), .B2(new_n819_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n591_), .A2(G134gat), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n845_), .A2(new_n846_), .B1(new_n848_), .B2(new_n849_), .ZN(G1343gat));
  NOR4_X1   g649(.A1(new_n272_), .A2(new_n355_), .A3(new_n377_), .A4(new_n336_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n813_), .A2(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n852_), .A2(new_n563_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(new_n202_), .ZN(G1344gat));
  NOR2_X1   g653(.A1(new_n852_), .A2(new_n694_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(new_n203_), .ZN(G1345gat));
  NAND3_X1  g655(.A1(new_n813_), .A2(new_n577_), .A3(new_n851_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT126), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n813_), .A2(KEYINPUT126), .A3(new_n577_), .A4(new_n851_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT61), .B(G155gat), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n859_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n861_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(G1346gat));
  INV_X1    g663(.A(G162gat), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n657_), .A2(new_n658_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n852_), .A2(new_n865_), .A3(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n813_), .A2(new_n485_), .A3(new_n851_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n865_), .B2(new_n869_), .ZN(G1347gat));
  NOR2_X1   g669(.A1(new_n378_), .A2(new_n337_), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n638_), .A2(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n847_), .A2(new_n562_), .A3(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(KEYINPUT62), .B1(new_n873_), .B2(KEYINPUT22), .ZN(new_n874_));
  OAI21_X1  g673(.A(G169gat), .B1(new_n873_), .B2(KEYINPUT62), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  OAI211_X1 g675(.A(KEYINPUT62), .B(G169gat), .C1(new_n873_), .C2(KEYINPUT22), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1348gat));
  NAND3_X1  g677(.A1(new_n847_), .A2(new_n522_), .A3(new_n872_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n691_), .B1(new_n807_), .B2(new_n812_), .ZN(new_n880_));
  AND3_X1   g679(.A1(new_n871_), .A2(G176gat), .A3(new_n522_), .ZN(new_n881_));
  AOI22_X1  g680(.A1(new_n879_), .A2(new_n289_), .B1(new_n880_), .B2(new_n881_), .ZN(G1349gat));
  NAND2_X1  g681(.A1(new_n847_), .A2(new_n872_), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n883_), .A2(new_n578_), .A3(new_n304_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n880_), .A2(new_n577_), .A3(new_n871_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n293_), .B2(new_n885_), .ZN(G1350gat));
  INV_X1    g685(.A(new_n591_), .ZN(new_n887_));
  OAI21_X1  g686(.A(G190gat), .B1(new_n883_), .B2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n485_), .A2(new_n305_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n883_), .B2(new_n889_), .ZN(G1351gat));
  NAND3_X1  g689(.A1(new_n403_), .A2(new_n400_), .A3(new_n336_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n891_), .B1(new_n807_), .B2(new_n812_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n562_), .ZN(new_n893_));
  XOR2_X1   g692(.A(KEYINPUT127), .B(G197gat), .Z(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1352gat));
  NAND2_X1  g694(.A1(new_n892_), .A2(new_n522_), .ZN(new_n896_));
  MUX2_X1   g695(.A(new_n229_), .B(G204gat), .S(new_n896_), .Z(G1353gat));
  INV_X1    g696(.A(new_n892_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(KEYINPUT63), .B(G211gat), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n898_), .A2(new_n578_), .A3(new_n899_), .ZN(new_n900_));
  AOI211_X1 g699(.A(KEYINPUT63), .B(G211gat), .C1(new_n892_), .C2(new_n577_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n900_), .A2(new_n901_), .ZN(G1354gat));
  OR3_X1    g701(.A1(new_n898_), .A2(G218gat), .A3(new_n484_), .ZN(new_n903_));
  OAI21_X1  g702(.A(G218gat), .B1(new_n898_), .B2(new_n887_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1355gat));
endmodule


