//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n871_, new_n872_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n921_, new_n922_, new_n923_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_, new_n940_;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G92gat), .Z(new_n202_));
  INV_X1    g001(.A(KEYINPUT9), .ZN(new_n203_));
  NAND3_X1  g002(.A1(new_n202_), .A2(new_n203_), .A3(G85gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT6), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(KEYINPUT10), .B(G99gat), .Z(new_n209_));
  INV_X1    g008(.A(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(G85gat), .B(G92gat), .Z(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT9), .ZN(new_n213_));
  NAND4_X1  g012(.A1(new_n204_), .A2(new_n208_), .A3(new_n211_), .A4(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT7), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n212_), .B1(new_n217_), .B2(new_n207_), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n218_), .A2(KEYINPUT8), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(KEYINPUT8), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n214_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G57gat), .B(G64gat), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n222_), .A2(KEYINPUT11), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(KEYINPUT11), .ZN(new_n224_));
  XOR2_X1   g023(.A(G71gat), .B(G78gat), .Z(new_n225_));
  NAND3_X1  g024(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n224_), .A2(new_n225_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n221_), .A2(new_n229_), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n228_), .B(new_n214_), .C1(new_n219_), .C2(new_n220_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT12), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G230gat), .A2(G233gat), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT12), .B1(new_n221_), .B2(new_n229_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n233_), .A2(new_n234_), .A3(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT65), .ZN(new_n238_));
  INV_X1    g037(.A(new_n234_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n232_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT12), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n241_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n242_), .A2(new_n235_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(new_n244_), .A3(new_n234_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n238_), .A2(new_n240_), .A3(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G120gat), .B(G148gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT5), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G176gat), .B(G204gat), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n248_), .B(new_n249_), .Z(new_n250_));
  OR2_X1    g049(.A1(new_n246_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n246_), .A2(new_n250_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n251_), .A2(KEYINPUT13), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT13), .B1(new_n251_), .B2(new_n252_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT66), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT66), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n258_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  XOR2_X1   g059(.A(G29gat), .B(G36gat), .Z(new_n261_));
  XOR2_X1   g060(.A(G43gat), .B(G50gat), .Z(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G15gat), .B(G22gat), .ZN(new_n265_));
  INV_X1    g064(.A(G1gat), .ZN(new_n266_));
  INV_X1    g065(.A(G8gat), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT14), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G1gat), .B(G8gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  OR2_X1    g070(.A1(new_n264_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n263_), .B(KEYINPUT15), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n273_), .B1(new_n271_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G229gat), .A2(G233gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n264_), .B(new_n271_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n276_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G113gat), .B(G141gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G169gat), .B(G197gat), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n281_), .B(new_n282_), .Z(new_n283_));
  NAND3_X1  g082(.A1(new_n277_), .A2(new_n280_), .A3(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n283_), .B1(new_n277_), .B2(new_n280_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT69), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n260_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G155gat), .B(G162gat), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n290_), .A2(KEYINPUT1), .ZN(new_n291_));
  INV_X1    g090(.A(G141gat), .ZN(new_n292_));
  INV_X1    g091(.A(G148gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G141gat), .A2(G148gat), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n294_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n291_), .A2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n292_), .A2(new_n293_), .A3(KEYINPUT3), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT3), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n300_), .B1(G141gat), .B2(G148gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n296_), .A2(KEYINPUT76), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT2), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT2), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n296_), .A2(KEYINPUT76), .A3(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n302_), .A2(new_n304_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT77), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n290_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n302_), .A2(new_n304_), .A3(KEYINPUT77), .A4(new_n306_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n298_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(G134gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(G127gat), .ZN(new_n313_));
  INV_X1    g112(.A(G127gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(G134gat), .ZN(new_n315_));
  AND3_X1   g114(.A1(new_n313_), .A2(new_n315_), .A3(KEYINPUT74), .ZN(new_n316_));
  AOI21_X1  g115(.A(KEYINPUT74), .B1(new_n313_), .B2(new_n315_), .ZN(new_n317_));
  XOR2_X1   g116(.A(G113gat), .B(G120gat), .Z(new_n318_));
  NOR3_X1   g117(.A1(new_n316_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G113gat), .B(G120gat), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT74), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n314_), .A2(G134gat), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n312_), .A2(G127gat), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n321_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n313_), .A2(new_n315_), .A3(KEYINPUT74), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n320_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT89), .B1(new_n319_), .B2(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n318_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n324_), .A2(new_n325_), .A3(new_n320_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT89), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n328_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n311_), .A2(KEYINPUT90), .A3(new_n327_), .A4(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n298_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n307_), .A2(new_n308_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n290_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(new_n335_), .A3(new_n310_), .ZN(new_n336_));
  AND4_X1   g135(.A1(new_n333_), .A2(new_n327_), .A3(new_n336_), .A4(new_n331_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT90), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n319_), .A2(new_n326_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n338_), .B1(new_n311_), .B2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n332_), .B1(new_n337_), .B2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT4), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G225gat), .A2(G233gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n336_), .A2(new_n333_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n339_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n347_), .A2(KEYINPUT4), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n342_), .A2(new_n344_), .A3(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n311_), .A2(new_n327_), .A3(new_n331_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n347_), .A2(new_n351_), .A3(new_n338_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n344_), .B1(new_n352_), .B2(new_n332_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n350_), .A2(new_n354_), .ZN(new_n355_));
  XOR2_X1   g154(.A(G1gat), .B(G29gat), .Z(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G57gat), .B(G85gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n355_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n350_), .A2(new_n360_), .A3(new_n354_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G8gat), .B(G36gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT18), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G64gat), .B(G92gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT32), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G226gat), .A2(G233gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT19), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT22), .B(G169gat), .ZN(new_n373_));
  INV_X1    g172(.A(G176gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G169gat), .A2(G176gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G183gat), .A2(G190gat), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT23), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  OR2_X1    g178(.A1(G183gat), .A2(G190gat), .ZN(new_n380_));
  NAND3_X1  g179(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n375_), .A2(new_n376_), .A3(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(G169gat), .A2(G176gat), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT24), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n386_), .B1(G169gat), .B2(G176gat), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT87), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n385_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n376_), .A2(new_n388_), .A3(KEYINPUT24), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT25), .B(G183gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT26), .B(G190gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n379_), .A2(new_n381_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n384_), .A2(new_n386_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n383_), .B1(new_n391_), .B2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT93), .ZN(new_n399_));
  OR2_X1    g198(.A1(KEYINPUT80), .A2(G197gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(KEYINPUT80), .A2(G197gat), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n400_), .A2(G204gat), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT82), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT82), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n400_), .A2(new_n404_), .A3(G204gat), .A4(new_n401_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(KEYINPUT81), .A2(G204gat), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(KEYINPUT81), .A2(G204gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(G197gat), .A3(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n403_), .A2(new_n405_), .A3(new_n409_), .ZN(new_n410_));
  XOR2_X1   g209(.A(G211gat), .B(G218gat), .Z(new_n411_));
  AND2_X1   g210(.A1(new_n411_), .A2(KEYINPUT21), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(G204gat), .ZN(new_n415_));
  AND2_X1   g214(.A1(KEYINPUT80), .A2(G197gat), .ZN(new_n416_));
  NOR2_X1   g215(.A1(KEYINPUT80), .A2(G197gat), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n415_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(G197gat), .ZN(new_n419_));
  AND2_X1   g218(.A1(KEYINPUT81), .A2(G204gat), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n419_), .B1(new_n420_), .B2(new_n406_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n418_), .A2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n411_), .B1(new_n422_), .B2(KEYINPUT21), .ZN(new_n423_));
  XOR2_X1   g222(.A(KEYINPUT83), .B(KEYINPUT21), .Z(new_n424_));
  NAND4_X1  g223(.A1(new_n403_), .A2(new_n424_), .A3(new_n405_), .A4(new_n409_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT84), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n423_), .A2(new_n425_), .A3(KEYINPUT84), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n414_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n399_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(KEYINPUT70), .A2(G169gat), .ZN(new_n432_));
  AOI21_X1  g231(.A(G176gat), .B1(new_n432_), .B2(KEYINPUT22), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT22), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n434_), .A2(KEYINPUT70), .A3(G169gat), .ZN(new_n435_));
  AOI22_X1  g234(.A1(new_n433_), .A2(new_n435_), .B1(G169gat), .B2(G176gat), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT71), .ZN(new_n437_));
  AOI22_X1  g236(.A1(new_n436_), .A2(new_n437_), .B1(new_n395_), .B2(new_n380_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(new_n437_), .B2(new_n436_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n397_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n387_), .A2(new_n385_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n439_), .A2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT20), .B1(new_n430_), .B2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n372_), .B1(new_n431_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n430_), .A2(new_n443_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n423_), .A2(new_n425_), .A3(KEYINPUT84), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT84), .B1(new_n423_), .B2(new_n425_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n413_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(new_n398_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n372_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n446_), .A2(new_n450_), .A3(KEYINPUT20), .A4(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n370_), .B1(new_n445_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n398_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n454_), .B(new_n413_), .C1(new_n447_), .C2(new_n448_), .ZN(new_n455_));
  OAI211_X1 g254(.A(new_n455_), .B(KEYINPUT20), .C1(new_n430_), .C2(new_n443_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n451_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n446_), .A2(new_n450_), .A3(KEYINPUT20), .A4(new_n372_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n453_), .B1(new_n459_), .B2(new_n370_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n364_), .A2(new_n460_), .ZN(new_n461_));
  AOI211_X1 g260(.A(new_n344_), .B(new_n348_), .C1(new_n341_), .C2(KEYINPUT4), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n341_), .A2(new_n344_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n361_), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT92), .B1(new_n462_), .B2(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n348_), .B1(new_n341_), .B2(KEYINPUT4), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n343_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT92), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n360_), .B1(new_n341_), .B2(new_n344_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n465_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n457_), .A2(new_n458_), .A3(new_n368_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT88), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n368_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n457_), .A2(new_n458_), .A3(new_n368_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n475_), .B1(new_n476_), .B2(KEYINPUT88), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n471_), .A2(new_n474_), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT33), .ZN(new_n479_));
  AND4_X1   g278(.A1(new_n479_), .A2(new_n350_), .A3(new_n360_), .A4(new_n354_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n353_), .B1(new_n466_), .B2(new_n344_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n479_), .B1(new_n481_), .B2(new_n360_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n461_), .B1(new_n478_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n345_), .A2(KEYINPUT29), .ZN(new_n485_));
  NAND2_X1  g284(.A1(KEYINPUT79), .A2(G233gat), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(KEYINPUT79), .A2(G233gat), .ZN(new_n488_));
  OAI21_X1  g287(.A(G228gat), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n449_), .A2(new_n485_), .A3(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n489_), .B1(new_n449_), .B2(new_n485_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G78gat), .B(G106gat), .ZN(new_n492_));
  NOR3_X1   g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n492_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n489_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT29), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n311_), .A2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n495_), .B1(new_n430_), .B2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n449_), .A2(new_n485_), .A3(new_n489_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n494_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n493_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT86), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n492_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT85), .ZN(new_n505_));
  XOR2_X1   g304(.A(KEYINPUT78), .B(KEYINPUT28), .Z(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n336_), .A2(new_n496_), .A3(new_n333_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G22gat), .B(G50gat), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n509_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n511_), .B1(new_n311_), .B2(new_n496_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n507_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n508_), .A2(new_n509_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n311_), .A2(new_n496_), .A3(new_n511_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(new_n506_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n513_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n503_), .B1(new_n505_), .B2(new_n518_), .ZN(new_n519_));
  AOI211_X1 g318(.A(KEYINPUT86), .B(new_n517_), .C1(new_n504_), .C2(KEYINPUT85), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n502_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT85), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n518_), .B1(new_n500_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT86), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n505_), .A2(new_n503_), .A3(new_n518_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n524_), .A2(new_n525_), .A3(new_n501_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n521_), .A2(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n364_), .B1(new_n521_), .B2(new_n526_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n475_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n457_), .A2(new_n458_), .A3(KEYINPUT88), .A4(new_n368_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n474_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT27), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n445_), .A2(new_n452_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(new_n368_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n475_), .A2(new_n532_), .ZN(new_n535_));
  AOI22_X1  g334(.A1(new_n531_), .A2(new_n532_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  AOI22_X1  g335(.A1(new_n484_), .A2(new_n527_), .B1(new_n528_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G227gat), .A2(G233gat), .ZN(new_n538_));
  INV_X1    g337(.A(G15gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(G71gat), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n541_), .B(G99gat), .Z(new_n542_));
  XOR2_X1   g341(.A(KEYINPUT72), .B(G43gat), .Z(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n439_), .A2(new_n442_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT30), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT73), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n544_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT75), .ZN(new_n550_));
  XOR2_X1   g349(.A(new_n339_), .B(KEYINPUT31), .Z(new_n551_));
  AOI21_X1  g350(.A(new_n549_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n551_), .A2(new_n550_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n546_), .A2(new_n547_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n554_), .A2(new_n544_), .A3(new_n548_), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n552_), .A2(new_n553_), .A3(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n553_), .B1(new_n552_), .B2(new_n555_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT94), .B1(new_n537_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT94), .ZN(new_n560_));
  INV_X1    g359(.A(new_n558_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n528_), .A2(new_n536_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n521_), .A2(new_n526_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n363_), .A2(KEYINPUT33), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n481_), .A2(new_n479_), .A3(new_n360_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n474_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(new_n567_), .A3(new_n471_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n563_), .B1(new_n568_), .B2(new_n461_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n560_), .B(new_n561_), .C1(new_n562_), .C2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n561_), .A2(new_n364_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n536_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n572_), .A2(new_n563_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n559_), .A2(new_n570_), .A3(new_n574_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n289_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n274_), .A2(new_n221_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT34), .ZN(new_n579_));
  OAI221_X1 g378(.A(new_n577_), .B1(KEYINPUT35), .B2(new_n579_), .C1(new_n264_), .C2(new_n221_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(KEYINPUT35), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n581_), .B(KEYINPUT67), .Z(new_n582_));
  XNOR2_X1  g381(.A(new_n580_), .B(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G190gat), .B(G218gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G134gat), .B(G162gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n586_), .A2(KEYINPUT36), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n586_), .A2(KEYINPUT36), .ZN(new_n588_));
  OR3_X1    g387(.A1(new_n583_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n583_), .A2(new_n587_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT37), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G231gat), .A2(G233gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n228_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT68), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n596_), .B(new_n271_), .Z(new_n597_));
  XOR2_X1   g396(.A(G127gat), .B(G155gat), .Z(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT16), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G183gat), .B(G211gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT17), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n601_), .A2(new_n602_), .ZN(new_n604_));
  OR3_X1    g403(.A1(new_n597_), .A2(new_n603_), .A3(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n597_), .A2(new_n603_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n593_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n576_), .A2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n611_), .A2(new_n266_), .A3(new_n364_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n612_), .A2(KEYINPUT95), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(KEYINPUT95), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT38), .ZN(new_n615_));
  OR3_X1    g414(.A1(new_n613_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n615_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n591_), .B(KEYINPUT96), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n618_), .A2(new_n607_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n576_), .A2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT97), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n621_), .A2(new_n364_), .ZN(new_n622_));
  OAI211_X1 g421(.A(new_n616_), .B(new_n617_), .C1(new_n266_), .C2(new_n622_), .ZN(G1324gat));
  NAND3_X1  g422(.A1(new_n611_), .A2(new_n267_), .A3(new_n572_), .ZN(new_n624_));
  OAI21_X1  g423(.A(G8gat), .B1(new_n620_), .B2(new_n536_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n625_), .A2(KEYINPUT39), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(KEYINPUT39), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n624_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g428(.A1(new_n611_), .A2(new_n539_), .A3(new_n558_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n621_), .A2(new_n558_), .ZN(new_n631_));
  XOR2_X1   g430(.A(KEYINPUT98), .B(KEYINPUT41), .Z(new_n632_));
  AND3_X1   g431(.A1(new_n631_), .A2(G15gat), .A3(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n632_), .B1(new_n631_), .B2(G15gat), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n630_), .B1(new_n633_), .B2(new_n634_), .ZN(G1326gat));
  INV_X1    g434(.A(G22gat), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n611_), .A2(new_n636_), .A3(new_n563_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n621_), .A2(new_n563_), .ZN(new_n638_));
  XOR2_X1   g437(.A(KEYINPUT99), .B(KEYINPUT42), .Z(new_n639_));
  AND3_X1   g438(.A1(new_n638_), .A2(G22gat), .A3(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n639_), .B1(new_n638_), .B2(G22gat), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n637_), .B1(new_n640_), .B2(new_n641_), .ZN(G1327gat));
  NAND2_X1  g441(.A1(new_n289_), .A2(new_n607_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT101), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n593_), .A2(KEYINPUT43), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n575_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n575_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n593_), .B1(new_n575_), .B2(KEYINPUT100), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT100), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n559_), .A2(new_n570_), .A3(new_n653_), .A4(new_n574_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n651_), .B1(new_n652_), .B2(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n644_), .B1(new_n650_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT44), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  OAI211_X1 g457(.A(KEYINPUT44), .B(new_n644_), .C1(new_n650_), .C2(new_n655_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n364_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G29gat), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n591_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n608_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n576_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n576_), .A2(KEYINPUT102), .A3(new_n664_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(G29gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(new_n670_), .A3(new_n364_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n662_), .A2(new_n671_), .ZN(G1328gat));
  NOR2_X1   g471(.A1(new_n536_), .A2(G36gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n667_), .A2(new_n668_), .A3(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT45), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n575_), .A2(KEYINPUT100), .ZN(new_n677_));
  INV_X1    g476(.A(new_n593_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n677_), .A2(new_n678_), .A3(new_n654_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(KEYINPUT43), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n575_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n681_), .A2(new_n647_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT44), .B1(new_n683_), .B2(new_n644_), .ZN(new_n684_));
  AOI211_X1 g483(.A(new_n657_), .B(new_n643_), .C1(new_n680_), .C2(new_n682_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n676_), .B1(new_n686_), .B2(new_n572_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n658_), .A2(new_n676_), .A3(new_n572_), .A4(new_n659_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(G36gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n675_), .B1(new_n687_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT46), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  OAI211_X1 g491(.A(KEYINPUT46), .B(new_n675_), .C1(new_n687_), .C2(new_n689_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1329gat));
  NAND3_X1  g493(.A1(new_n667_), .A2(new_n558_), .A3(new_n668_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n696_));
  XOR2_X1   g495(.A(KEYINPUT104), .B(G43gat), .Z(new_n697_));
  AND3_X1   g496(.A1(new_n695_), .A2(new_n696_), .A3(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n696_), .B1(new_n695_), .B2(new_n697_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n558_), .A2(G43gat), .ZN(new_n700_));
  OAI22_X1  g499(.A1(new_n698_), .A2(new_n699_), .B1(new_n660_), .B2(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g501(.A(G50gat), .B1(new_n669_), .B2(new_n563_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n563_), .A2(G50gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n686_), .B2(new_n704_), .ZN(G1331gat));
  INV_X1    g504(.A(G57gat), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n260_), .A2(new_n288_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n575_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n709_), .A2(new_n609_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n706_), .B1(new_n711_), .B2(new_n661_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n712_), .A2(KEYINPUT106), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n712_), .A2(KEYINPUT106), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n708_), .A2(new_n575_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n715_), .A2(KEYINPUT107), .A3(new_n619_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n717_));
  INV_X1    g516(.A(new_n619_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n717_), .B1(new_n709_), .B2(new_n718_), .ZN(new_n719_));
  XOR2_X1   g518(.A(KEYINPUT108), .B(G57gat), .Z(new_n720_));
  AND4_X1   g519(.A1(new_n364_), .A2(new_n716_), .A3(new_n719_), .A4(new_n720_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n713_), .A2(new_n714_), .A3(new_n721_), .ZN(G1332gat));
  NAND3_X1  g521(.A1(new_n716_), .A2(new_n572_), .A3(new_n719_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT48), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n723_), .A2(new_n724_), .A3(G64gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n723_), .B2(G64gat), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n536_), .A2(G64gat), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT109), .Z(new_n728_));
  OAI22_X1  g527(.A1(new_n725_), .A2(new_n726_), .B1(new_n711_), .B2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT110), .ZN(G1333gat));
  OR3_X1    g529(.A1(new_n711_), .A2(G71gat), .A3(new_n561_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n716_), .A2(new_n558_), .A3(new_n719_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT49), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n732_), .A2(new_n733_), .A3(G71gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n732_), .B2(G71gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n731_), .B1(new_n734_), .B2(new_n735_), .ZN(G1334gat));
  OR3_X1    g535(.A1(new_n711_), .A2(G78gat), .A3(new_n527_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n716_), .A2(new_n563_), .A3(new_n719_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n738_), .A2(G78gat), .A3(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n738_), .B2(G78gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n740_), .B2(new_n741_), .ZN(G1335gat));
  INV_X1    g541(.A(G85gat), .ZN(new_n743_));
  AOI211_X1 g542(.A(new_n608_), .B(new_n707_), .C1(new_n680_), .C2(new_n682_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n744_), .B2(new_n364_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n715_), .A2(new_n664_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n746_), .A2(G85gat), .A3(new_n661_), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n745_), .A2(new_n747_), .ZN(G1336gat));
  INV_X1    g547(.A(G92gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n749_), .B1(new_n746_), .B2(new_n536_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT112), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n572_), .A2(new_n202_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n744_), .B2(new_n752_), .ZN(G1337gat));
  NAND2_X1  g552(.A1(new_n558_), .A2(new_n209_), .ZN(new_n754_));
  OAI21_X1  g553(.A(KEYINPUT113), .B1(new_n746_), .B2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n744_), .A2(new_n558_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(G99gat), .ZN(new_n757_));
  XNOR2_X1  g556(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n757_), .B(new_n758_), .ZN(G1338gat));
  NOR3_X1   g558(.A1(new_n746_), .A2(G106gat), .A3(new_n527_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT115), .Z(new_n761_));
  AOI21_X1  g560(.A(new_n210_), .B1(new_n744_), .B2(new_n563_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT52), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n762_), .A2(KEYINPUT52), .ZN(new_n765_));
  OAI21_X1  g564(.A(KEYINPUT53), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n765_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n767_), .A2(new_n768_), .A3(new_n763_), .A4(new_n761_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n766_), .A2(new_n769_), .ZN(G1339gat));
  NAND3_X1  g569(.A1(new_n610_), .A2(new_n288_), .A3(new_n256_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT54), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n771_), .B(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT57), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n283_), .B1(new_n278_), .B2(new_n276_), .ZN(new_n775_));
  AOI22_X1  g574(.A1(new_n275_), .A2(new_n279_), .B1(new_n775_), .B2(KEYINPUT118), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n776_), .B1(KEYINPUT118), .B2(new_n775_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n777_), .A2(new_n284_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n779_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n251_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n782_));
  NOR4_X1   g581(.A1(new_n242_), .A2(new_n782_), .A3(new_n239_), .A4(new_n235_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT116), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n784_), .B1(new_n243_), .B2(new_n234_), .ZN(new_n785_));
  OAI211_X1 g584(.A(KEYINPUT116), .B(new_n239_), .C1(new_n242_), .C2(new_n235_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n783_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n238_), .A2(new_n782_), .A3(new_n245_), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n787_), .A2(KEYINPUT117), .A3(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT117), .B1(new_n787_), .B2(new_n788_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n250_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT56), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT117), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n233_), .A2(new_n236_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT116), .B1(new_n795_), .B2(new_n239_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n786_), .ZN(new_n797_));
  OAI22_X1  g596(.A1(new_n796_), .A2(new_n797_), .B1(new_n782_), .B2(new_n237_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n244_), .B1(new_n243_), .B2(new_n234_), .ZN(new_n799_));
  NOR4_X1   g598(.A1(new_n242_), .A2(KEYINPUT65), .A3(new_n239_), .A4(new_n235_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n799_), .A2(KEYINPUT55), .A3(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n794_), .B1(new_n798_), .B2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n787_), .A2(new_n788_), .A3(KEYINPUT117), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n804_), .A2(KEYINPUT56), .A3(new_n250_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n781_), .B1(new_n793_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n288_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n780_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n774_), .B1(new_n808_), .B2(new_n591_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT119), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT56), .B1(new_n804_), .B2(new_n250_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n250_), .ZN(new_n813_));
  AOI211_X1 g612(.A(new_n792_), .B(new_n813_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n251_), .B(new_n778_), .C1(new_n812_), .C2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT58), .ZN(new_n816_));
  OAI21_X1  g615(.A(KEYINPUT120), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n593_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n806_), .A2(new_n819_), .A3(KEYINPUT58), .A4(new_n778_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n817_), .A2(new_n818_), .A3(new_n820_), .ZN(new_n821_));
  AOI211_X1 g620(.A(new_n288_), .B(new_n781_), .C1(new_n793_), .C2(new_n805_), .ZN(new_n822_));
  OAI211_X1 g621(.A(KEYINPUT57), .B(new_n663_), .C1(new_n822_), .C2(new_n780_), .ZN(new_n823_));
  OAI211_X1 g622(.A(KEYINPUT119), .B(new_n774_), .C1(new_n808_), .C2(new_n591_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n811_), .A2(new_n821_), .A3(new_n823_), .A4(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n773_), .B1(new_n825_), .B2(new_n607_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n573_), .A2(new_n364_), .A3(new_n558_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(G113gat), .B1(new_n828_), .B2(new_n807_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n821_), .A2(new_n823_), .A3(new_n809_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n607_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT121), .ZN(new_n832_));
  INV_X1    g631(.A(new_n773_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT121), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n830_), .A2(new_n834_), .A3(new_n607_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n832_), .A2(new_n833_), .A3(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT59), .ZN(new_n837_));
  INV_X1    g636(.A(new_n827_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n836_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT59), .B1(new_n826_), .B2(new_n827_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(KEYINPUT122), .A3(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT122), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n836_), .A2(new_n842_), .A3(new_n837_), .A4(new_n838_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n807_), .A2(G113gat), .ZN(new_n845_));
  XOR2_X1   g644(.A(new_n845_), .B(KEYINPUT123), .Z(new_n846_));
  AOI21_X1  g645(.A(new_n829_), .B1(new_n844_), .B2(new_n846_), .ZN(G1340gat));
  INV_X1    g646(.A(G120gat), .ZN(new_n848_));
  INV_X1    g647(.A(new_n260_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(KEYINPUT60), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n828_), .B(new_n850_), .C1(KEYINPUT60), .C2(new_n848_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n849_), .B1(new_n841_), .B2(new_n843_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n852_), .B2(new_n848_), .ZN(G1341gat));
  NAND3_X1  g652(.A1(new_n828_), .A2(new_n314_), .A3(new_n608_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n607_), .B1(new_n841_), .B2(new_n843_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n314_), .ZN(G1342gat));
  NAND3_X1  g655(.A1(new_n828_), .A2(new_n312_), .A3(new_n618_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n593_), .B1(new_n841_), .B2(new_n843_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n312_), .ZN(G1343gat));
  NOR2_X1   g658(.A1(new_n826_), .A2(new_n558_), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n527_), .A2(new_n572_), .A3(new_n661_), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT124), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT124), .ZN(new_n863_));
  INV_X1    g662(.A(new_n861_), .ZN(new_n864_));
  NOR4_X1   g663(.A1(new_n826_), .A2(new_n863_), .A3(new_n558_), .A4(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n807_), .B1(new_n862_), .B2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(G141gat), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n292_), .B(new_n807_), .C1(new_n862_), .C2(new_n865_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1344gat));
  OAI21_X1  g668(.A(new_n260_), .B1(new_n862_), .B2(new_n865_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(G148gat), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n293_), .B(new_n260_), .C1(new_n862_), .C2(new_n865_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1345gat));
  OAI21_X1  g672(.A(new_n608_), .B1(new_n862_), .B2(new_n865_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(KEYINPUT61), .B(G155gat), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n875_), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n608_), .B(new_n877_), .C1(new_n862_), .C2(new_n865_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(G1346gat));
  INV_X1    g678(.A(G162gat), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n880_), .B(new_n618_), .C1(new_n862_), .C2(new_n865_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n862_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n865_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n593_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n881_), .B1(new_n884_), .B2(new_n880_), .ZN(G1347gat));
  INV_X1    g684(.A(KEYINPUT62), .ZN(new_n886_));
  INV_X1    g685(.A(G169gat), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n571_), .A2(new_n572_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(new_n563_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n773_), .B1(new_n831_), .B2(KEYINPUT121), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n835_), .ZN(new_n892_));
  AOI211_X1 g691(.A(KEYINPUT125), .B(new_n887_), .C1(new_n892_), .C2(new_n807_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT125), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n836_), .A2(new_n807_), .A3(new_n889_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(G169gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n886_), .B1(new_n893_), .B2(new_n896_), .ZN(new_n897_));
  AOI211_X1 g696(.A(new_n288_), .B(new_n890_), .C1(new_n891_), .C2(new_n835_), .ZN(new_n898_));
  OAI21_X1  g697(.A(KEYINPUT125), .B1(new_n898_), .B2(new_n887_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n895_), .A2(new_n894_), .A3(G169gat), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n899_), .A2(KEYINPUT62), .A3(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n898_), .A2(new_n373_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n897_), .A2(new_n901_), .A3(new_n902_), .ZN(G1348gat));
  AOI21_X1  g702(.A(G176gat), .B1(new_n892_), .B2(new_n260_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n260_), .A2(G176gat), .ZN(new_n905_));
  NOR4_X1   g704(.A1(new_n826_), .A2(new_n563_), .A3(new_n888_), .A4(new_n905_), .ZN(new_n906_));
  OR3_X1    g705(.A1(new_n904_), .A2(new_n906_), .A3(KEYINPUT126), .ZN(new_n907_));
  OAI21_X1  g706(.A(KEYINPUT126), .B1(new_n904_), .B2(new_n906_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1349gat));
  INV_X1    g708(.A(new_n392_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n892_), .A2(new_n910_), .A3(new_n608_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT127), .ZN(new_n912_));
  AND2_X1   g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n826_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(new_n527_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n571_), .A2(new_n572_), .A3(new_n608_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n917_), .A2(G183gat), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n911_), .A2(new_n912_), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n913_), .A2(new_n918_), .A3(new_n919_), .ZN(G1350gat));
  INV_X1    g719(.A(new_n892_), .ZN(new_n921_));
  OAI21_X1  g720(.A(G190gat), .B1(new_n921_), .B2(new_n593_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n892_), .A2(new_n393_), .A3(new_n618_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(G1351gat));
  NAND2_X1  g723(.A1(new_n914_), .A2(new_n561_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n572_), .A2(new_n528_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n925_), .A2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(new_n807_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(G197gat), .ZN(G1352gat));
  NAND4_X1  g728(.A1(new_n860_), .A2(new_n260_), .A3(new_n572_), .A4(new_n528_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n930_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n931_), .B1(new_n415_), .B2(new_n930_), .ZN(G1353gat));
  NOR3_X1   g731(.A1(new_n925_), .A2(new_n607_), .A3(new_n926_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n934_));
  AND2_X1   g733(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n933_), .B1(new_n934_), .B2(new_n935_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n936_), .B1(new_n933_), .B2(new_n934_), .ZN(G1354gat));
  INV_X1    g736(.A(G218gat), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n927_), .A2(new_n938_), .A3(new_n618_), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n925_), .A2(new_n593_), .A3(new_n926_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n938_), .B2(new_n940_), .ZN(G1355gat));
endmodule


