//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 1 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n617_,
    new_n618_, new_n619_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n854_, new_n855_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_;
  INV_X1    g000(.A(KEYINPUT101), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT13), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G230gat), .A2(G233gat), .ZN(new_n204_));
  INV_X1    g003(.A(G64gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G57gat), .ZN(new_n206_));
  INV_X1    g005(.A(G57gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G64gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT11), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n210_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G71gat), .B(G78gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(KEYINPUT68), .B1(new_n212_), .B2(new_n214_), .ZN(new_n215_));
  AOI21_X1  g014(.A(KEYINPUT11), .B1(new_n206_), .B2(new_n208_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT68), .ZN(new_n217_));
  NOR3_X1   g016(.A1(new_n216_), .A2(new_n217_), .A3(new_n213_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n211_), .B1(new_n215_), .B2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n212_), .A2(KEYINPUT68), .A3(new_n214_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n217_), .B1(new_n216_), .B2(new_n213_), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n220_), .B(new_n221_), .C1(new_n210_), .C2(new_n209_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n219_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G99gat), .A2(G106gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G99gat), .A2(G106gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT6), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n231_));
  OAI22_X1  g030(.A1(KEYINPUT66), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n227_), .A2(new_n230_), .A3(new_n231_), .A4(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(G85gat), .ZN(new_n234_));
  INV_X1    g033(.A(G92gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G85gat), .A2(G92gat), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n233_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT8), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(G85gat), .B1(KEYINPUT65), .B2(G92gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT65), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n242_), .B1(new_n243_), .B2(new_n235_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT9), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT64), .B(G106gat), .ZN(new_n247_));
  OR2_X1    g046(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n247_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n230_), .A2(new_n231_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n236_), .A2(new_n243_), .A3(KEYINPUT9), .A4(new_n237_), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n246_), .A2(new_n250_), .A3(new_n251_), .A4(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n233_), .A2(KEYINPUT8), .A3(new_n238_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n241_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n224_), .A2(KEYINPUT12), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(KEYINPUT67), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n241_), .A2(new_n258_), .A3(new_n253_), .A4(new_n254_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n257_), .A2(new_n223_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n256_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  AND3_X1   g061(.A1(new_n233_), .A2(KEYINPUT8), .A3(new_n238_), .ZN(new_n263_));
  AOI21_X1  g062(.A(KEYINPUT8), .B1(new_n233_), .B2(new_n238_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n258_), .B1(new_n265_), .B2(new_n253_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n259_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n224_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT12), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT69), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n223_), .B1(new_n257_), .B2(new_n259_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n272_));
  NOR3_X1   g071(.A1(new_n271_), .A2(new_n272_), .A3(KEYINPUT12), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n204_), .B(new_n262_), .C1(new_n270_), .C2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n268_), .A2(new_n260_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n204_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G120gat), .B(G148gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT5), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G176gat), .B(G204gat), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n279_), .B(new_n280_), .Z(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n274_), .A2(new_n277_), .A3(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT70), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n274_), .A2(new_n277_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n281_), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n284_), .A2(KEYINPUT71), .A3(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT71), .B1(new_n284_), .B2(new_n286_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n203_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n284_), .A2(new_n286_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n284_), .A2(KEYINPUT71), .A3(new_n286_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n292_), .A2(KEYINPUT13), .A3(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n289_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G15gat), .B(G22gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G1gat), .A2(G8gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT14), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n296_), .B1(new_n298_), .B2(KEYINPUT77), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n298_), .A2(KEYINPUT77), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G1gat), .B(G8gat), .ZN(new_n301_));
  OR3_X1    g100(.A1(new_n299_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n301_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G29gat), .B(G36gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G43gat), .B(G50gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  AND3_X1   g105(.A1(new_n302_), .A2(new_n303_), .A3(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n302_), .A2(new_n303_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n306_), .B(KEYINPUT15), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n307_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G229gat), .A2(G233gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n308_), .B(new_n306_), .Z(new_n314_));
  OAI21_X1  g113(.A(new_n313_), .B1(new_n311_), .B2(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(G113gat), .B(G141gat), .Z(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT80), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n317_), .B(KEYINPUT81), .Z(new_n318_));
  XNOR2_X1  g117(.A(G169gat), .B(G197gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n315_), .B(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n202_), .B1(new_n295_), .B2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G232gat), .A2(G233gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT73), .B(KEYINPUT35), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n309_), .A2(new_n255_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT74), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n257_), .A2(new_n306_), .A3(new_n259_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n327_), .A2(new_n328_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n329_), .B1(new_n331_), .B2(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(new_n329_), .B(KEYINPUT76), .Z(new_n336_));
  NAND4_X1  g135(.A1(new_n336_), .A2(new_n332_), .A3(new_n333_), .A4(new_n330_), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G190gat), .B(G218gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT75), .ZN(new_n340_));
  XOR2_X1   g139(.A(G134gat), .B(G162gat), .Z(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT36), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n342_), .A2(new_n343_), .ZN(new_n345_));
  NOR3_X1   g144(.A1(new_n338_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n338_), .A2(new_n344_), .ZN(new_n347_));
  OR2_X1    g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G169gat), .A2(G176gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT24), .ZN(new_n351_));
  NOR2_X1   g150(.A1(G169gat), .A2(G176gat), .ZN(new_n352_));
  MUX2_X1   g151(.A(new_n351_), .B(KEYINPUT24), .S(new_n352_), .Z(new_n353_));
  NAND2_X1  g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT23), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT25), .B(G183gat), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n356_), .A2(KEYINPUT82), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT26), .B(G190gat), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT82), .ZN(new_n359_));
  INV_X1    g158(.A(G183gat), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n360_), .A2(KEYINPUT25), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n358_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n353_), .B(new_n355_), .C1(new_n357_), .C2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n355_), .B1(G183gat), .B2(G190gat), .ZN(new_n364_));
  INV_X1    g163(.A(G176gat), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT22), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT83), .B1(new_n366_), .B2(G169gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT22), .B(G169gat), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n365_), .B(new_n367_), .C1(new_n368_), .C2(KEYINPUT83), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n364_), .A2(new_n369_), .A3(new_n350_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n363_), .A2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT30), .ZN(new_n372_));
  XOR2_X1   g171(.A(G71gat), .B(G99gat), .Z(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(G43gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G227gat), .A2(G233gat), .ZN(new_n375_));
  INV_X1    g174(.A(G15gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n374_), .B(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n372_), .B(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT84), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  XOR2_X1   g180(.A(G127gat), .B(G134gat), .Z(new_n382_));
  XNOR2_X1  g181(.A(G113gat), .B(G120gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n384_), .B(KEYINPUT31), .Z(new_n385_));
  NOR2_X1   g184(.A1(new_n381_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n379_), .A2(new_n380_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n379_), .A2(new_n380_), .A3(new_n385_), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G226gat), .A2(G233gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT19), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n368_), .A2(new_n365_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n350_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT93), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n393_), .A2(KEYINPUT93), .A3(new_n350_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n396_), .A2(new_n364_), .A3(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n356_), .A2(new_n358_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n353_), .A2(new_n355_), .A3(new_n399_), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(G197gat), .ZN(new_n402_));
  INV_X1    g201(.A(G204gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G197gat), .A2(G204gat), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n404_), .A2(KEYINPUT21), .A3(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G211gat), .B(G218gat), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n404_), .A2(new_n405_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT21), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT92), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n411_), .A2(KEYINPUT92), .A3(new_n406_), .A4(new_n407_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n408_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT20), .B1(new_n401_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n416_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n418_), .A2(new_n371_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n392_), .B1(new_n417_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n401_), .A2(new_n416_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n418_), .A2(new_n371_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n392_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n421_), .A2(new_n422_), .A3(KEYINPUT20), .A4(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G8gat), .B(G36gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT18), .ZN(new_n426_));
  XOR2_X1   g225(.A(G64gat), .B(G92gat), .Z(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT32), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n420_), .A2(new_n424_), .A3(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n423_), .B1(new_n417_), .B2(new_n419_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n421_), .A2(KEYINPUT20), .A3(new_n422_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n431_), .B1(new_n423_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G141gat), .A2(G148gat), .ZN(new_n434_));
  INV_X1    g233(.A(G141gat), .ZN(new_n435_));
  INV_X1    g234(.A(G148gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G155gat), .A2(G162gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT1), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT85), .ZN(new_n440_));
  INV_X1    g239(.A(G155gat), .ZN(new_n441_));
  INV_X1    g240(.A(G162gat), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT85), .B1(G155gat), .B2(G162gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n434_), .B(new_n437_), .C1(new_n439_), .C2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n435_), .A2(new_n436_), .A3(KEYINPUT86), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT3), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n434_), .A2(KEYINPUT2), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT2), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n450_), .A2(G141gat), .A3(G148gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n449_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT3), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n453_), .A2(new_n435_), .A3(new_n436_), .A4(KEYINPUT86), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n448_), .A2(new_n452_), .A3(new_n454_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n443_), .A2(new_n444_), .A3(new_n438_), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n455_), .A2(KEYINPUT87), .A3(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(KEYINPUT87), .B1(new_n455_), .B2(new_n456_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n446_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT88), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT88), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n461_), .B(new_n446_), .C1(new_n457_), .C2(new_n458_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n460_), .A2(new_n384_), .A3(new_n462_), .ZN(new_n463_));
  OR2_X1    g262(.A1(new_n463_), .A2(KEYINPUT4), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G225gat), .A2(G233gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT94), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n459_), .A2(new_n384_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n463_), .A2(KEYINPUT4), .A3(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n464_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n463_), .A2(new_n465_), .A3(new_n467_), .ZN(new_n470_));
  XOR2_X1   g269(.A(G1gat), .B(G29gat), .Z(new_n471_));
  XNOR2_X1  g270(.A(G57gat), .B(G85gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n474_));
  XOR2_X1   g273(.A(new_n473_), .B(new_n474_), .Z(new_n475_));
  NAND3_X1  g274(.A1(new_n469_), .A2(new_n470_), .A3(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n475_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n478_));
  OAI221_X1 g277(.A(new_n430_), .B1(new_n433_), .B2(new_n429_), .C1(new_n477_), .C2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT33), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n476_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n420_), .A2(new_n424_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(new_n428_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n469_), .A2(KEYINPUT33), .A3(new_n470_), .A4(new_n475_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n464_), .A2(new_n465_), .A3(new_n468_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n475_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n463_), .A2(new_n467_), .A3(new_n466_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n485_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n481_), .A2(new_n483_), .A3(new_n484_), .A4(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(KEYINPUT89), .B(KEYINPUT28), .Z(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G78gat), .B(G106gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G228gat), .A2(G233gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT91), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n418_), .A2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n460_), .A2(KEYINPUT29), .A3(new_n462_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT90), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n460_), .A2(KEYINPUT90), .A3(KEYINPUT29), .A4(new_n462_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n495_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n459_), .A2(KEYINPUT29), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n493_), .B1(new_n501_), .B2(new_n418_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n492_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NOR3_X1   g303(.A1(new_n500_), .A2(new_n502_), .A3(new_n492_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n491_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n460_), .A2(new_n462_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT29), .ZN(new_n508_));
  XOR2_X1   g307(.A(G22gat), .B(G50gat), .Z(new_n509_));
  NAND3_X1  g308(.A1(new_n507_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n509_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n500_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n502_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n492_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(new_n503_), .A3(new_n490_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n506_), .A2(new_n513_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n513_), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n517_), .A2(new_n503_), .A3(new_n490_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n490_), .B1(new_n517_), .B2(new_n503_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n520_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  AOI221_X4 g322(.A(new_n390_), .B1(new_n479_), .B2(new_n489_), .C1(new_n519_), .C2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(KEYINPUT97), .B(KEYINPUT27), .Z(new_n526_));
  NOR2_X1   g325(.A1(new_n483_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n420_), .A2(new_n428_), .A3(new_n424_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n528_), .A2(KEYINPUT27), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n529_), .B1(new_n428_), .B2(new_n433_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT96), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n529_), .B(KEYINPUT96), .C1(new_n428_), .C2(new_n433_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n527_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n477_), .A2(new_n478_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n388_), .A2(new_n389_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n523_), .A2(new_n538_), .A3(new_n519_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n538_), .B1(new_n523_), .B2(new_n519_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n537_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n349_), .B1(new_n525_), .B2(new_n542_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n289_), .A2(new_n294_), .A3(KEYINPUT101), .A4(new_n322_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G231gat), .A2(G233gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n308_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(new_n224_), .ZN(new_n547_));
  XOR2_X1   g346(.A(G127gat), .B(G155gat), .Z(new_n548_));
  XNOR2_X1  g347(.A(G183gat), .B(G211gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT17), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n547_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n547_), .A2(KEYINPUT17), .A3(new_n552_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n324_), .A2(new_n543_), .A3(new_n544_), .A4(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(G1gat), .B1(new_n558_), .B2(new_n535_), .ZN(new_n559_));
  NOR3_X1   g358(.A1(new_n521_), .A2(new_n522_), .A3(new_n520_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n513_), .B1(new_n506_), .B2(new_n518_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n390_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n536_), .B1(new_n562_), .B2(new_n539_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n322_), .B1(new_n563_), .B2(new_n524_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT98), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n289_), .A2(new_n294_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT37), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n348_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n556_), .B(KEYINPUT79), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  OAI211_X1 g370(.A(KEYINPUT98), .B(new_n322_), .C1(new_n563_), .C2(new_n524_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n566_), .A2(new_n567_), .A3(new_n571_), .A4(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT99), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n572_), .A2(new_n567_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n576_), .A2(KEYINPUT99), .A3(new_n571_), .A4(new_n566_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n575_), .A2(new_n577_), .A3(KEYINPUT100), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(KEYINPUT100), .B1(new_n575_), .B2(new_n577_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT38), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n535_), .A2(G1gat), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n581_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n582_), .B1(new_n581_), .B2(new_n583_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n559_), .B1(new_n584_), .B2(new_n585_), .ZN(G1324gat));
  INV_X1    g385(.A(KEYINPUT40), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n575_), .A2(new_n577_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT100), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n534_), .A2(G8gat), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n590_), .A2(new_n578_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT103), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n324_), .A2(new_n544_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n532_), .A2(new_n533_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n527_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n594_), .A2(new_n557_), .A3(new_n597_), .A4(new_n543_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT102), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT39), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n598_), .A2(new_n599_), .A3(new_n600_), .A4(G8gat), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n600_), .B(G8gat), .C1(new_n558_), .C2(new_n534_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT102), .ZN(new_n603_));
  OAI21_X1  g402(.A(G8gat), .B1(new_n558_), .B2(new_n534_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT39), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n601_), .A2(new_n603_), .A3(new_n605_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n592_), .A2(new_n593_), .A3(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n593_), .B1(new_n592_), .B2(new_n606_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n587_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n591_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n579_), .A2(new_n580_), .A3(new_n610_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n601_), .A2(new_n603_), .A3(new_n605_), .ZN(new_n612_));
  OAI21_X1  g411(.A(KEYINPUT103), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n592_), .A2(new_n593_), .A3(new_n606_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n613_), .A2(KEYINPUT40), .A3(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n609_), .A2(new_n615_), .ZN(G1325gat));
  OAI21_X1  g415(.A(G15gat), .B1(new_n558_), .B2(new_n538_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT41), .Z(new_n618_));
  NAND2_X1  g417(.A1(new_n390_), .A2(new_n376_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n618_), .B1(new_n588_), .B2(new_n619_), .ZN(G1326gat));
  NOR2_X1   g419(.A1(new_n560_), .A2(new_n561_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(G22gat), .B1(new_n558_), .B2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT42), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n622_), .A2(G22gat), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n624_), .B1(new_n588_), .B2(new_n625_), .ZN(G1327gat));
  OAI21_X1  g425(.A(new_n569_), .B1(new_n563_), .B2(new_n524_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT43), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(new_n594_), .A3(new_n570_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT44), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n535_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n629_), .A2(new_n630_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n631_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT104), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(G29gat), .B1(new_n634_), .B2(new_n635_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n349_), .A2(new_n570_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n576_), .A2(new_n566_), .A3(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n535_), .A2(G29gat), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT105), .Z(new_n642_));
  OAI22_X1  g441(.A1(new_n636_), .A2(new_n637_), .B1(new_n640_), .B2(new_n642_), .ZN(G1328gat));
  NAND3_X1  g442(.A1(new_n631_), .A2(new_n597_), .A3(new_n633_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(G36gat), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n534_), .A2(G36gat), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n640_), .A2(new_n646_), .ZN(new_n647_));
  XOR2_X1   g446(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n648_));
  XOR2_X1   g447(.A(new_n647_), .B(new_n648_), .Z(new_n649_));
  NAND2_X1  g448(.A1(new_n645_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT46), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n645_), .A2(new_n649_), .A3(KEYINPUT46), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1329gat));
  NAND3_X1  g453(.A1(new_n631_), .A2(new_n390_), .A3(new_n633_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(G43gat), .ZN(new_n656_));
  OR3_X1    g455(.A1(new_n640_), .A2(G43gat), .A3(new_n538_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT47), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n656_), .A2(KEYINPUT47), .A3(new_n657_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1330gat));
  NAND3_X1  g461(.A1(new_n631_), .A2(new_n621_), .A3(new_n633_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(G50gat), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n622_), .A2(G50gat), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT107), .Z(new_n666_));
  OAI21_X1  g465(.A(new_n664_), .B1(new_n640_), .B2(new_n666_), .ZN(G1331gat));
  AOI21_X1  g466(.A(new_n322_), .B1(new_n525_), .B2(new_n542_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT108), .ZN(new_n669_));
  OR2_X1    g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n669_), .ZN(new_n671_));
  AND4_X1   g470(.A1(new_n295_), .A2(new_n670_), .A3(new_n571_), .A4(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n672_), .A2(new_n207_), .A3(new_n632_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n295_), .A2(new_n323_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n570_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n675_), .A2(new_n543_), .A3(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(G57gat), .B1(new_n678_), .B2(new_n535_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n673_), .A2(new_n679_), .ZN(G1332gat));
  AOI21_X1  g479(.A(new_n205_), .B1(new_n677_), .B2(new_n597_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT48), .Z(new_n682_));
  NAND3_X1  g481(.A1(new_n672_), .A2(new_n205_), .A3(new_n597_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1333gat));
  INV_X1    g483(.A(G71gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n685_), .B1(new_n677_), .B2(new_n390_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT49), .Z(new_n687_));
  NAND3_X1  g486(.A1(new_n672_), .A2(new_n685_), .A3(new_n390_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1334gat));
  INV_X1    g488(.A(G78gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n690_), .B1(new_n677_), .B2(new_n621_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n691_), .B(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n672_), .A2(new_n690_), .A3(new_n621_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1335gat));
  NAND3_X1  g494(.A1(new_n628_), .A2(new_n570_), .A3(new_n675_), .ZN(new_n696_));
  OAI21_X1  g495(.A(G85gat), .B1(new_n696_), .B2(new_n535_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n670_), .A2(new_n295_), .A3(new_n639_), .A4(new_n671_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n632_), .A2(new_n234_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n697_), .B1(new_n698_), .B2(new_n699_), .ZN(G1336gat));
  INV_X1    g499(.A(new_n698_), .ZN(new_n701_));
  AOI21_X1  g500(.A(G92gat), .B1(new_n701_), .B2(new_n597_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n696_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n534_), .A2(new_n235_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT110), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n702_), .B1(new_n703_), .B2(new_n705_), .ZN(G1337gat));
  NAND4_X1  g505(.A1(new_n701_), .A2(new_n248_), .A3(new_n249_), .A4(new_n390_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n628_), .A2(new_n390_), .A3(new_n570_), .A4(new_n675_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT111), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n708_), .A2(new_n709_), .A3(G99gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n708_), .B2(G99gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND2_X1  g512(.A1(new_n621_), .A2(new_n247_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n698_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT112), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n715_), .B(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G106gat), .B1(new_n696_), .B2(new_n622_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT52), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n719_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n717_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n722_));
  XOR2_X1   g521(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n723_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n717_), .A2(new_n721_), .A3(new_n720_), .A4(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1339gat));
  NAND2_X1  g526(.A1(new_n322_), .A2(G113gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n567_), .A2(new_n571_), .A3(new_n323_), .ZN(new_n729_));
  XOR2_X1   g528(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n730_));
  XNOR2_X1  g529(.A(new_n729_), .B(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n315_), .A2(new_n321_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n314_), .A2(new_n311_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n310_), .A2(new_n312_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n320_), .A2(new_n734_), .A3(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT119), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT119), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n320_), .A2(new_n734_), .A3(new_n738_), .A4(new_n735_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n733_), .A2(new_n737_), .A3(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT120), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n733_), .A2(new_n737_), .A3(KEYINPUT120), .A4(new_n739_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n284_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n262_), .B1(new_n270_), .B2(new_n273_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n746_), .A2(KEYINPUT116), .A3(new_n276_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT116), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n268_), .A2(KEYINPUT69), .A3(new_n269_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n272_), .B1(new_n271_), .B2(KEYINPUT12), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n261_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n748_), .B1(new_n751_), .B2(new_n204_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n747_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT117), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT55), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT115), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n274_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n274_), .A2(new_n756_), .A3(new_n755_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n753_), .A2(new_n754_), .A3(new_n758_), .A4(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n759_), .A2(new_n752_), .A3(new_n747_), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT117), .B1(new_n761_), .B2(new_n757_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n282_), .B1(new_n760_), .B2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT56), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n745_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n759_), .A2(new_n752_), .A3(new_n747_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n754_), .B1(new_n766_), .B2(new_n758_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n761_), .A2(KEYINPUT117), .A3(new_n757_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n281_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT56), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT121), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n765_), .A2(new_n770_), .A3(new_n771_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n772_), .A2(KEYINPUT122), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n765_), .A2(new_n770_), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT121), .B1(KEYINPUT122), .B2(KEYINPUT58), .ZN(new_n775_));
  OAI22_X1  g574(.A1(new_n773_), .A2(KEYINPUT58), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n744_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n284_), .A2(new_n322_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n760_), .A2(new_n762_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT118), .B1(new_n780_), .B2(new_n281_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n779_), .B1(new_n781_), .B2(KEYINPUT56), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n764_), .B1(new_n763_), .B2(KEYINPUT118), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n778_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(KEYINPUT57), .B1(new_n784_), .B2(new_n349_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT118), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n769_), .A2(new_n786_), .A3(KEYINPUT56), .ZN(new_n787_));
  INV_X1    g586(.A(new_n779_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n783_), .A3(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n777_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT57), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n791_), .A3(new_n348_), .ZN(new_n792_));
  AOI22_X1  g591(.A1(new_n776_), .A2(new_n569_), .B1(new_n785_), .B2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n732_), .B1(new_n793_), .B2(new_n676_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n597_), .A2(new_n535_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n796_), .A2(new_n562_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n794_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT59), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT58), .B1(new_n772_), .B2(KEYINPUT122), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n775_), .B1(new_n765_), .B2(new_n770_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n569_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n791_), .B1(new_n790_), .B2(new_n348_), .ZN(new_n804_));
  AOI211_X1 g603(.A(KEYINPUT57), .B(new_n349_), .C1(new_n789_), .C2(new_n777_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n803_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n731_), .B1(new_n806_), .B2(new_n556_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n797_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT59), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n728_), .B1(new_n800_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n732_), .B1(new_n793_), .B2(new_n557_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n812_), .A2(new_n322_), .A3(new_n797_), .ZN(new_n813_));
  INV_X1    g612(.A(G113gat), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n813_), .A2(KEYINPUT123), .A3(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT123), .B1(new_n813_), .B2(new_n814_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n811_), .A2(new_n815_), .A3(new_n816_), .ZN(G1340gat));
  INV_X1    g616(.A(KEYINPUT60), .ZN(new_n818_));
  INV_X1    g617(.A(G120gat), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n295_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n820_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n809_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n567_), .B1(new_n800_), .B2(new_n810_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n823_), .B2(new_n819_), .ZN(G1341gat));
  NAND2_X1  g623(.A1(new_n557_), .A2(G127gat), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n825_), .B1(new_n800_), .B2(new_n810_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n812_), .A2(new_n676_), .A3(new_n797_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT124), .ZN(new_n828_));
  INV_X1    g627(.A(G127gat), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n827_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n828_), .B1(new_n827_), .B2(new_n829_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n826_), .A2(new_n830_), .A3(new_n831_), .ZN(G1342gat));
  INV_X1    g631(.A(G134gat), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n809_), .A2(new_n833_), .A3(new_n349_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n569_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(new_n800_), .B2(new_n810_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n834_), .B1(new_n836_), .B2(new_n833_), .ZN(G1343gat));
  NAND2_X1  g636(.A1(new_n806_), .A2(new_n556_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n539_), .B1(new_n838_), .B2(new_n732_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT125), .B1(new_n839_), .B2(new_n795_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT125), .ZN(new_n841_));
  NOR4_X1   g640(.A1(new_n807_), .A2(new_n841_), .A3(new_n539_), .A4(new_n796_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n322_), .B1(new_n840_), .B2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(G141gat), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n785_), .A2(new_n792_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n557_), .B1(new_n845_), .B2(new_n803_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n540_), .B(new_n795_), .C1(new_n846_), .C2(new_n731_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n841_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n812_), .A2(KEYINPUT125), .A3(new_n540_), .A4(new_n795_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n850_), .A2(new_n435_), .A3(new_n322_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n844_), .A2(new_n851_), .ZN(G1344gat));
  OAI21_X1  g651(.A(new_n295_), .B1(new_n840_), .B2(new_n842_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(G148gat), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n850_), .A2(new_n436_), .A3(new_n295_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(G1345gat));
  XNOR2_X1  g655(.A(KEYINPUT61), .B(G155gat), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(new_n850_), .B2(new_n676_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n857_), .ZN(new_n859_));
  AOI211_X1 g658(.A(new_n570_), .B(new_n859_), .C1(new_n848_), .C2(new_n849_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n858_), .A2(new_n860_), .ZN(G1346gat));
  NAND3_X1  g660(.A1(new_n850_), .A2(new_n442_), .A3(new_n349_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n835_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n442_), .B2(new_n863_), .ZN(G1347gat));
  NOR2_X1   g663(.A1(new_n534_), .A2(new_n632_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n390_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(KEYINPUT126), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(new_n621_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n794_), .A2(new_n322_), .A3(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT62), .ZN(new_n870_));
  AND3_X1   g669(.A1(new_n869_), .A2(new_n870_), .A3(G169gat), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n869_), .B2(G169gat), .ZN(new_n872_));
  INV_X1    g671(.A(new_n368_), .ZN(new_n873_));
  OAI22_X1  g672(.A1(new_n871_), .A2(new_n872_), .B1(new_n873_), .B2(new_n869_), .ZN(G1348gat));
  NAND2_X1  g673(.A1(new_n794_), .A2(new_n868_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(G176gat), .B1(new_n876_), .B2(new_n295_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n807_), .A2(new_n621_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n867_), .A2(new_n365_), .A3(new_n567_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n877_), .B1(new_n878_), .B2(new_n879_), .ZN(G1349gat));
  NOR3_X1   g679(.A1(new_n875_), .A2(new_n556_), .A3(new_n356_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n867_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n878_), .A2(new_n676_), .A3(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n881_), .B1(new_n360_), .B2(new_n883_), .ZN(G1350gat));
  OAI21_X1  g683(.A(G190gat), .B1(new_n875_), .B2(new_n835_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n349_), .A2(new_n358_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n875_), .B2(new_n886_), .ZN(G1351gat));
  NAND2_X1  g686(.A1(new_n839_), .A2(new_n865_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(new_n323_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(new_n402_), .ZN(G1352gat));
  NOR2_X1   g689(.A1(new_n888_), .A2(new_n567_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(new_n403_), .ZN(G1353gat));
  AOI21_X1  g691(.A(new_n556_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n893_));
  XOR2_X1   g692(.A(new_n893_), .B(KEYINPUT127), .Z(new_n894_));
  NOR2_X1   g693(.A1(new_n888_), .A2(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1354gat));
  OAI21_X1  g696(.A(G218gat), .B1(new_n888_), .B2(new_n835_), .ZN(new_n898_));
  OR2_X1    g697(.A1(new_n348_), .A2(G218gat), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n888_), .B2(new_n899_), .ZN(G1355gat));
endmodule


