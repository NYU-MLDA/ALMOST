//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n891_, new_n892_, new_n894_, new_n895_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G113gat), .B(G120gat), .Z(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n206_));
  AND2_X1   g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207_));
  MUX2_X1   g006(.A(KEYINPUT23), .B(new_n206_), .S(new_n207_), .Z(new_n208_));
  OAI21_X1  g007(.A(new_n208_), .B1(G183gat), .B2(G190gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT82), .ZN(new_n211_));
  INV_X1    g010(.A(G176gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT22), .B(G169gat), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n211_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n209_), .A2(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n211_), .A2(new_n216_), .ZN(new_n217_));
  NOR3_X1   g016(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT23), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n207_), .A2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n221_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n222_));
  INV_X1    g021(.A(G183gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT25), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT80), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT26), .B(G190gat), .ZN(new_n226_));
  OR3_X1    g025(.A1(new_n223_), .A2(KEYINPUT81), .A3(KEYINPUT25), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n223_), .A2(KEYINPUT25), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT81), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .A4(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n219_), .A2(new_n222_), .A3(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n215_), .A2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT84), .B(KEYINPUT30), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G227gat), .A2(G233gat), .ZN(new_n236_));
  INV_X1    g035(.A(G15gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(G43gat), .ZN(new_n239_));
  XOR2_X1   g038(.A(G71gat), .B(G99gat), .Z(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n235_), .A2(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(new_n242_), .B(KEYINPUT86), .Z(new_n243_));
  INV_X1    g042(.A(KEYINPUT31), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n235_), .A2(new_n241_), .ZN(new_n245_));
  XOR2_X1   g044(.A(new_n245_), .B(KEYINPUT85), .Z(new_n246_));
  NAND3_X1  g045(.A1(new_n243_), .A2(new_n244_), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n244_), .B1(new_n243_), .B2(new_n246_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n205_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n249_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n251_), .A2(new_n204_), .A3(new_n247_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(G155gat), .B(G162gat), .Z(new_n255_));
  INV_X1    g054(.A(G141gat), .ZN(new_n256_));
  INV_X1    g055(.A(G148gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT3), .ZN(new_n259_));
  OR3_X1    g058(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G141gat), .A2(G148gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT87), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n259_), .B(new_n260_), .C1(KEYINPUT2), .C2(new_n263_), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n263_), .A2(KEYINPUT2), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n255_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT1), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n255_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n268_), .A2(new_n261_), .A3(new_n258_), .A4(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n266_), .A2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n271_), .A2(KEYINPUT29), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT89), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n272_), .B(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G22gat), .B(G50gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(G218gat), .ZN(new_n278_));
  AOI21_X1  g077(.A(KEYINPUT90), .B1(new_n278_), .B2(G211gat), .ZN(new_n279_));
  XOR2_X1   g078(.A(G197gat), .B(G204gat), .Z(new_n280_));
  OAI221_X1 g079(.A(new_n279_), .B1(G211gat), .B2(new_n278_), .C1(new_n280_), .C2(KEYINPUT21), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(KEYINPUT21), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n283_), .B1(KEYINPUT29), .B2(new_n271_), .ZN(new_n284_));
  INV_X1    g083(.A(G78gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(G106gat), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n287_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G228gat), .A2(G233gat), .ZN(new_n290_));
  INV_X1    g089(.A(new_n283_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n290_), .B1(new_n291_), .B2(KEYINPUT91), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n288_), .A2(new_n289_), .A3(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n293_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n277_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n288_), .A2(new_n289_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(new_n292_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n277_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n299_), .A2(new_n300_), .A3(new_n294_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n297_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G1gat), .B(G29gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(G85gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT0), .B(G57gat), .ZN(new_n305_));
  XOR2_X1   g104(.A(new_n304_), .B(new_n305_), .Z(new_n306_));
  INV_X1    g105(.A(new_n271_), .ZN(new_n307_));
  NOR3_X1   g106(.A1(new_n307_), .A2(new_n205_), .A3(KEYINPUT4), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n271_), .B(new_n205_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n308_), .B1(new_n309_), .B2(KEYINPUT4), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G225gat), .A2(G233gat), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n311_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n309_), .A2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n306_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT33), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n309_), .A2(KEYINPUT95), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n309_), .A2(KEYINPUT95), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n318_), .A2(new_n319_), .A3(new_n313_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n306_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n315_), .A2(new_n316_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n317_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n229_), .A2(new_n224_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n218_), .B1(new_n325_), .B2(new_n226_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n210_), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n326_), .B(new_n208_), .C1(new_n327_), .C2(new_n216_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n222_), .B1(G183gat), .B2(G190gat), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n329_), .A2(KEYINPUT92), .A3(new_n214_), .ZN(new_n330_));
  AOI21_X1  g129(.A(KEYINPUT92), .B1(new_n329_), .B2(new_n214_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n328_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n332_), .A2(new_n291_), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n333_), .A2(KEYINPUT93), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(KEYINPUT93), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n283_), .A2(new_n215_), .A3(new_n232_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n334_), .A2(KEYINPUT20), .A3(new_n335_), .A4(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G226gat), .A2(G233gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT19), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n283_), .B1(new_n215_), .B2(new_n232_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT20), .ZN(new_n342_));
  NOR3_X1   g141(.A1(new_n341_), .A2(new_n342_), .A3(new_n339_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n343_), .B1(new_n291_), .B2(new_n332_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n340_), .A2(new_n344_), .ZN(new_n345_));
  XOR2_X1   g144(.A(G8gat), .B(G36gat), .Z(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G64gat), .B(G92gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n345_), .A2(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n350_), .B1(new_n340_), .B2(new_n344_), .ZN(new_n353_));
  OR3_X1    g152(.A1(new_n324_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n329_), .A2(new_n214_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n283_), .A2(new_n355_), .A3(new_n328_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT20), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n339_), .B1(new_n357_), .B2(new_n341_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n358_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n350_), .A2(KEYINPUT32), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  OR3_X1    g161(.A1(new_n312_), .A2(new_n306_), .A3(new_n314_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(new_n315_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n362_), .B(new_n364_), .C1(new_n361_), .C2(new_n345_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n302_), .B1(new_n354_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n364_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n302_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT27), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n369_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n359_), .A2(new_n351_), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n371_), .B(KEYINPUT27), .C1(new_n351_), .C2(new_n345_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n368_), .A2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n254_), .B1(new_n366_), .B2(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n373_), .A2(new_n302_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n376_), .A2(new_n367_), .A3(new_n253_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G29gat), .B(G36gat), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n379_), .A2(KEYINPUT73), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n379_), .A2(KEYINPUT73), .ZN(new_n381_));
  XOR2_X1   g180(.A(G43gat), .B(G50gat), .Z(new_n382_));
  OR3_X1    g181(.A1(new_n380_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n382_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT74), .B(KEYINPUT15), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  OR2_X1    g186(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n388_));
  NAND2_X1  g187(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n388_), .A2(G85gat), .A3(G92gat), .A4(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(G85gat), .ZN(new_n391_));
  INV_X1    g190(.A(G92gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G85gat), .A2(G92gat), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n393_), .A2(KEYINPUT65), .A3(KEYINPUT9), .A4(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G99gat), .A2(G106gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT6), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT6), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(G99gat), .A3(G106gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  OR2_X1    g199(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(new_n287_), .A3(new_n402_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n390_), .A2(new_n395_), .A3(new_n400_), .A4(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT7), .ZN(new_n406_));
  INV_X1    g205(.A(G99gat), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(new_n407_), .A3(new_n287_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n400_), .A2(new_n405_), .A3(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT8), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n393_), .A2(new_n394_), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n409_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n410_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n404_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n387_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n404_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n397_), .A2(new_n399_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n408_), .A2(new_n405_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n411_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT8), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n409_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n416_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n422_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G232gat), .A2(G233gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT34), .ZN(new_n425_));
  OR2_X1    g224(.A1(new_n425_), .A2(KEYINPUT35), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n415_), .A2(new_n423_), .A3(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n425_), .A2(KEYINPUT35), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G190gat), .B(G218gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G134gat), .B(G162gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n433_), .A2(KEYINPUT36), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n427_), .A2(KEYINPUT35), .A3(new_n425_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n430_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(new_n433_), .B(KEYINPUT36), .Z(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n438_), .B1(new_n430_), .B2(new_n435_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n436_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n378_), .A2(new_n441_), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n442_), .A2(KEYINPUT98), .ZN(new_n443_));
  XOR2_X1   g242(.A(G127gat), .B(G155gat), .Z(new_n444_));
  XNOR2_X1  g243(.A(G183gat), .B(G211gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT17), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT67), .ZN(new_n450_));
  INV_X1    g249(.A(G64gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(G57gat), .ZN(new_n452_));
  INV_X1    g251(.A(G57gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(G64gat), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(new_n454_), .A3(KEYINPUT11), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT66), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n452_), .A2(new_n454_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT11), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT66), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n452_), .A2(new_n454_), .A3(new_n460_), .A4(KEYINPUT11), .ZN(new_n461_));
  AND2_X1   g260(.A1(G71gat), .A2(G78gat), .ZN(new_n462_));
  NOR2_X1   g261(.A1(G71gat), .A2(G78gat), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n456_), .A2(new_n459_), .A3(new_n461_), .A4(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  AOI22_X1  g265(.A1(new_n456_), .A2(new_n461_), .B1(new_n459_), .B2(new_n464_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n450_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G57gat), .B(G64gat), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n464_), .B1(new_n469_), .B2(KEYINPUT11), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n460_), .B1(new_n469_), .B2(KEYINPUT11), .ZN(new_n471_));
  AND4_X1   g270(.A1(new_n460_), .A2(new_n452_), .A3(new_n454_), .A4(KEYINPUT11), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n470_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(new_n465_), .A3(KEYINPUT67), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n468_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G15gat), .B(G22gat), .ZN(new_n477_));
  INV_X1    g276(.A(G1gat), .ZN(new_n478_));
  INV_X1    g277(.A(G8gat), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT14), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G1gat), .B(G8gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G231gat), .A2(G233gat), .ZN(new_n484_));
  XOR2_X1   g283(.A(new_n484_), .B(KEYINPUT76), .Z(new_n485_));
  XNOR2_X1  g284(.A(new_n483_), .B(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n449_), .B1(new_n476_), .B2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n487_), .B1(new_n476_), .B2(new_n486_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n466_), .A2(new_n467_), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n486_), .B(new_n489_), .Z(new_n490_));
  XOR2_X1   g289(.A(KEYINPUT78), .B(KEYINPUT17), .Z(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n448_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n488_), .A2(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n493_), .B1(new_n442_), .B2(KEYINPUT98), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n473_), .A2(new_n465_), .A3(KEYINPUT12), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT68), .B1(new_n422_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT68), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n414_), .A2(new_n489_), .A3(new_n497_), .A4(KEYINPUT12), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n473_), .A2(new_n465_), .A3(KEYINPUT67), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT67), .B1(new_n473_), .B2(new_n465_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n414_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT12), .ZN(new_n502_));
  AOI22_X1  g301(.A1(new_n496_), .A2(new_n498_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n468_), .A2(new_n422_), .A3(new_n474_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G230gat), .A2(G233gat), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n505_), .B(KEYINPUT64), .Z(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n504_), .A2(KEYINPUT69), .A3(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT69), .B1(new_n504_), .B2(new_n507_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n503_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT70), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n504_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n501_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n506_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n503_), .B(KEYINPUT70), .C1(new_n508_), .C2(new_n509_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n512_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  XOR2_X1   g316(.A(G120gat), .B(G148gat), .Z(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT72), .ZN(new_n519_));
  XOR2_X1   g318(.A(G176gat), .B(G204gat), .Z(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n521_), .B(new_n522_), .Z(new_n523_));
  XNOR2_X1  g322(.A(new_n517_), .B(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT13), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n524_), .A2(new_n525_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n387_), .A2(new_n483_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n385_), .A2(new_n483_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G229gat), .A2(G233gat), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n530_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n385_), .B(new_n483_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n532_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G113gat), .B(G141gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G169gat), .B(G197gat), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n537_), .B(new_n538_), .Z(new_n539_));
  NAND3_X1  g338(.A1(new_n533_), .A2(new_n536_), .A3(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT79), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n539_), .B1(new_n533_), .B2(new_n536_), .ZN(new_n543_));
  OR3_X1    g342(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n542_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n529_), .A2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n443_), .A2(new_n494_), .A3(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(G1gat), .B1(new_n549_), .B2(new_n367_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT99), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT37), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n552_), .A2(KEYINPUT75), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(KEYINPUT75), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n440_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n493_), .ZN(new_n556_));
  OAI211_X1 g355(.A(KEYINPUT75), .B(new_n552_), .C1(new_n436_), .C2(new_n439_), .ZN(new_n557_));
  AND3_X1   g356(.A1(new_n555_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n528_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n302_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n365_), .ZN(new_n561_));
  NOR3_X1   g360(.A1(new_n324_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n560_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n302_), .A2(new_n370_), .A3(new_n367_), .A4(new_n372_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n253_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n204_), .B1(new_n251_), .B2(new_n247_), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n248_), .A2(new_n205_), .A3(new_n249_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n367_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n560_), .A2(new_n370_), .A3(new_n372_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n546_), .B1(new_n565_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT96), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  OAI211_X1 g372(.A(KEYINPUT96), .B(new_n546_), .C1(new_n565_), .C2(new_n570_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n559_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n575_), .A2(KEYINPUT97), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(KEYINPUT97), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n578_), .A2(G1gat), .A3(new_n367_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT38), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NOR4_X1   g380(.A1(new_n578_), .A2(KEYINPUT38), .A3(G1gat), .A4(new_n367_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n551_), .B1(new_n581_), .B2(new_n582_), .ZN(G1324gat));
  XNOR2_X1  g382(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n443_), .A2(new_n494_), .A3(new_n548_), .A4(new_n373_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(G8gat), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT39), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT39), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n585_), .A2(new_n588_), .A3(G8gat), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n576_), .A2(new_n479_), .A3(new_n373_), .A4(new_n577_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n584_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n585_), .A2(new_n588_), .A3(G8gat), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n588_), .B1(new_n585_), .B2(G8gat), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n591_), .B(new_n584_), .C1(new_n593_), .C2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n592_), .A2(new_n596_), .ZN(G1325gat));
  OAI21_X1  g396(.A(G15gat), .B1(new_n549_), .B2(new_n254_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT101), .B(KEYINPUT41), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n599_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n253_), .A2(new_n237_), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n600_), .B(new_n601_), .C1(new_n578_), .C2(new_n602_), .ZN(G1326gat));
  OAI21_X1  g402(.A(G22gat), .B1(new_n549_), .B2(new_n560_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n604_), .A2(KEYINPUT42), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(KEYINPUT42), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n560_), .A2(G22gat), .ZN(new_n607_));
  OAI22_X1  g406(.A1(new_n605_), .A2(new_n606_), .B1(new_n578_), .B2(new_n607_), .ZN(G1327gat));
  NAND2_X1  g407(.A1(new_n555_), .A2(new_n557_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n378_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT43), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n378_), .A2(KEYINPUT43), .A3(new_n609_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n612_), .A2(new_n548_), .A3(new_n493_), .A4(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT44), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n556_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n617_), .A2(KEYINPUT44), .A3(new_n548_), .A4(new_n613_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n616_), .A2(new_n364_), .A3(new_n618_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n619_), .A2(KEYINPUT102), .ZN(new_n620_));
  OAI21_X1  g419(.A(G29gat), .B1(new_n619_), .B2(KEYINPUT102), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n441_), .A2(new_n556_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n528_), .A2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n623_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT103), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  AOI211_X1 g425(.A(KEYINPUT103), .B(new_n623_), .C1(new_n573_), .C2(new_n574_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n367_), .A2(G29gat), .ZN(new_n630_));
  OAI22_X1  g429(.A1(new_n620_), .A2(new_n621_), .B1(new_n629_), .B2(new_n630_), .ZN(G1328gat));
  NAND3_X1  g430(.A1(new_n616_), .A2(new_n373_), .A3(new_n618_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(G36gat), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT45), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n373_), .A2(KEYINPUT104), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n373_), .A2(KEYINPUT104), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n637_), .A2(G36gat), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n634_), .B1(new_n628_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n638_), .ZN(new_n640_));
  NOR4_X1   g439(.A1(new_n626_), .A2(new_n627_), .A3(KEYINPUT45), .A4(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n633_), .B1(new_n639_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT46), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  OAI211_X1 g443(.A(new_n633_), .B(KEYINPUT46), .C1(new_n639_), .C2(new_n641_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(G1329gat));
  NAND3_X1  g445(.A1(new_n616_), .A2(new_n253_), .A3(new_n618_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(G43gat), .ZN(new_n648_));
  INV_X1    g447(.A(G43gat), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n628_), .A2(new_n649_), .A3(new_n253_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT47), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n648_), .A2(KEYINPUT47), .A3(new_n650_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1330gat));
  NAND3_X1  g454(.A1(new_n616_), .A2(new_n302_), .A3(new_n618_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n656_), .A2(KEYINPUT105), .ZN(new_n657_));
  OAI21_X1  g456(.A(G50gat), .B1(new_n656_), .B2(KEYINPUT105), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n560_), .A2(G50gat), .ZN(new_n659_));
  OAI22_X1  g458(.A1(new_n657_), .A2(new_n658_), .B1(new_n629_), .B2(new_n659_), .ZN(G1331gat));
  NOR2_X1   g459(.A1(new_n528_), .A2(new_n546_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n378_), .A2(new_n558_), .A3(new_n661_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT106), .Z(new_n663_));
  NAND3_X1  g462(.A1(new_n663_), .A2(new_n453_), .A3(new_n364_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n443_), .A2(new_n494_), .A3(new_n661_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G57gat), .B1(new_n665_), .B2(new_n367_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(G1332gat));
  INV_X1    g466(.A(new_n637_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n663_), .A2(new_n451_), .A3(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(G64gat), .B1(new_n665_), .B2(new_n637_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n670_), .A2(KEYINPUT48), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n670_), .A2(KEYINPUT48), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n669_), .B1(new_n671_), .B2(new_n672_), .ZN(G1333gat));
  INV_X1    g472(.A(G71gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n663_), .A2(new_n674_), .A3(new_n253_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n443_), .A2(new_n494_), .A3(new_n253_), .A4(new_n661_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT49), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n676_), .A2(new_n677_), .A3(G71gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n677_), .B1(new_n676_), .B2(G71gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n675_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT107), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(G1334gat));
  NAND3_X1  g481(.A1(new_n663_), .A2(new_n285_), .A3(new_n302_), .ZN(new_n683_));
  OAI21_X1  g482(.A(G78gat), .B1(new_n665_), .B2(new_n560_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n684_), .A2(KEYINPUT50), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n684_), .A2(KEYINPUT50), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n683_), .B1(new_n685_), .B2(new_n686_), .ZN(G1335gat));
  AND2_X1   g486(.A1(new_n617_), .A2(new_n613_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n688_), .A2(G85gat), .A3(new_n364_), .A4(new_n661_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n378_), .A2(new_n622_), .A3(new_n661_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT108), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n690_), .B(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(new_n364_), .ZN(new_n693_));
  AOI21_X1  g492(.A(KEYINPUT109), .B1(new_n693_), .B2(new_n391_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT109), .ZN(new_n695_));
  AOI211_X1 g494(.A(new_n695_), .B(G85gat), .C1(new_n692_), .C2(new_n364_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n689_), .B1(new_n694_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT110), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n689_), .B(KEYINPUT110), .C1(new_n694_), .C2(new_n696_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1336gat));
  NAND2_X1  g500(.A1(new_n688_), .A2(new_n661_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n702_), .A2(new_n392_), .A3(new_n637_), .ZN(new_n703_));
  AOI21_X1  g502(.A(G92gat), .B1(new_n692_), .B2(new_n373_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT111), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n705_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n703_), .B1(new_n706_), .B2(new_n707_), .ZN(G1337gat));
  OAI21_X1  g507(.A(G99gat), .B1(new_n702_), .B2(new_n254_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n401_), .A2(new_n402_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n692_), .A2(new_n710_), .A3(new_n253_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT112), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n711_), .A2(new_n712_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n709_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT51), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT51), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n717_), .B(new_n709_), .C1(new_n713_), .C2(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(G1338gat));
  NAND3_X1  g518(.A1(new_n692_), .A2(new_n287_), .A3(new_n302_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n617_), .A2(new_n302_), .A3(new_n613_), .A4(new_n661_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT52), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n721_), .A2(new_n722_), .A3(G106gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n721_), .B2(G106gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n720_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g525(.A1(new_n376_), .A2(new_n364_), .A3(new_n253_), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n517_), .A2(new_n523_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n546_), .A2(new_n728_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n503_), .B(KEYINPUT55), .C1(new_n508_), .C2(new_n509_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT114), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n504_), .A2(new_n507_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT69), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n504_), .A2(KEYINPUT69), .A3(new_n507_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n737_), .A2(KEYINPUT114), .A3(KEYINPUT55), .A4(new_n503_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n732_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT55), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n512_), .A2(new_n740_), .A3(new_n516_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n503_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n506_), .B1(new_n742_), .B2(new_n513_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n739_), .A2(new_n741_), .A3(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n744_), .A2(KEYINPUT56), .A3(new_n523_), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT56), .B1(new_n744_), .B2(new_n523_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n746_), .B2(KEYINPUT115), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT115), .ZN(new_n748_));
  AOI211_X1 g547(.A(new_n748_), .B(KEYINPUT56), .C1(new_n744_), .C2(new_n523_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n729_), .B1(new_n747_), .B2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n530_), .A2(new_n531_), .A3(new_n535_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n539_), .B1(new_n534_), .B2(new_n532_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n541_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n524_), .A2(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n440_), .B1(new_n750_), .B2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n744_), .A2(new_n523_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT56), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(KEYINPUT116), .A3(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n728_), .A2(new_n753_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT116), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n745_), .A2(new_n761_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n758_), .B(new_n760_), .C1(new_n762_), .C2(new_n746_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT58), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n609_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n756_), .A2(new_n757_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n766_), .A2(new_n761_), .A3(new_n745_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n759_), .B1(new_n746_), .B2(KEYINPUT116), .ZN(new_n768_));
  AOI21_X1  g567(.A(KEYINPUT58), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  OAI22_X1  g568(.A1(new_n755_), .A2(KEYINPUT57), .B1(new_n765_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT57), .ZN(new_n771_));
  AOI211_X1 g570(.A(new_n771_), .B(new_n440_), .C1(new_n750_), .C2(new_n754_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n493_), .B1(new_n770_), .B2(new_n772_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n774_), .B1(new_n559_), .B2(new_n546_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(KEYINPUT113), .A2(KEYINPUT54), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n558_), .A2(new_n547_), .A3(new_n528_), .A4(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n727_), .B1(new_n773_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT59), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT117), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n775_), .A2(new_n777_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n766_), .A2(new_n748_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n746_), .A2(KEYINPUT115), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n784_), .A2(new_n785_), .A3(new_n745_), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n786_), .A2(new_n729_), .B1(new_n524_), .B2(new_n753_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n771_), .B1(new_n787_), .B2(new_n440_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n763_), .A2(new_n764_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n767_), .A2(new_n768_), .A3(KEYINPUT58), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n609_), .A3(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n755_), .A2(KEYINPUT57), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n788_), .A2(new_n791_), .A3(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n783_), .B1(new_n793_), .B2(new_n493_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n782_), .B(KEYINPUT59), .C1(new_n794_), .C2(new_n727_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT118), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n750_), .A2(new_n754_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT57), .B1(new_n797_), .B2(new_n441_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n765_), .A2(new_n769_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n796_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n791_), .B(KEYINPUT118), .C1(new_n755_), .C2(KEYINPUT57), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n800_), .A2(new_n792_), .A3(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n493_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n778_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n727_), .A2(KEYINPUT59), .ZN(new_n805_));
  AOI22_X1  g604(.A1(new_n781_), .A2(new_n795_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n546_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(G113gat), .ZN(new_n808_));
  INV_X1    g607(.A(new_n779_), .ZN(new_n809_));
  OR2_X1    g608(.A1(new_n547_), .A2(G113gat), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n808_), .B1(new_n809_), .B2(new_n810_), .ZN(G1340gat));
  INV_X1    g610(.A(KEYINPUT121), .ZN(new_n812_));
  XOR2_X1   g611(.A(KEYINPUT119), .B(G120gat), .Z(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(new_n806_), .B2(new_n529_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT120), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n528_), .A2(KEYINPUT60), .ZN(new_n816_));
  MUX2_X1   g615(.A(KEYINPUT60), .B(new_n816_), .S(new_n813_), .Z(new_n817_));
  AND3_X1   g616(.A1(new_n779_), .A2(new_n815_), .A3(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n815_), .B1(new_n779_), .B2(new_n817_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n812_), .B1(new_n814_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n781_), .A2(new_n795_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n804_), .A2(new_n805_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n822_), .A2(new_n529_), .A3(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n813_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n820_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(KEYINPUT121), .A3(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n821_), .A2(new_n828_), .ZN(G1341gat));
  NAND2_X1  g628(.A1(new_n806_), .A2(new_n556_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(G127gat), .ZN(new_n831_));
  OR2_X1    g630(.A1(new_n493_), .A2(G127gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n809_), .B2(new_n832_), .ZN(G1342gat));
  NAND2_X1  g632(.A1(new_n806_), .A2(new_n609_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(G134gat), .ZN(new_n835_));
  OR2_X1    g634(.A1(new_n441_), .A2(G134gat), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n809_), .B2(new_n836_), .ZN(G1343gat));
  NOR2_X1   g636(.A1(new_n794_), .A2(new_n253_), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n668_), .A2(new_n367_), .A3(new_n560_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n840_), .A2(new_n547_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(new_n256_), .ZN(G1344gat));
  NOR2_X1   g641(.A1(new_n840_), .A2(new_n528_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(new_n257_), .ZN(G1345gat));
  OAI21_X1  g643(.A(KEYINPUT122), .B1(new_n840_), .B2(new_n493_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n838_), .A2(new_n846_), .A3(new_n556_), .A4(new_n839_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT61), .B(G155gat), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n848_), .B(new_n850_), .ZN(G1346gat));
  INV_X1    g650(.A(new_n609_), .ZN(new_n852_));
  OAI21_X1  g651(.A(G162gat), .B1(new_n840_), .B2(new_n852_), .ZN(new_n853_));
  OR2_X1    g652(.A1(new_n441_), .A2(G162gat), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n840_), .B2(new_n854_), .ZN(G1347gat));
  NOR2_X1   g654(.A1(new_n637_), .A2(new_n568_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n560_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(new_n803_), .B2(new_n778_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n858_), .A2(new_n546_), .A3(new_n213_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n857_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n772_), .B1(new_n770_), .B2(new_n796_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n556_), .B1(new_n861_), .B2(new_n801_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n546_), .B(new_n860_), .C1(new_n862_), .C2(new_n783_), .ZN(new_n863_));
  XOR2_X1   g662(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n864_));
  NAND3_X1  g663(.A1(new_n863_), .A2(G169gat), .A3(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT124), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n863_), .A2(KEYINPUT124), .A3(G169gat), .A4(new_n864_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT125), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n864_), .B1(new_n863_), .B2(G169gat), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n867_), .B(new_n868_), .C1(new_n869_), .C2(new_n870_), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n870_), .A2(new_n869_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n859_), .B1(new_n871_), .B2(new_n872_), .ZN(G1348gat));
  NOR2_X1   g672(.A1(new_n794_), .A2(new_n302_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n874_), .A2(G176gat), .A3(new_n529_), .A4(new_n856_), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n529_), .B(new_n860_), .C1(new_n862_), .C2(new_n783_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT126), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n876_), .A2(new_n877_), .A3(new_n212_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n876_), .B2(new_n212_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n875_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(KEYINPUT127), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT127), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n882_), .B(new_n875_), .C1(new_n878_), .C2(new_n879_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n883_), .ZN(G1349gat));
  NAND2_X1  g683(.A1(new_n856_), .A2(new_n556_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(G183gat), .B1(new_n874_), .B2(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n493_), .A2(new_n325_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n858_), .B2(new_n888_), .ZN(G1350gat));
  NAND2_X1  g688(.A1(new_n858_), .A2(new_n609_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(G190gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n858_), .A2(new_n226_), .A3(new_n440_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1351gat));
  NOR4_X1   g692(.A1(new_n794_), .A2(new_n368_), .A3(new_n253_), .A4(new_n637_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n546_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n529_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g697(.A1(new_n894_), .A2(new_n556_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n900_));
  AND2_X1   g699(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n899_), .A2(new_n900_), .A3(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n902_), .B1(new_n899_), .B2(new_n900_), .ZN(G1354gat));
  NAND3_X1  g702(.A1(new_n894_), .A2(new_n278_), .A3(new_n440_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n894_), .A2(new_n609_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n905_), .B2(new_n278_), .ZN(G1355gat));
endmodule


