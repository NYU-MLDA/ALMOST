//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 1 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 1 1 1 1 1 1 0 1 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n813_, new_n815_, new_n816_, new_n818_,
    new_n819_, new_n820_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n841_, new_n842_, new_n843_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT65), .B(G85gat), .Z(new_n203_));
  INV_X1    g002(.A(G92gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(KEYINPUT9), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G85gat), .A2(G92gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  AOI22_X1  g008(.A1(new_n203_), .A2(new_n205_), .B1(new_n209_), .B2(KEYINPUT9), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT10), .B(G99gat), .ZN(new_n211_));
  OR3_X1    g010(.A1(new_n211_), .A2(KEYINPUT64), .A3(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G99gat), .A2(G106gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n216_), .A2(KEYINPUT66), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n213_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(KEYINPUT66), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n220_));
  AND2_X1   g019(.A1(G99gat), .A2(G106gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n218_), .A2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT64), .B1(new_n211_), .B2(G106gat), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n210_), .A2(new_n212_), .A3(new_n223_), .A4(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G57gat), .B(G64gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT11), .ZN(new_n227_));
  XOR2_X1   g026(.A(G71gat), .B(G78gat), .Z(new_n228_));
  OR2_X1    g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n226_), .A2(KEYINPUT11), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n227_), .A2(new_n228_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n229_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT7), .ZN(new_n233_));
  INV_X1    g032(.A(G99gat), .ZN(new_n234_));
  INV_X1    g033(.A(G106gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n238_), .B1(new_n218_), .B2(new_n222_), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT67), .B1(new_n207_), .B2(new_n208_), .ZN(new_n240_));
  INV_X1    g039(.A(G85gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(new_n204_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n242_), .A2(new_n243_), .A3(new_n206_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n240_), .A2(new_n244_), .ZN(new_n245_));
  NOR3_X1   g044(.A1(new_n239_), .A2(KEYINPUT8), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT8), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n236_), .A2(new_n237_), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n221_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n248_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n240_), .A2(new_n244_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n247_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n225_), .B(new_n232_), .C1(new_n246_), .C2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(KEYINPUT8), .B1(new_n239_), .B2(new_n245_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n251_), .A2(new_n247_), .A3(new_n252_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n232_), .B1(new_n258_), .B2(new_n225_), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT12), .B1(new_n255_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G230gat), .A2(G233gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT12), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n210_), .A2(new_n223_), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n212_), .A2(new_n224_), .ZN(new_n264_));
  AOI22_X1  g063(.A1(new_n263_), .A2(new_n264_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n262_), .B1(new_n265_), .B2(new_n232_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n260_), .A2(new_n261_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT68), .ZN(new_n268_));
  OAI211_X1 g067(.A(G230gat), .B(G233gat), .C1(new_n255_), .C2(new_n259_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n260_), .A2(new_n270_), .A3(new_n261_), .A4(new_n266_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n268_), .A2(new_n269_), .A3(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT69), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n268_), .A2(new_n274_), .A3(new_n269_), .A4(new_n271_), .ZN(new_n275_));
  XOR2_X1   g074(.A(G120gat), .B(G148gat), .Z(new_n276_));
  XNOR2_X1  g075(.A(G176gat), .B(G204gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n279_));
  XOR2_X1   g078(.A(new_n278_), .B(new_n279_), .Z(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  AND4_X1   g080(.A1(new_n202_), .A2(new_n273_), .A3(new_n275_), .A4(new_n281_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n268_), .A2(new_n269_), .A3(new_n271_), .A4(new_n280_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT71), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n280_), .B1(new_n272_), .B2(KEYINPUT69), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n284_), .B1(new_n285_), .B2(new_n275_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT72), .B1(new_n282_), .B2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n273_), .A2(new_n275_), .A3(new_n281_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n284_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n285_), .A2(new_n202_), .A3(new_n275_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  AND3_X1   g092(.A1(new_n287_), .A2(KEYINPUT13), .A3(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT13), .B1(new_n287_), .B2(new_n293_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT77), .B(G1gat), .ZN(new_n297_));
  INV_X1    g096(.A(G8gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT14), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G15gat), .B(G22gat), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G1gat), .B(G8gat), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n302_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(G29gat), .B(G36gat), .Z(new_n306_));
  XOR2_X1   g105(.A(G43gat), .B(G50gat), .Z(new_n307_));
  XOR2_X1   g106(.A(new_n306_), .B(new_n307_), .Z(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n305_), .B(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G229gat), .A2(G233gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n308_), .B(KEYINPUT15), .Z(new_n313_));
  INV_X1    g112(.A(new_n305_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n312_), .B1(new_n305_), .B2(new_n309_), .ZN(new_n316_));
  AOI22_X1  g115(.A1(new_n310_), .A2(new_n312_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G113gat), .B(G141gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT80), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G169gat), .B(G197gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n317_), .B(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n296_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT25), .B(G183gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT26), .B(G190gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(G169gat), .ZN(new_n328_));
  INV_X1    g127(.A(G176gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G169gat), .A2(G176gat), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n330_), .A2(KEYINPUT24), .A3(new_n331_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n327_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT81), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G183gat), .A2(G190gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT23), .ZN(new_n336_));
  OR2_X1    g135(.A1(new_n330_), .A2(KEYINPUT24), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n327_), .A2(new_n332_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT81), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n334_), .A2(new_n338_), .A3(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(new_n328_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  OR2_X1    g144(.A1(G183gat), .A2(G190gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n336_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n342_), .A2(KEYINPUT30), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(KEYINPUT30), .B1(new_n342_), .B2(new_n348_), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT83), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n342_), .A2(new_n348_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT30), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT83), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n342_), .A2(KEYINPUT30), .A3(new_n348_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G71gat), .B(G99gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(G43gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT82), .B(G15gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G227gat), .A2(G233gat), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n361_), .B(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n351_), .A2(new_n357_), .A3(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n361_), .B(new_n362_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n366_), .A2(new_n355_), .A3(new_n354_), .A4(new_n356_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT85), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT85), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n365_), .A2(new_n370_), .A3(new_n367_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G127gat), .B(G134gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G113gat), .B(G120gat), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT84), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n372_), .A2(new_n373_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n372_), .A2(new_n373_), .A3(KEYINPUT84), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT31), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n369_), .A2(new_n371_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n380_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n368_), .A2(KEYINPUT85), .A3(new_n382_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n381_), .A2(KEYINPUT86), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(KEYINPUT86), .B1(new_n381_), .B2(new_n383_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G78gat), .B(G106gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT95), .ZN(new_n388_));
  INV_X1    g187(.A(G141gat), .ZN(new_n389_));
  INV_X1    g188(.A(G148gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G141gat), .A2(G148gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G155gat), .A2(G162gat), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT87), .B1(new_n393_), .B2(KEYINPUT1), .ZN(new_n394_));
  OR2_X1    g193(.A1(G155gat), .A2(G162gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(KEYINPUT1), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  NOR3_X1   g196(.A1(new_n393_), .A2(KEYINPUT87), .A3(KEYINPUT1), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n391_), .B(new_n392_), .C1(new_n397_), .C2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT2), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n392_), .A2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT3), .ZN(new_n403_));
  NOR2_X1   g202(.A1(G141gat), .A2(G148gat), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n401_), .B(new_n402_), .C1(new_n403_), .C2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT88), .ZN(new_n406_));
  AOI21_X1  g205(.A(KEYINPUT3), .B1(new_n391_), .B2(new_n406_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n407_), .B(KEYINPUT89), .C1(new_n406_), .C2(new_n391_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT89), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n391_), .A2(new_n406_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n403_), .B1(new_n404_), .B2(KEYINPUT88), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n409_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n405_), .B1(new_n408_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n395_), .A2(new_n393_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n399_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT29), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G197gat), .B(G204gat), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT21), .ZN(new_n418_));
  OR2_X1    g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G211gat), .B(G218gat), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n417_), .A2(new_n418_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT94), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n417_), .A2(KEYINPUT94), .A3(new_n418_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n424_), .A2(new_n419_), .A3(new_n425_), .A4(new_n420_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n421_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(G233gat), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n428_), .A2(KEYINPUT92), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(KEYINPUT92), .ZN(new_n430_));
  OAI21_X1  g229(.A(G228gat), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT93), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT91), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n416_), .A2(new_n427_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n431_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n415_), .A2(KEYINPUT91), .A3(KEYINPUT29), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n421_), .A2(new_n426_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n438_), .A2(new_n432_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n436_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n388_), .B1(new_n435_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT96), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT29), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n443_), .B(new_n399_), .C1(new_n413_), .C2(new_n414_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G22gat), .B(G50gat), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  XOR2_X1   g245(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n447_));
  NAND2_X1  g246(.A1(new_n444_), .A2(new_n445_), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n446_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n447_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n442_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n388_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n437_), .A2(new_n439_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n453_), .B(new_n434_), .C1(new_n454_), .C2(new_n436_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n441_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n452_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT96), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n451_), .A2(new_n455_), .A3(new_n458_), .A4(new_n441_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G225gat), .A2(G233gat), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n413_), .A2(new_n414_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT101), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n374_), .A2(new_n376_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n463_), .A2(new_n464_), .A3(new_n399_), .A4(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n415_), .A2(new_n379_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n465_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT101), .B1(new_n415_), .B2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n466_), .A2(new_n467_), .A3(new_n469_), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n470_), .A2(KEYINPUT4), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT4), .B1(new_n415_), .B2(new_n379_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n462_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G1gat), .B(G29gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(G85gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT0), .B(G57gat), .ZN(new_n476_));
  XOR2_X1   g275(.A(new_n475_), .B(new_n476_), .Z(new_n477_));
  AND3_X1   g276(.A1(new_n466_), .A2(new_n467_), .A3(new_n469_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n461_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n473_), .A2(KEYINPUT33), .A3(new_n477_), .A4(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n472_), .B1(new_n470_), .B2(KEYINPUT4), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n479_), .B(new_n477_), .C1(new_n481_), .C2(new_n461_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT33), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT99), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n344_), .B1(new_n347_), .B2(KEYINPUT98), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT98), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n336_), .A2(new_n487_), .A3(new_n346_), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n486_), .A2(new_n488_), .B1(new_n333_), .B2(new_n338_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n485_), .B1(new_n438_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n347_), .A2(KEYINPUT98), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n491_), .A2(new_n345_), .A3(new_n488_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n333_), .A2(new_n338_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n494_), .A2(KEYINPUT99), .A3(new_n427_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n438_), .A2(new_n342_), .A3(new_n348_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n490_), .A2(new_n495_), .A3(new_n496_), .A4(KEYINPUT20), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G226gat), .A2(G233gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n438_), .B1(new_n348_), .B2(new_n342_), .ZN(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT20), .B1(new_n494_), .B2(new_n427_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n500_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  XOR2_X1   g305(.A(G8gat), .B(G36gat), .Z(new_n507_));
  XNOR2_X1  g306(.A(G64gat), .B(G92gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(KEYINPUT100), .B(KEYINPUT18), .Z(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  AND3_X1   g310(.A1(new_n501_), .A2(new_n506_), .A3(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n511_), .B1(new_n501_), .B2(new_n506_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n477_), .B1(new_n478_), .B2(new_n462_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n515_), .B1(new_n462_), .B2(new_n481_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n480_), .A2(new_n484_), .A3(new_n514_), .A4(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n479_), .B1(new_n481_), .B2(new_n461_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n477_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(new_n482_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n500_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n522_), .B1(new_n497_), .B2(new_n500_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n511_), .A2(KEYINPUT32), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n524_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n501_), .A2(new_n506_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n525_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n521_), .A2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n460_), .B1(new_n517_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n459_), .ZN(new_n531_));
  AOI22_X1  g330(.A1(new_n442_), .A2(new_n451_), .B1(new_n455_), .B2(new_n441_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT103), .B(KEYINPUT27), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n534_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n511_), .B(KEYINPUT102), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n523_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n501_), .A2(new_n506_), .A3(new_n511_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n537_), .A2(KEYINPUT27), .A3(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n535_), .A2(new_n539_), .ZN(new_n540_));
  NOR3_X1   g339(.A1(new_n533_), .A2(new_n540_), .A3(new_n521_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n386_), .B1(new_n530_), .B2(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n460_), .A2(new_n540_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n521_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n381_), .A2(new_n383_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n542_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n265_), .A2(new_n308_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n548_), .B1(new_n313_), .B2(new_n265_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT73), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G232gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n551_), .A2(new_n554_), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n551_), .B(new_n554_), .C1(KEYINPUT35), .C2(new_n549_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G190gat), .B(G218gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT74), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G134gat), .B(G162gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n561_), .A2(KEYINPUT36), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT75), .Z(new_n563_));
  NAND3_X1  g362(.A1(new_n555_), .A2(new_n556_), .A3(new_n563_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n555_), .A2(new_n556_), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n560_), .B(KEYINPUT36), .Z(new_n566_));
  OAI21_X1  g365(.A(new_n564_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT37), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT76), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n568_), .B1(new_n564_), .B2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n567_), .A2(new_n570_), .ZN(new_n571_));
  OAI221_X1 g370(.A(new_n564_), .B1(new_n569_), .B2(new_n568_), .C1(new_n565_), .C2(new_n566_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  XOR2_X1   g373(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT79), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G127gat), .B(G155gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G183gat), .B(G211gat), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n578_), .B(new_n579_), .Z(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT17), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G231gat), .A2(G233gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n232_), .B(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(new_n305_), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n581_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(KEYINPUT17), .A3(new_n580_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n574_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n324_), .A2(new_n547_), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(new_n521_), .A3(new_n297_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(KEYINPUT105), .A2(KEYINPUT38), .ZN(new_n592_));
  AND2_X1   g391(.A1(KEYINPUT105), .A2(KEYINPUT38), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n591_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n594_), .B1(new_n592_), .B2(new_n591_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n567_), .ZN(new_n596_));
  AOI211_X1 g395(.A(new_n596_), .B(new_n587_), .C1(new_n542_), .C2(new_n546_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n324_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT104), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(new_n521_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n595_), .B1(G1gat), .B2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT106), .ZN(G1324gat));
  INV_X1    g401(.A(new_n540_), .ZN(new_n603_));
  OAI21_X1  g402(.A(G8gat), .B1(new_n598_), .B2(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT39), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n590_), .A2(new_n298_), .A3(new_n540_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n607_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g407(.A(G15gat), .ZN(new_n609_));
  INV_X1    g408(.A(new_n386_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n609_), .B1(new_n599_), .B2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT41), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT107), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n613_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n589_), .A2(G15gat), .A3(new_n386_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT108), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n614_), .A2(new_n615_), .A3(new_n617_), .ZN(G1326gat));
  INV_X1    g417(.A(G22gat), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n619_), .B1(new_n599_), .B2(new_n460_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT42), .Z(new_n621_));
  NAND3_X1  g420(.A1(new_n590_), .A2(new_n619_), .A3(new_n460_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(G1327gat));
  INV_X1    g422(.A(new_n587_), .ZN(new_n624_));
  AOI211_X1 g423(.A(new_n567_), .B(new_n624_), .C1(new_n542_), .C2(new_n546_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n324_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(G29gat), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(new_n628_), .A3(new_n521_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT111), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n547_), .A2(new_n574_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(KEYINPUT43), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT43), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n547_), .A2(new_n633_), .A3(new_n574_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n635_), .A2(KEYINPUT44), .A3(new_n324_), .A4(new_n587_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT110), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n633_), .B1(new_n547_), .B2(new_n574_), .ZN(new_n638_));
  AOI211_X1 g437(.A(KEYINPUT43), .B(new_n573_), .C1(new_n542_), .C2(new_n546_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n587_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT110), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n641_), .A2(new_n642_), .A3(KEYINPUT44), .A4(new_n324_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n637_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT44), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n294_), .A2(new_n295_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(new_n322_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n645_), .B1(new_n640_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT109), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  OAI211_X1 g449(.A(KEYINPUT109), .B(new_n645_), .C1(new_n640_), .C2(new_n647_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n644_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(new_n521_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n630_), .B1(new_n653_), .B2(G29gat), .ZN(new_n654_));
  AOI211_X1 g453(.A(KEYINPUT111), .B(new_n628_), .C1(new_n652_), .C2(new_n521_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n629_), .B1(new_n654_), .B2(new_n655_), .ZN(G1328gat));
  NOR3_X1   g455(.A1(new_n626_), .A2(G36gat), .A3(new_n603_), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n657_), .B(KEYINPUT45), .Z(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT112), .B1(new_n652_), .B2(new_n540_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n637_), .A2(new_n643_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n650_), .A2(new_n651_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n660_), .A2(KEYINPUT112), .A3(new_n540_), .A4(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(G36gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n658_), .B1(new_n659_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT46), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  OAI211_X1 g465(.A(KEYINPUT46), .B(new_n658_), .C1(new_n659_), .C2(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1329gat));
  NAND2_X1  g467(.A1(new_n660_), .A2(new_n661_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n545_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G43gat), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  OR3_X1    g470(.A1(new_n626_), .A2(G43gat), .A3(new_n386_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT47), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(G1330gat));
  AOI21_X1  g474(.A(G50gat), .B1(new_n627_), .B2(new_n460_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n460_), .A2(G50gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n652_), .B2(new_n677_), .ZN(G1331gat));
  NAND2_X1  g477(.A1(new_n296_), .A2(new_n588_), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n679_), .A2(KEYINPUT113), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(KEYINPUT113), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n680_), .A2(new_n323_), .A3(new_n547_), .A4(new_n681_), .ZN(new_n682_));
  AOI211_X1 g481(.A(G57gat), .B(new_n544_), .C1(new_n682_), .C2(KEYINPUT114), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n683_), .B1(KEYINPUT114), .B2(new_n682_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n646_), .A2(new_n322_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(new_n597_), .ZN(new_n686_));
  OAI21_X1  g485(.A(G57gat), .B1(new_n686_), .B2(new_n544_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n684_), .A2(new_n687_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT115), .ZN(G1332gat));
  OAI21_X1  g488(.A(G64gat), .B1(new_n686_), .B2(new_n603_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT48), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n603_), .A2(G64gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(new_n682_), .B2(new_n692_), .ZN(G1333gat));
  OAI21_X1  g492(.A(G71gat), .B1(new_n686_), .B2(new_n386_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT49), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n386_), .A2(G71gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n682_), .B2(new_n696_), .ZN(G1334gat));
  OAI21_X1  g496(.A(G78gat), .B1(new_n686_), .B2(new_n533_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT50), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n533_), .A2(G78gat), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n699_), .B1(new_n682_), .B2(new_n700_), .ZN(G1335gat));
  NAND2_X1  g500(.A1(new_n685_), .A2(new_n625_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT116), .Z(new_n703_));
  AOI21_X1  g502(.A(G85gat), .B1(new_n703_), .B2(new_n521_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n640_), .A2(new_n322_), .A3(new_n646_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n521_), .A2(new_n203_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n704_), .B1(new_n705_), .B2(new_n706_), .ZN(G1336gat));
  NAND3_X1  g506(.A1(new_n703_), .A2(new_n204_), .A3(new_n540_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n705_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G92gat), .B1(new_n709_), .B2(new_n603_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(G1337gat));
  AOI21_X1  g510(.A(new_n234_), .B1(new_n705_), .B2(new_n610_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n670_), .A2(new_n211_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n703_), .B2(new_n713_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g514(.A1(new_n703_), .A2(new_n235_), .A3(new_n460_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT117), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n705_), .A2(new_n717_), .A3(new_n460_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n718_), .A2(G106gat), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT52), .ZN(new_n720_));
  OAI21_X1  g519(.A(KEYINPUT117), .B1(new_n709_), .B2(new_n533_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n719_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n720_), .B1(new_n719_), .B2(new_n721_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n716_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT53), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT53), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n726_), .B(new_n716_), .C1(new_n722_), .C2(new_n723_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1339gat));
  INV_X1    g527(.A(KEYINPUT122), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n543_), .A2(new_n521_), .A3(new_n545_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT119), .Z(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n732_), .A2(KEYINPUT59), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n646_), .A2(new_n323_), .A3(new_n588_), .A4(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n735_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n588_), .A2(new_n323_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n737_), .B1(new_n296_), .B2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n736_), .A2(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n321_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n315_), .B(new_n312_), .C1(new_n314_), .C2(new_n308_), .ZN(new_n742_));
  AOI22_X1  g541(.A1(new_n317_), .A2(new_n321_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n743_), .A2(new_n283_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT55), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n268_), .A2(new_n745_), .A3(new_n271_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n260_), .A2(new_n266_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n747_), .A2(G230gat), .A3(G233gat), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n746_), .B(new_n748_), .C1(new_n745_), .C2(new_n267_), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n749_), .A2(KEYINPUT56), .A3(new_n281_), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT56), .B1(new_n749_), .B2(new_n281_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n744_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT58), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  OAI211_X1 g553(.A(KEYINPUT58), .B(new_n744_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n754_), .A2(new_n574_), .A3(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n287_), .A2(new_n293_), .A3(new_n743_), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n322_), .B(new_n283_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n596_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n756_), .B1(new_n759_), .B2(KEYINPUT57), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT120), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT57), .ZN(new_n763_));
  AOI211_X1 g562(.A(new_n763_), .B(new_n596_), .C1(new_n757_), .C2(new_n758_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  OAI211_X1 g564(.A(KEYINPUT120), .B(new_n756_), .C1(new_n759_), .C2(KEYINPUT57), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n762_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(new_n587_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n740_), .B1(new_n768_), .B2(KEYINPUT121), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n764_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n624_), .B1(new_n770_), .B2(new_n766_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT121), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n734_), .B1(new_n769_), .B2(new_n773_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n760_), .A2(new_n764_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n775_), .A2(new_n624_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n776_), .A2(new_n740_), .ZN(new_n777_));
  OAI21_X1  g576(.A(KEYINPUT59), .B1(new_n777_), .B2(new_n732_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n729_), .B1(new_n774_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n773_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n740_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n782_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n733_), .B1(new_n781_), .B2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n784_), .A2(KEYINPUT122), .A3(new_n778_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n780_), .A2(new_n322_), .A3(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(G113gat), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n777_), .A2(new_n732_), .ZN(new_n788_));
  INV_X1    g587(.A(G113gat), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n322_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n787_), .A2(new_n790_), .ZN(G1340gat));
  NOR2_X1   g590(.A1(new_n646_), .A2(KEYINPUT60), .ZN(new_n792_));
  MUX2_X1   g591(.A(new_n792_), .B(KEYINPUT60), .S(G120gat), .Z(new_n793_));
  NAND2_X1  g592(.A1(new_n788_), .A2(new_n793_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n774_), .A2(new_n779_), .A3(new_n646_), .ZN(new_n795_));
  INV_X1    g594(.A(G120gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n794_), .B1(new_n795_), .B2(new_n796_), .ZN(G1341gat));
  NAND3_X1  g596(.A1(new_n780_), .A2(new_n624_), .A3(new_n785_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(G127gat), .ZN(new_n799_));
  INV_X1    g598(.A(G127gat), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n788_), .A2(new_n800_), .A3(new_n624_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(G1342gat));
  NAND3_X1  g601(.A1(new_n780_), .A2(new_n574_), .A3(new_n785_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(G134gat), .ZN(new_n804_));
  INV_X1    g603(.A(G134gat), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n788_), .A2(new_n805_), .A3(new_n596_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(G1343gat));
  NAND4_X1  g606(.A1(new_n386_), .A2(new_n521_), .A3(new_n460_), .A4(new_n603_), .ZN(new_n808_));
  XOR2_X1   g607(.A(new_n808_), .B(KEYINPUT123), .Z(new_n809_));
  NOR2_X1   g608(.A1(new_n777_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n322_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n296_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g613(.A1(new_n810_), .A2(new_n624_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(KEYINPUT61), .B(G155gat), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n815_), .B(new_n816_), .ZN(G1346gat));
  INV_X1    g616(.A(G162gat), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n810_), .A2(new_n818_), .A3(new_n596_), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n777_), .A2(new_n573_), .A3(new_n809_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n819_), .B1(new_n820_), .B2(new_n818_), .ZN(G1347gat));
  NOR2_X1   g620(.A1(new_n603_), .A2(new_n521_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n610_), .A2(new_n533_), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n823_), .B1(new_n769_), .B2(new_n773_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n322_), .ZN(new_n825_));
  XOR2_X1   g624(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n826_));
  INV_X1    g625(.A(KEYINPUT125), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n328_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n825_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n828_), .B1(new_n825_), .B2(new_n829_), .ZN(new_n831_));
  XOR2_X1   g630(.A(KEYINPUT22), .B(G169gat), .Z(new_n832_));
  OAI22_X1  g631(.A1(new_n830_), .A2(new_n831_), .B1(new_n825_), .B2(new_n832_), .ZN(G1348gat));
  AOI21_X1  g632(.A(G176gat), .B1(new_n824_), .B2(new_n296_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n777_), .A2(new_n823_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n646_), .A2(new_n329_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n834_), .B1(new_n835_), .B2(new_n836_), .ZN(G1349gat));
  AOI21_X1  g636(.A(G183gat), .B1(new_n835_), .B2(new_n624_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n587_), .A2(new_n325_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n838_), .B1(new_n824_), .B2(new_n839_), .ZN(G1350gat));
  NAND2_X1  g639(.A1(new_n824_), .A2(new_n574_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(G190gat), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n824_), .A2(new_n326_), .A3(new_n596_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(G1351gat));
  NAND3_X1  g643(.A1(new_n386_), .A2(new_n460_), .A3(new_n822_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n777_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n322_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n296_), .ZN(new_n849_));
  INV_X1    g648(.A(G204gat), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n850_), .A2(KEYINPUT126), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n849_), .B(new_n851_), .ZN(G1353gat));
  NAND2_X1  g651(.A1(new_n846_), .A2(new_n624_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n854_));
  AND2_X1   g653(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n853_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(new_n853_), .B2(new_n854_), .ZN(G1354gat));
  INV_X1    g656(.A(G218gat), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n846_), .A2(new_n858_), .A3(new_n596_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n777_), .A2(new_n573_), .A3(new_n845_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(new_n858_), .ZN(G1355gat));
endmodule


