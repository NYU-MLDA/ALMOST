//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n949_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_,
    new_n959_;
  XOR2_X1   g000(.A(G71gat), .B(G78gat), .Z(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G57gat), .B(G64gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT65), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT11), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n203_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n206_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT65), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n204_), .B(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(KEYINPUT11), .A3(new_n202_), .ZN(new_n211_));
  AND3_X1   g010(.A1(new_n207_), .A2(new_n208_), .A3(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G85gat), .B(G92gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT7), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT6), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n213_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n218_));
  OR3_X1    g017(.A1(new_n218_), .A2(KEYINPUT64), .A3(KEYINPUT8), .ZN(new_n219_));
  INV_X1    g018(.A(new_n213_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT7), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n214_), .B(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT6), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n216_), .B(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n220_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n218_), .A2(KEYINPUT64), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(KEYINPUT8), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n220_), .A2(KEYINPUT9), .ZN(new_n230_));
  XOR2_X1   g029(.A(KEYINPUT10), .B(G99gat), .Z(new_n231_));
  INV_X1    g030(.A(G106gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT9), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n234_), .A2(G85gat), .A3(G92gat), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n230_), .A2(new_n233_), .A3(new_n217_), .A4(new_n235_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n212_), .A2(new_n219_), .A3(new_n229_), .A4(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n229_), .A2(new_n219_), .A3(new_n236_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n207_), .A2(new_n208_), .A3(new_n211_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n237_), .A2(new_n240_), .A3(KEYINPUT12), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT12), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n238_), .A2(new_n242_), .A3(new_n239_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G230gat), .A2(G233gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n237_), .A2(new_n240_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n245_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G176gat), .B(G204gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G120gat), .B(G148gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n254_));
  XOR2_X1   g053(.A(new_n253_), .B(new_n254_), .Z(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT66), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n250_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n246_), .A2(new_n249_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n259_), .A2(KEYINPUT66), .A3(new_n256_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT13), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n258_), .A2(KEYINPUT13), .A3(new_n260_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G29gat), .B(G36gat), .ZN(new_n266_));
  INV_X1    g065(.A(G43gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(G50gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G15gat), .B(G22gat), .ZN(new_n270_));
  INV_X1    g069(.A(G1gat), .ZN(new_n271_));
  INV_X1    g070(.A(G8gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT14), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G1gat), .B(G8gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n269_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(G50gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n268_), .B(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT15), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT15), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n269_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n277_), .B1(new_n283_), .B2(new_n276_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G229gat), .A2(G233gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n269_), .A2(new_n276_), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n287_), .A2(new_n277_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n285_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G113gat), .B(G141gat), .ZN(new_n291_));
  INV_X1    g090(.A(G169gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(G197gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n286_), .A2(new_n290_), .A3(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n296_), .B1(new_n286_), .B2(new_n290_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(new_n299_), .B(KEYINPUT72), .Z(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT25), .B(G183gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT26), .B(G190gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G183gat), .A2(G190gat), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT23), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(G176gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n292_), .A2(new_n309_), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n310_), .A2(KEYINPUT24), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n310_), .A2(KEYINPUT24), .A3(new_n312_), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n303_), .A2(new_n308_), .A3(new_n311_), .A4(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT73), .B(G176gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT22), .B(G169gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  OAI211_X1 g116(.A(new_n306_), .B(new_n307_), .C1(G183gat), .C2(G190gat), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n317_), .A2(new_n318_), .A3(new_n312_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n314_), .A2(new_n319_), .A3(KEYINPUT74), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(KEYINPUT74), .B1(new_n314_), .B2(new_n319_), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT30), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n314_), .A2(new_n319_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT74), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT30), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n326_), .A2(new_n327_), .A3(new_n320_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n323_), .A2(new_n328_), .A3(KEYINPUT75), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G71gat), .B(G99gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G15gat), .B(G43gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G227gat), .A2(G233gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n332_), .B(new_n333_), .Z(new_n334_));
  NAND2_X1  g133(.A1(new_n329_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT31), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT31), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n329_), .A2(new_n337_), .A3(new_n334_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n323_), .A2(new_n328_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n340_));
  INV_X1    g139(.A(G120gat), .ZN(new_n341_));
  OR2_X1    g140(.A1(G127gat), .A2(G134gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G127gat), .A2(G134gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  AND2_X1   g144(.A1(G127gat), .A2(G134gat), .ZN(new_n346_));
  NOR2_X1   g145(.A1(G127gat), .A2(G134gat), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT76), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(G113gat), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n345_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n349_), .B1(new_n345_), .B2(new_n348_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n341_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NOR3_X1   g151(.A1(new_n346_), .A2(new_n347_), .A3(KEYINPUT76), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n343_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n354_));
  OAI21_X1  g153(.A(G113gat), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n345_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n355_), .A2(G120gat), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n352_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n339_), .A2(new_n340_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n358_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n336_), .B(new_n338_), .C1(new_n360_), .C2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n339_), .A2(new_n340_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n358_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n329_), .A2(new_n337_), .A3(new_n334_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n337_), .B1(new_n329_), .B2(new_n334_), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n359_), .B(new_n365_), .C1(new_n366_), .C2(new_n367_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n362_), .A2(new_n368_), .A3(KEYINPUT77), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT77), .B1(new_n362_), .B2(new_n368_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT83), .B1(new_n294_), .B2(G204gat), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT83), .ZN(new_n373_));
  INV_X1    g172(.A(G204gat), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(new_n374_), .A3(G197gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n372_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT21), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n294_), .A2(G204gat), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n376_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT84), .ZN(new_n380_));
  AOI22_X1  g179(.A1(new_n372_), .A2(new_n375_), .B1(new_n294_), .B2(G204gat), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT84), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n381_), .A2(new_n382_), .A3(new_n377_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT85), .ZN(new_n384_));
  AND2_X1   g183(.A1(G211gat), .A2(G218gat), .ZN(new_n385_));
  NOR2_X1   g184(.A1(G211gat), .A2(G218gat), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n384_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n386_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G211gat), .A2(G218gat), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(KEYINPUT85), .A3(new_n389_), .ZN(new_n390_));
  AOI22_X1  g189(.A1(new_n380_), .A2(new_n383_), .B1(new_n387_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT82), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n378_), .A2(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n393_), .B1(new_n294_), .B2(G204gat), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n378_), .A2(new_n392_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT21), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n376_), .A2(new_n378_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT87), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT87), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n381_), .A2(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n377_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n390_), .A2(new_n387_), .A3(KEYINPUT86), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT86), .B1(new_n390_), .B2(new_n387_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  AOI22_X1  g203(.A1(new_n391_), .A2(new_n396_), .B1(new_n401_), .B2(new_n404_), .ZN(new_n405_));
  OAI211_X1 g204(.A(G228gat), .B(G233gat), .C1(new_n405_), .C2(KEYINPUT88), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT29), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT3), .ZN(new_n408_));
  INV_X1    g207(.A(G141gat), .ZN(new_n409_));
  INV_X1    g208(.A(G148gat), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n408_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G141gat), .A2(G148gat), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT2), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n411_), .A2(new_n414_), .A3(new_n415_), .A4(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT79), .ZN(new_n418_));
  AND2_X1   g217(.A1(G155gat), .A2(G162gat), .ZN(new_n419_));
  NOR2_X1   g218(.A1(G155gat), .A2(G162gat), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n418_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(G155gat), .ZN(new_n422_));
  INV_X1    g221(.A(G162gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G155gat), .A2(G162gat), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n424_), .A2(KEYINPUT79), .A3(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n417_), .A2(new_n421_), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT80), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n417_), .A2(KEYINPUT80), .A3(new_n421_), .A4(new_n426_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n409_), .A2(new_n410_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT1), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT78), .B1(new_n419_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT78), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n425_), .A2(new_n435_), .A3(KEYINPUT1), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n434_), .A2(new_n424_), .A3(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n425_), .A2(KEYINPUT1), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n412_), .B(new_n432_), .C1(new_n437_), .C2(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n407_), .B1(new_n431_), .B2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G78gat), .B(G106gat), .ZN(new_n441_));
  NOR3_X1   g240(.A1(new_n405_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n441_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n421_), .A2(new_n426_), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT80), .B1(new_n444_), .B2(new_n417_), .ZN(new_n445_));
  AND4_X1   g244(.A1(KEYINPUT80), .A2(new_n417_), .A3(new_n421_), .A4(new_n426_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n439_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT29), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n398_), .A2(new_n400_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n404_), .A2(new_n449_), .A3(KEYINPUT21), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n390_), .A2(new_n387_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n379_), .A2(KEYINPUT84), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n382_), .B1(new_n381_), .B2(new_n377_), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n396_), .B(new_n451_), .C1(new_n452_), .C2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n450_), .A2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n443_), .B1(new_n448_), .B2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n406_), .B1(new_n442_), .B2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n441_), .B1(new_n405_), .B2(new_n440_), .ZN(new_n458_));
  INV_X1    g257(.A(G228gat), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT88), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n459_), .B1(new_n455_), .B2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n448_), .A2(new_n455_), .A3(new_n443_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n458_), .A2(new_n461_), .A3(new_n462_), .A4(G233gat), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n457_), .A2(new_n463_), .A3(KEYINPUT81), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT28), .B1(new_n447_), .B2(KEYINPUT29), .ZN(new_n465_));
  XOR2_X1   g264(.A(G22gat), .B(G50gat), .Z(new_n466_));
  INV_X1    g265(.A(KEYINPUT28), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n431_), .A2(new_n467_), .A3(new_n407_), .A4(new_n439_), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n465_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n466_), .B1(new_n465_), .B2(new_n468_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n464_), .A2(new_n472_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n471_), .A2(new_n457_), .A3(KEYINPUT81), .A4(new_n463_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n371_), .A2(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(G57gat), .B(G85gat), .Z(new_n478_));
  XNOR2_X1  g277(.A(G1gat), .B(G29gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n480_), .B(new_n481_), .Z(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n447_), .A2(new_n358_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n431_), .A2(new_n357_), .A3(new_n352_), .A4(new_n439_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n484_), .A2(KEYINPUT4), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT92), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G225gat), .A2(G233gat), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n484_), .A2(KEYINPUT4), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT92), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n484_), .A2(new_n485_), .A3(new_n491_), .A4(KEYINPUT4), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n487_), .A2(new_n489_), .A3(new_n490_), .A4(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT93), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n484_), .A2(new_n485_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(new_n488_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n494_), .B1(new_n493_), .B2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n483_), .B1(new_n495_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT96), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n493_), .A2(new_n494_), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n493_), .A2(new_n497_), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n482_), .B(new_n501_), .C1(new_n502_), .C2(new_n494_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT96), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n504_), .B(new_n483_), .C1(new_n495_), .C2(new_n498_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n500_), .A2(new_n503_), .A3(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT91), .B(KEYINPUT24), .ZN(new_n507_));
  INV_X1    g306(.A(new_n310_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n310_), .A2(new_n312_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n509_), .B1(new_n507_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n303_), .A2(new_n308_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n318_), .A2(new_n312_), .ZN(new_n514_));
  AOI22_X1  g313(.A1(new_n512_), .A2(new_n513_), .B1(new_n514_), .B2(new_n317_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n450_), .A2(new_n454_), .A3(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n321_), .A2(new_n322_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n516_), .B(KEYINPUT20), .C1(new_n405_), .C2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT95), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G226gat), .A2(G233gat), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n520_), .B(KEYINPUT90), .Z(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT89), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT19), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  AND3_X1   g324(.A1(new_n518_), .A2(new_n519_), .A3(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n519_), .B1(new_n518_), .B2(new_n525_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n515_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n455_), .A2(new_n528_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n450_), .A2(new_n454_), .A3(new_n326_), .A4(new_n320_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n529_), .A2(new_n524_), .A3(KEYINPUT20), .A4(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NOR3_X1   g331(.A1(new_n526_), .A2(new_n527_), .A3(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G8gat), .B(G36gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT18), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(G64gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(G92gat), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT32), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n533_), .A2(new_n539_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n525_), .A2(KEYINPUT20), .A3(new_n530_), .A4(new_n529_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n518_), .A2(new_n524_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n540_), .B1(new_n543_), .B2(new_n539_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n506_), .A2(new_n544_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n487_), .A2(new_n488_), .A3(new_n490_), .A4(new_n492_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n496_), .A2(new_n489_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n546_), .A2(new_n483_), .A3(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n543_), .A2(new_n538_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n543_), .A2(new_n538_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT33), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n495_), .A2(new_n498_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n553_), .B1(new_n554_), .B2(new_n482_), .ZN(new_n555_));
  NOR4_X1   g354(.A1(new_n495_), .A2(new_n498_), .A3(KEYINPUT33), .A4(new_n483_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n548_), .B(new_n552_), .C1(new_n555_), .C2(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n477_), .B1(new_n545_), .B2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n362_), .A2(new_n368_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n475_), .A2(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n560_), .B1(new_n371_), .B2(new_n475_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT97), .B1(new_n533_), .B2(new_n538_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n518_), .A2(new_n525_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT95), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n518_), .A2(new_n519_), .A3(new_n525_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n564_), .A2(new_n531_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT97), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(new_n567_), .A3(new_n537_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n562_), .A2(KEYINPUT27), .A3(new_n549_), .A4(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT98), .B(KEYINPUT27), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n570_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  NOR3_X1   g371(.A1(new_n561_), .A2(new_n572_), .A3(new_n506_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n300_), .B1(new_n558_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(KEYINPUT99), .ZN(new_n575_));
  INV_X1    g374(.A(new_n506_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n569_), .A2(new_n571_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT77), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n559_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n362_), .A2(new_n368_), .A3(KEYINPUT77), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n579_), .A2(new_n475_), .A3(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n581_), .B1(new_n475_), .B2(new_n559_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n576_), .A2(new_n577_), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n552_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n503_), .A2(KEYINPUT33), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n554_), .A2(new_n553_), .A3(new_n482_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n584_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  AOI22_X1  g386(.A1(new_n587_), .A2(new_n548_), .B1(new_n506_), .B2(new_n544_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n583_), .B1(new_n588_), .B2(new_n477_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT99), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n589_), .A2(new_n590_), .A3(new_n300_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n265_), .B1(new_n575_), .B2(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(G190gat), .B(G218gat), .Z(new_n593_));
  XNOR2_X1  g392(.A(G134gat), .B(G162gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(KEYINPUT36), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT36), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n283_), .A2(new_n238_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n238_), .A2(new_n269_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G232gat), .A2(G233gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT68), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT34), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT35), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n598_), .A2(new_n599_), .A3(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n602_), .A2(new_n603_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n606_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n598_), .A2(new_n599_), .A3(new_n608_), .A4(new_n604_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n597_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n596_), .B1(new_n610_), .B2(new_n595_), .ZN(new_n611_));
  AOI21_X1  g410(.A(KEYINPUT69), .B1(new_n607_), .B2(new_n609_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n612_), .ZN(new_n614_));
  OAI211_X1 g413(.A(new_n614_), .B(new_n596_), .C1(new_n610_), .C2(new_n595_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT37), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n613_), .A2(new_n615_), .A3(KEYINPUT37), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(G231gat), .A2(G233gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n276_), .B(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(new_n239_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G183gat), .B(G211gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G127gat), .B(G155gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  XOR2_X1   g425(.A(KEYINPUT71), .B(KEYINPUT16), .Z(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT17), .ZN(new_n629_));
  OR3_X1    g428(.A1(new_n628_), .A2(KEYINPUT70), .A3(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n623_), .A2(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n623_), .B1(new_n629_), .B2(new_n628_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n631_), .B1(new_n633_), .B2(new_n630_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n620_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n592_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n637_), .A2(new_n271_), .A3(new_n506_), .ZN(new_n638_));
  XOR2_X1   g437(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  OR3_X1    g439(.A1(new_n638_), .A2(KEYINPUT101), .A3(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n558_), .A2(new_n573_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n265_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n299_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n616_), .ZN(new_n646_));
  NOR4_X1   g445(.A1(new_n642_), .A2(new_n645_), .A3(new_n634_), .A4(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n271_), .B1(new_n647_), .B2(new_n506_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n638_), .B1(new_n648_), .B2(new_n640_), .ZN(new_n649_));
  OAI21_X1  g448(.A(KEYINPUT101), .B1(new_n638_), .B2(new_n640_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n641_), .A2(new_n649_), .A3(new_n650_), .ZN(G1324gat));
  NAND3_X1  g450(.A1(new_n637_), .A2(new_n272_), .A3(new_n572_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n272_), .B1(new_n647_), .B2(new_n572_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n653_), .A2(new_n654_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n652_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g458(.A(G15gat), .ZN(new_n660_));
  INV_X1    g459(.A(new_n371_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n647_), .B2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT41), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n637_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(G1326gat));
  INV_X1    g466(.A(G22gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n668_), .B1(new_n647_), .B2(new_n475_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT42), .Z(new_n670_));
  NAND2_X1  g469(.A1(new_n475_), .A2(new_n668_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n670_), .B1(new_n636_), .B2(new_n671_), .ZN(G1327gat));
  INV_X1    g471(.A(new_n645_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n589_), .B2(new_n620_), .ZN(new_n675_));
  OAI211_X1 g474(.A(new_n674_), .B(new_n620_), .C1(new_n558_), .C2(new_n573_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n634_), .B(new_n673_), .C1(new_n675_), .C2(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(KEYINPUT103), .A2(KEYINPUT44), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n620_), .B1(new_n558_), .B2(new_n573_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT43), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n645_), .B1(new_n683_), .B2(new_n676_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(new_n634_), .A3(new_n679_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n576_), .B1(new_n681_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(G29gat), .ZN(new_n687_));
  INV_X1    g486(.A(new_n634_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n616_), .A2(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT104), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n592_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n506_), .A2(new_n687_), .ZN(new_n692_));
  OAI22_X1  g491(.A1(new_n686_), .A2(new_n687_), .B1(new_n691_), .B2(new_n692_), .ZN(G1328gat));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n694_));
  INV_X1    g493(.A(G36gat), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n592_), .A2(new_n695_), .A3(new_n572_), .A4(new_n690_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n696_), .B(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n681_), .A2(new_n685_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n695_), .B1(new_n700_), .B2(new_n572_), .ZN(new_n701_));
  OAI211_X1 g500(.A(new_n694_), .B(KEYINPUT46), .C1(new_n699_), .C2(new_n701_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n678_), .A2(new_n680_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n679_), .B1(new_n684_), .B2(new_n634_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n572_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(G36gat), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n696_), .B(new_n697_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n694_), .A2(KEYINPUT46), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n694_), .A2(KEYINPUT46), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n706_), .A2(new_n707_), .A3(new_n708_), .A4(new_n709_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n702_), .A2(new_n710_), .ZN(G1329gat));
  INV_X1    g510(.A(new_n559_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n700_), .A2(G43gat), .A3(new_n712_), .ZN(new_n713_));
  XOR2_X1   g512(.A(KEYINPUT107), .B(G43gat), .Z(new_n714_));
  OAI21_X1  g513(.A(new_n714_), .B1(new_n691_), .B2(new_n371_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g516(.A(new_n476_), .B1(new_n681_), .B2(new_n685_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n475_), .A2(new_n278_), .ZN(new_n719_));
  OAI22_X1  g518(.A1(new_n718_), .A2(new_n278_), .B1(new_n691_), .B2(new_n719_), .ZN(G1331gat));
  NOR2_X1   g519(.A1(new_n643_), .A2(new_n644_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n589_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(new_n635_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(G57gat), .B1(new_n724_), .B2(new_n506_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n300_), .A2(new_n634_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n589_), .A2(new_n616_), .A3(new_n265_), .A4(new_n726_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT108), .Z(new_n728_));
  AND2_X1   g527(.A1(new_n506_), .A2(G57gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(G1332gat));
  OR3_X1    g529(.A1(new_n723_), .A2(G64gat), .A3(new_n577_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n728_), .A2(new_n572_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT48), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n732_), .A2(new_n733_), .A3(G64gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n732_), .B2(G64gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n731_), .B1(new_n734_), .B2(new_n735_), .ZN(G1333gat));
  INV_X1    g535(.A(KEYINPUT49), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n728_), .A2(new_n661_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n738_), .B2(G71gat), .ZN(new_n739_));
  INV_X1    g538(.A(G71gat), .ZN(new_n740_));
  AOI211_X1 g539(.A(KEYINPUT49), .B(new_n740_), .C1(new_n728_), .C2(new_n661_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n661_), .A2(new_n740_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT109), .ZN(new_n743_));
  OAI22_X1  g542(.A1(new_n739_), .A2(new_n741_), .B1(new_n723_), .B2(new_n743_), .ZN(G1334gat));
  OR3_X1    g543(.A1(new_n723_), .A2(G78gat), .A3(new_n476_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n728_), .A2(new_n475_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n746_), .A2(G78gat), .A3(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n746_), .B2(G78gat), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n745_), .B1(new_n749_), .B2(new_n750_), .ZN(G1335gat));
  NAND2_X1  g550(.A1(new_n722_), .A2(new_n690_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(G85gat), .B1(new_n753_), .B2(new_n506_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n721_), .A2(new_n634_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n683_), .B2(new_n676_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n757_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n576_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n754_), .B1(new_n760_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g560(.A(G92gat), .B1(new_n753_), .B2(new_n572_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n577_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(G92gat), .ZN(G1337gat));
  NAND2_X1  g563(.A1(new_n756_), .A2(new_n661_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(G99gat), .ZN(new_n766_));
  XOR2_X1   g565(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n767_));
  NAND2_X1  g566(.A1(new_n712_), .A2(new_n231_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n766_), .B(new_n767_), .C1(new_n752_), .C2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT114), .ZN(new_n770_));
  INV_X1    g569(.A(new_n766_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n752_), .A2(new_n768_), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT51), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT112), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n773_), .A2(new_n774_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n770_), .B1(new_n775_), .B2(new_n776_), .ZN(G1338gat));
  NAND3_X1  g576(.A1(new_n753_), .A2(new_n232_), .A3(new_n475_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n755_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n475_), .B(new_n779_), .C1(new_n675_), .C2(new_n677_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n780_), .A2(new_n781_), .A3(G106gat), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n780_), .B2(G106gat), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n782_), .A2(new_n783_), .A3(KEYINPUT52), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785_));
  AOI211_X1 g584(.A(new_n476_), .B(new_n755_), .C1(new_n683_), .C2(new_n676_), .ZN(new_n786_));
  OAI21_X1  g585(.A(KEYINPUT115), .B1(new_n786_), .B2(new_n232_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n780_), .A2(new_n781_), .A3(G106gat), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n785_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n778_), .B1(new_n784_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT53), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n792_), .B(new_n778_), .C1(new_n784_), .C2(new_n789_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(G1339gat));
  NOR2_X1   g593(.A1(new_n265_), .A2(new_n300_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n795_), .A2(new_n688_), .A3(new_n619_), .A4(new_n618_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n796_), .B(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n299_), .B1(new_n250_), .B2(new_n255_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n800_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n801_));
  AOI211_X1 g600(.A(KEYINPUT55), .B(new_n248_), .C1(new_n241_), .C2(new_n243_), .ZN(new_n802_));
  OAI22_X1  g601(.A1(new_n801_), .A2(new_n802_), .B1(new_n245_), .B2(new_n244_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n803_), .A2(KEYINPUT116), .A3(KEYINPUT56), .A4(new_n256_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n799_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT56), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n244_), .A2(new_n245_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n246_), .A2(KEYINPUT55), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n244_), .A2(new_n800_), .A3(new_n245_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n807_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n806_), .B1(new_n810_), .B2(new_n255_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n803_), .A2(KEYINPUT56), .A3(new_n256_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n811_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n805_), .A2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n296_), .B1(new_n288_), .B2(new_n285_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT117), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n284_), .A2(new_n289_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n297_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n261_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n815_), .A2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n821_), .A2(KEYINPUT57), .A3(new_n616_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT118), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n824_));
  AOI22_X1  g623(.A1(new_n805_), .A2(new_n814_), .B1(new_n261_), .B2(new_n819_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n825_), .B2(new_n646_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n811_), .A2(new_n813_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n250_), .A2(new_n255_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n827_), .A2(new_n819_), .A3(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT58), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n827_), .A2(KEYINPUT58), .A3(new_n819_), .A4(new_n828_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n620_), .A3(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n646_), .B1(new_n815_), .B2(new_n820_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n834_), .A2(new_n835_), .A3(KEYINPUT57), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n823_), .A2(new_n826_), .A3(new_n833_), .A4(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n798_), .B1(new_n837_), .B2(new_n634_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n576_), .A2(new_n572_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n560_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(KEYINPUT119), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n838_), .A2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(G113gat), .B1(new_n843_), .B2(new_n644_), .ZN(new_n844_));
  XOR2_X1   g643(.A(KEYINPUT121), .B(G113gat), .Z(new_n845_));
  INV_X1    g644(.A(KEYINPUT120), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT59), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n846_), .B(new_n847_), .C1(new_n838_), .C2(new_n842_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n798_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n826_), .A2(new_n833_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n835_), .B1(new_n834_), .B2(KEYINPUT57), .ZN(new_n851_));
  NOR4_X1   g650(.A1(new_n825_), .A2(KEYINPUT118), .A3(new_n824_), .A4(new_n646_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n850_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n849_), .B1(new_n853_), .B2(new_n688_), .ZN(new_n854_));
  XOR2_X1   g653(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n855_));
  NAND3_X1  g654(.A1(new_n854_), .A2(new_n841_), .A3(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n845_), .B1(new_n848_), .B2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n844_), .B1(new_n857_), .B2(new_n300_), .ZN(G1340gat));
  INV_X1    g657(.A(KEYINPUT60), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n643_), .B2(G120gat), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n854_), .A2(new_n841_), .A3(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n846_), .A2(new_n847_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n862_), .B1(new_n854_), .B2(new_n841_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n855_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n838_), .A2(new_n842_), .A3(new_n864_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n265_), .B(new_n861_), .C1(new_n863_), .C2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(G120gat), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n843_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1341gat));
  INV_X1    g668(.A(G127gat), .ZN(new_n870_));
  AOI211_X1 g669(.A(new_n870_), .B(new_n634_), .C1(new_n848_), .C2(new_n856_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT122), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n843_), .A2(new_n688_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(new_n870_), .ZN(new_n874_));
  AOI211_X1 g673(.A(KEYINPUT122), .B(G127gat), .C1(new_n843_), .C2(new_n688_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n871_), .A2(new_n874_), .A3(new_n875_), .ZN(G1342gat));
  AOI21_X1  g675(.A(G134gat), .B1(new_n843_), .B2(new_n646_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n620_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n878_), .B1(new_n848_), .B2(new_n856_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n877_), .B1(new_n879_), .B2(G134gat), .ZN(G1343gat));
  NOR2_X1   g679(.A1(new_n838_), .A2(new_n581_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n839_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n883_), .A2(new_n409_), .A3(new_n644_), .ZN(new_n884_));
  OAI21_X1  g683(.A(G141gat), .B1(new_n882_), .B2(new_n299_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1344gat));
  NAND3_X1  g685(.A1(new_n883_), .A2(new_n410_), .A3(new_n265_), .ZN(new_n887_));
  OAI21_X1  g686(.A(G148gat), .B1(new_n882_), .B2(new_n643_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1345gat));
  XNOR2_X1  g688(.A(KEYINPUT61), .B(G155gat), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n890_), .B1(new_n883_), .B2(new_n688_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n890_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n882_), .A2(new_n634_), .A3(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n891_), .A2(new_n893_), .ZN(G1346gat));
  NOR3_X1   g693(.A1(new_n882_), .A2(new_n423_), .A3(new_n878_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n883_), .A2(new_n646_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n895_), .B1(new_n423_), .B2(new_n896_), .ZN(G1347gat));
  INV_X1    g696(.A(KEYINPUT124), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n577_), .A2(new_n506_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n661_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n644_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n902_), .B(new_n903_), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n838_), .A2(new_n475_), .A3(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n898_), .B1(new_n905_), .B2(new_n292_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n854_), .A2(new_n476_), .ZN(new_n907_));
  OAI211_X1 g706(.A(KEYINPUT124), .B(G169gat), .C1(new_n907_), .C2(new_n904_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n906_), .A2(new_n908_), .A3(KEYINPUT62), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n838_), .A2(new_n475_), .ZN(new_n910_));
  NAND4_X1  g709(.A1(new_n910_), .A2(new_n316_), .A3(new_n644_), .A4(new_n901_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n898_), .B(new_n912_), .C1(new_n905_), .C2(new_n292_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n909_), .A2(new_n911_), .A3(new_n913_), .ZN(G1348gat));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n915_), .B1(new_n838_), .B2(new_n475_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n851_), .A2(new_n852_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n850_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n688_), .B1(new_n917_), .B2(new_n918_), .ZN(new_n919_));
  OAI211_X1 g718(.A(KEYINPUT125), .B(new_n476_), .C1(new_n919_), .C2(new_n798_), .ZN(new_n920_));
  AND3_X1   g719(.A1(new_n916_), .A2(new_n901_), .A3(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n643_), .A2(new_n309_), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n838_), .A2(new_n475_), .A3(new_n900_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n265_), .ZN(new_n924_));
  AOI22_X1  g723(.A1(new_n921_), .A2(new_n922_), .B1(new_n315_), .B2(new_n924_), .ZN(G1349gat));
  NAND4_X1  g724(.A1(new_n916_), .A2(new_n920_), .A3(new_n688_), .A4(new_n901_), .ZN(new_n926_));
  INV_X1    g725(.A(G183gat), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n301_), .ZN(new_n929_));
  NAND4_X1  g728(.A1(new_n854_), .A2(new_n929_), .A3(new_n476_), .A4(new_n901_), .ZN(new_n930_));
  OAI21_X1  g729(.A(KEYINPUT126), .B1(new_n930_), .B2(new_n634_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n932_));
  NAND4_X1  g731(.A1(new_n923_), .A2(new_n932_), .A3(new_n688_), .A4(new_n929_), .ZN(new_n933_));
  AND3_X1   g732(.A1(new_n928_), .A2(new_n931_), .A3(new_n933_), .ZN(G1350gat));
  AND2_X1   g733(.A1(new_n646_), .A2(new_n302_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n910_), .A2(new_n901_), .A3(new_n935_), .ZN(new_n936_));
  NOR4_X1   g735(.A1(new_n838_), .A2(new_n475_), .A3(new_n878_), .A4(new_n900_), .ZN(new_n937_));
  INV_X1    g736(.A(G190gat), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n936_), .B1(new_n937_), .B2(new_n938_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(KEYINPUT127), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT127), .ZN(new_n941_));
  OAI211_X1 g740(.A(new_n936_), .B(new_n941_), .C1(new_n938_), .C2(new_n937_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n940_), .A2(new_n942_), .ZN(G1351gat));
  NAND2_X1  g742(.A1(new_n881_), .A2(new_n899_), .ZN(new_n944_));
  INV_X1    g743(.A(new_n944_), .ZN(new_n945_));
  AOI21_X1  g744(.A(G197gat), .B1(new_n945_), .B2(new_n644_), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n944_), .A2(new_n294_), .A3(new_n299_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n946_), .A2(new_n947_), .ZN(G1352gat));
  NAND3_X1  g747(.A1(new_n945_), .A2(new_n374_), .A3(new_n265_), .ZN(new_n949_));
  OAI21_X1  g748(.A(G204gat), .B1(new_n944_), .B2(new_n643_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n949_), .A2(new_n950_), .ZN(G1353gat));
  XOR2_X1   g750(.A(KEYINPUT63), .B(G211gat), .Z(new_n952_));
  NAND3_X1  g751(.A1(new_n945_), .A2(new_n688_), .A3(new_n952_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n954_), .B1(new_n944_), .B2(new_n634_), .ZN(new_n955_));
  AND2_X1   g754(.A1(new_n953_), .A2(new_n955_), .ZN(G1354gat));
  INV_X1    g755(.A(G218gat), .ZN(new_n957_));
  NOR3_X1   g756(.A1(new_n944_), .A2(new_n957_), .A3(new_n878_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n945_), .A2(new_n646_), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n958_), .B1(new_n957_), .B2(new_n959_), .ZN(G1355gat));
endmodule


