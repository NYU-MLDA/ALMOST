//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n904_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_;
  INV_X1    g000(.A(KEYINPUT67), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G230gat), .A2(G233gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT64), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT10), .B(G99gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G85gat), .A2(G92gat), .ZN(new_n206_));
  OAI22_X1  g005(.A1(new_n205_), .A2(G106gat), .B1(KEYINPUT9), .B2(new_n206_), .ZN(new_n207_));
  OR2_X1    g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n208_), .A2(KEYINPUT9), .A3(new_n206_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n209_), .A2(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n204_), .B1(new_n207_), .B2(new_n215_), .ZN(new_n216_));
  AND2_X1   g015(.A1(G85gat), .A2(G92gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G85gat), .A2(G92gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  AOI22_X1  g018(.A1(new_n219_), .A2(KEYINPUT9), .B1(new_n211_), .B2(new_n213_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n206_), .A2(KEYINPUT9), .ZN(new_n221_));
  INV_X1    g020(.A(G99gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT10), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT10), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(G99gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(G106gat), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n221_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n220_), .A2(new_n228_), .A3(KEYINPUT64), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n216_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT65), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n231_), .A2(new_n222_), .A3(new_n227_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT7), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT7), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n231_), .A2(new_n234_), .A3(new_n222_), .A4(new_n227_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n214_), .A3(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n236_), .A2(KEYINPUT8), .A3(new_n219_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n219_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT8), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G57gat), .B(G64gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT11), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G71gat), .B(G78gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n241_), .A2(KEYINPUT11), .ZN(new_n245_));
  XOR2_X1   g044(.A(G71gat), .B(G78gat), .Z(new_n246_));
  NAND3_X1  g045(.A1(new_n246_), .A2(KEYINPUT11), .A3(new_n241_), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n244_), .A2(new_n245_), .A3(new_n247_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n230_), .A2(new_n237_), .A3(new_n240_), .A4(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT12), .ZN(new_n250_));
  INV_X1    g049(.A(new_n237_), .ZN(new_n251_));
  AOI21_X1  g050(.A(KEYINPUT8), .B1(new_n236_), .B2(new_n219_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n248_), .B1(new_n253_), .B2(new_n230_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n250_), .A2(new_n254_), .ZN(new_n255_));
  NOR3_X1   g054(.A1(new_n207_), .A2(new_n215_), .A3(new_n204_), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT64), .B1(new_n220_), .B2(new_n228_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n240_), .B(new_n237_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT12), .ZN(new_n259_));
  INV_X1    g058(.A(new_n248_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n258_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n203_), .B1(new_n255_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n258_), .A2(new_n260_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT66), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n264_), .A2(new_n265_), .A3(new_n249_), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n230_), .A2(new_n237_), .A3(new_n240_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n267_), .A2(KEYINPUT66), .A3(new_n248_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n203_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n266_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n202_), .B1(new_n263_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n202_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G120gat), .B(G148gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT5), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(G176gat), .ZN(new_n276_));
  INV_X1    g075(.A(G204gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  NOR3_X1   g077(.A1(new_n271_), .A2(new_n273_), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n278_), .ZN(new_n280_));
  AND3_X1   g079(.A1(new_n266_), .A2(new_n269_), .A3(new_n268_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n264_), .A2(KEYINPUT12), .A3(new_n249_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n269_), .B1(new_n282_), .B2(new_n261_), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT67), .B1(new_n281_), .B2(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n280_), .B1(new_n284_), .B2(new_n272_), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n279_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT13), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G64gat), .B(G92gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G8gat), .B(G36gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n292_));
  XOR2_X1   g091(.A(new_n291_), .B(new_n292_), .Z(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G211gat), .B(G218gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n277_), .A2(G197gat), .ZN(new_n296_));
  INV_X1    g095(.A(G197gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G204gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n299_), .A2(KEYINPUT21), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n277_), .A2(KEYINPUT82), .A3(G197gat), .ZN(new_n301_));
  OAI211_X1 g100(.A(KEYINPUT21), .B(new_n301_), .C1(new_n299_), .C2(KEYINPUT82), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT83), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n302_), .A2(new_n303_), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n295_), .B(new_n300_), .C1(new_n304_), .C2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n295_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n307_), .A2(KEYINPUT21), .A3(new_n299_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT23), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n310_), .A2(G183gat), .A3(G190gat), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT75), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(G183gat), .ZN(new_n314_));
  INV_X1    g113(.A(G190gat), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT23), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n310_), .A2(KEYINPUT75), .A3(G183gat), .A4(G190gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n313_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n318_), .B1(G183gat), .B2(G190gat), .ZN(new_n319_));
  NOR2_X1   g118(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(G169gat), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  OR2_X1    g121(.A1(G169gat), .A2(G176gat), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n323_), .A2(KEYINPUT24), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n316_), .A2(new_n311_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G169gat), .A2(G176gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n323_), .A2(KEYINPUT24), .A3(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n324_), .A2(new_n325_), .A3(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT26), .B(G190gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT25), .B(G183gat), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n328_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n322_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n309_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G226gat), .A2(G233gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT19), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n318_), .A2(new_n324_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT76), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT74), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT26), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n338_), .B1(new_n339_), .B2(G190gat), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n340_), .B(new_n330_), .C1(new_n329_), .C2(new_n338_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT76), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n318_), .A2(new_n342_), .A3(new_n324_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n337_), .A2(new_n341_), .A3(new_n343_), .A4(new_n327_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n325_), .B1(G183gat), .B2(G190gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(new_n321_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n306_), .A2(new_n344_), .A3(new_n346_), .A4(new_n308_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n333_), .A2(KEYINPUT20), .A3(new_n335_), .A4(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT20), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n344_), .A2(new_n346_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n350_), .B1(new_n309_), .B2(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n322_), .A2(new_n331_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n353_), .A2(new_n306_), .A3(new_n308_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n335_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n294_), .B1(new_n349_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n335_), .ZN(new_n357_));
  AND4_X1   g156(.A1(KEYINPUT20), .A2(new_n333_), .A3(new_n357_), .A4(new_n347_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n357_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n293_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n356_), .A2(new_n360_), .A3(KEYINPUT27), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n352_), .A2(new_n354_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(new_n357_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(new_n348_), .A3(new_n293_), .ZN(new_n364_));
  AOI21_X1  g163(.A(KEYINPUT27), .B1(new_n356_), .B2(new_n364_), .ZN(new_n365_));
  NOR3_X1   g164(.A1(new_n361_), .A2(new_n365_), .A3(KEYINPUT93), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT93), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT27), .ZN(new_n368_));
  NOR3_X1   g167(.A1(new_n349_), .A2(new_n355_), .A3(new_n294_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n293_), .B1(new_n363_), .B2(new_n348_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n368_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n356_), .A2(new_n360_), .A3(KEYINPUT27), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n367_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n366_), .A2(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(G155gat), .A2(G162gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT78), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT3), .ZN(new_n377_));
  INV_X1    g176(.A(G141gat), .ZN(new_n378_));
  INV_X1    g177(.A(G148gat), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n377_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G141gat), .A2(G148gat), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT2), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n380_), .A2(new_n383_), .A3(new_n384_), .A4(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G155gat), .A2(G162gat), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n376_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n378_), .A2(new_n379_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n381_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT1), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n387_), .B(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n390_), .B1(new_n376_), .B2(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n388_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT29), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT79), .B(KEYINPUT28), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G22gat), .B(G50gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT29), .B1(new_n388_), .B2(new_n393_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n309_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G228gat), .A2(G233gat), .ZN(new_n403_));
  XOR2_X1   g202(.A(new_n403_), .B(KEYINPUT81), .Z(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  AOI22_X1  g204(.A1(new_n306_), .A2(new_n308_), .B1(new_n401_), .B2(KEYINPUT80), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT84), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n376_), .A2(new_n392_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n389_), .A2(new_n381_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n376_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n395_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT80), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n404_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n406_), .A2(new_n407_), .A3(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n407_), .B1(new_n406_), .B2(new_n414_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n405_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  XOR2_X1   g216(.A(G78gat), .B(G106gat), .Z(new_n418_));
  XOR2_X1   g217(.A(new_n418_), .B(KEYINPUT85), .Z(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n419_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n405_), .B(new_n421_), .C1(new_n415_), .C2(new_n416_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n420_), .A2(KEYINPUT86), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT86), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n417_), .A2(new_n424_), .A3(new_n419_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n400_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n400_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n418_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n417_), .A2(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n427_), .B1(new_n422_), .B2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT87), .B1(new_n426_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n422_), .A2(KEYINPUT86), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n406_), .A2(new_n414_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT84), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n406_), .A2(new_n407_), .A3(new_n414_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n421_), .B1(new_n436_), .B2(new_n405_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n432_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n425_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n427_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT87), .ZN(new_n441_));
  INV_X1    g240(.A(new_n430_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n374_), .A2(new_n431_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(G120gat), .ZN(new_n445_));
  OR2_X1    g244(.A1(G127gat), .A2(G134gat), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT77), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G127gat), .A2(G134gat), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n446_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n447_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n451_));
  NOR3_X1   g250(.A1(new_n450_), .A2(G113gat), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(G113gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n446_), .A2(new_n448_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT77), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n453_), .B1(new_n455_), .B2(new_n449_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n445_), .B1(new_n452_), .B2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(G113gat), .B1(new_n450_), .B2(new_n451_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n455_), .A2(new_n453_), .A3(new_n449_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(G120gat), .A3(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n457_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n410_), .A2(new_n411_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(KEYINPUT89), .A2(KEYINPUT4), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(KEYINPUT89), .A2(KEYINPUT4), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n461_), .A2(new_n462_), .A3(new_n464_), .A4(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT90), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n461_), .A2(new_n462_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n457_), .A2(new_n394_), .A3(new_n460_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(KEYINPUT4), .A3(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n394_), .B1(new_n457_), .B2(new_n460_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n472_), .A2(KEYINPUT90), .A3(new_n464_), .A4(new_n465_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G225gat), .A2(G233gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n468_), .A2(new_n471_), .A3(new_n473_), .A4(new_n475_), .ZN(new_n476_));
  XOR2_X1   g275(.A(KEYINPUT91), .B(KEYINPUT0), .Z(new_n477_));
  XNOR2_X1  g276(.A(G1gat), .B(G29gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G57gat), .B(G85gat), .ZN(new_n480_));
  XOR2_X1   g279(.A(new_n479_), .B(new_n480_), .Z(new_n481_));
  AND2_X1   g280(.A1(new_n469_), .A2(new_n470_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n474_), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n476_), .A2(new_n481_), .A3(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n481_), .B1(new_n476_), .B2(new_n483_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n351_), .B(new_n461_), .Z(new_n487_));
  XNOR2_X1  g286(.A(G15gat), .B(G43gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT31), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n487_), .B(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G71gat), .B(G99gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT30), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G227gat), .A2(G233gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n490_), .B(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n444_), .A2(KEYINPUT94), .A3(new_n486_), .A4(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT94), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n374_), .A2(new_n486_), .A3(new_n431_), .A4(new_n443_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n498_), .B1(new_n499_), .B2(new_n495_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n369_), .A2(new_n370_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n484_), .A2(KEYINPUT33), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n468_), .A2(new_n471_), .A3(new_n473_), .A4(new_n474_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n481_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n482_), .A2(new_n475_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n504_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n507_), .A2(KEYINPUT33), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n502_), .B(new_n503_), .C1(new_n484_), .C2(new_n508_), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n294_), .A2(KEYINPUT32), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n510_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n349_), .A2(new_n355_), .ZN(new_n512_));
  OAI221_X1 g311(.A(new_n511_), .B1(new_n512_), .B2(new_n510_), .C1(new_n484_), .C2(new_n485_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n509_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n443_), .A2(new_n431_), .A3(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT92), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n361_), .A2(new_n365_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n441_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n426_), .A2(KEYINPUT87), .A3(new_n430_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n486_), .B(new_n517_), .C1(new_n518_), .C2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT92), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n443_), .A2(new_n431_), .A3(new_n514_), .A4(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n516_), .A2(new_n520_), .A3(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n495_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n288_), .B1(new_n501_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT37), .ZN(new_n526_));
  INV_X1    g325(.A(G50gat), .ZN(new_n527_));
  INV_X1    g326(.A(G29gat), .ZN(new_n528_));
  INV_X1    g327(.A(G36gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(G43gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G29gat), .A2(G36gat), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n530_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n531_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n527_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n535_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n537_), .A2(G50gat), .A3(new_n533_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT15), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n258_), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n258_), .A2(new_n539_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G232gat), .A2(G233gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT34), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n545_), .B(KEYINPUT35), .Z(new_n546_));
  NAND3_X1  g345(.A1(new_n542_), .A2(new_n543_), .A3(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT68), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n542_), .A2(new_n543_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(KEYINPUT35), .A3(new_n545_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT68), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n542_), .A2(new_n543_), .A3(new_n551_), .A4(new_n546_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n548_), .A2(new_n550_), .A3(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G190gat), .B(G218gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(G134gat), .ZN(new_n555_));
  INV_X1    g354(.A(G162gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n558_), .A2(KEYINPUT36), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(KEYINPUT36), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n553_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n559_), .B1(new_n553_), .B2(new_n560_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n526_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n563_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n565_), .A2(KEYINPUT37), .A3(new_n561_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G127gat), .B(G155gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT16), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(G183gat), .ZN(new_n570_));
  INV_X1    g369(.A(G211gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT17), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n572_), .A2(new_n573_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G15gat), .B(G22gat), .ZN(new_n576_));
  INV_X1    g375(.A(G1gat), .ZN(new_n577_));
  INV_X1    g376(.A(G8gat), .ZN(new_n578_));
  OAI21_X1  g377(.A(KEYINPUT14), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G1gat), .B(G8gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(new_n260_), .ZN(new_n585_));
  OR3_X1    g384(.A1(new_n574_), .A2(new_n575_), .A3(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n575_), .A2(new_n585_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n567_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT70), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n541_), .A2(new_n590_), .A3(new_n582_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n539_), .A2(new_n540_), .ZN(new_n592_));
  AOI21_X1  g391(.A(KEYINPUT15), .B1(new_n536_), .B2(new_n538_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n582_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT70), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n539_), .A2(new_n582_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G229gat), .A2(G233gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT71), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n591_), .A2(new_n595_), .A3(new_n597_), .A4(new_n600_), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n539_), .A2(new_n582_), .ZN(new_n602_));
  OAI211_X1 g401(.A(G229gat), .B(G233gat), .C1(new_n602_), .C2(new_n596_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT69), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n603_), .A2(KEYINPUT69), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n601_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT72), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G113gat), .B(G141gat), .ZN(new_n608_));
  INV_X1    g407(.A(G169gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(new_n297_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n607_), .A2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n606_), .A2(KEYINPUT72), .A3(new_n611_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT73), .Z(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n525_), .A2(new_n589_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n486_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n618_), .A2(new_n577_), .A3(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT38), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n500_), .A2(new_n497_), .B1(new_n523_), .B2(new_n495_), .ZN(new_n622_));
  AOI21_X1  g421(.A(KEYINPUT96), .B1(new_n565_), .B2(new_n561_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT96), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n562_), .A2(new_n563_), .A3(new_n624_), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n622_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n588_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n287_), .A2(new_n615_), .A3(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(KEYINPUT95), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n629_), .A2(KEYINPUT95), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n627_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G1gat), .B1(new_n632_), .B2(new_n486_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n621_), .A2(new_n633_), .ZN(G1324gat));
  INV_X1    g433(.A(new_n374_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n618_), .A2(new_n578_), .A3(new_n635_), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n632_), .A2(new_n374_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT39), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n637_), .A2(new_n638_), .A3(G8gat), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n637_), .B2(G8gat), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n636_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT40), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(G1325gat));
  INV_X1    g442(.A(G15gat), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n618_), .A2(new_n644_), .A3(new_n496_), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n632_), .A2(new_n495_), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n646_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT41), .B1(new_n646_), .B2(G15gat), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n645_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT97), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(G1326gat));
  INV_X1    g450(.A(G22gat), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n443_), .A2(new_n431_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n618_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n653_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G22gat), .B1(new_n632_), .B2(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(KEYINPUT98), .B(KEYINPUT42), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n656_), .A2(new_n657_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n654_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT99), .Z(G1327gat));
  NAND2_X1  g460(.A1(new_n626_), .A2(new_n588_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(new_n664_));
  NOR4_X1   g463(.A1(new_n622_), .A2(new_n288_), .A3(new_n664_), .A4(new_n616_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(new_n528_), .A3(new_n619_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n615_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668_));
  AOI211_X1 g467(.A(new_n667_), .B(new_n288_), .C1(KEYINPUT100), .C2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT43), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n501_), .A2(new_n524_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n671_), .B2(new_n567_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n567_), .ZN(new_n673_));
  AOI211_X1 g472(.A(KEYINPUT43), .B(new_n673_), .C1(new_n501_), .C2(new_n524_), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n588_), .B(new_n669_), .C1(new_n672_), .C2(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n668_), .A2(KEYINPUT100), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(KEYINPUT43), .B1(new_n622_), .B2(new_n673_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n671_), .A2(new_n670_), .A3(new_n567_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n628_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n676_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n680_), .A2(new_n669_), .A3(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n677_), .A2(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n528_), .B1(new_n683_), .B2(new_n619_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT101), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n684_), .A2(new_n685_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n666_), .B1(new_n686_), .B2(new_n687_), .ZN(G1328gat));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n529_), .B1(new_n683_), .B2(new_n635_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n665_), .A2(new_n691_), .A3(new_n529_), .A4(new_n635_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n664_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n525_), .A2(new_n529_), .A3(new_n617_), .A4(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(KEYINPUT103), .B1(new_n694_), .B2(new_n374_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n692_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT45), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n692_), .A2(new_n695_), .A3(KEYINPUT45), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n689_), .B1(new_n690_), .B2(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  OAI211_X1 g503(.A(new_n689_), .B(new_n702_), .C1(new_n690_), .C2(new_n700_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1329gat));
  NAND3_X1  g505(.A1(new_n683_), .A2(G43gat), .A3(new_n496_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n665_), .A2(new_n496_), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n531_), .A2(KEYINPUT106), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n531_), .A2(KEYINPUT106), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n708_), .A2(new_n709_), .A3(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n707_), .A2(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g512(.A1(new_n665_), .A2(new_n527_), .A3(new_n653_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n655_), .B1(new_n677_), .B2(new_n682_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n714_), .B1(new_n715_), .B2(new_n527_), .ZN(G1331gat));
  AND4_X1   g515(.A1(new_n288_), .A2(new_n627_), .A3(new_n628_), .A4(new_n616_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n717_), .A2(G57gat), .A3(new_n619_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT107), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n719_), .B1(new_n622_), .B2(new_n615_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n671_), .A2(KEYINPUT107), .A3(new_n667_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n720_), .A2(new_n721_), .A3(new_n288_), .A4(new_n589_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n619_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n725_));
  INV_X1    g524(.A(G57gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n724_), .A2(new_n725_), .A3(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n725_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n718_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  OAI211_X1 g531(.A(KEYINPUT109), .B(new_n718_), .C1(new_n728_), .C2(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1332gat));
  INV_X1    g533(.A(G64gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n735_), .B1(new_n717_), .B2(new_n635_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT48), .Z(new_n737_));
  NAND3_X1  g536(.A1(new_n723_), .A2(new_n735_), .A3(new_n635_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1333gat));
  INV_X1    g538(.A(G71gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n717_), .B2(new_n496_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT49), .Z(new_n742_));
  NAND3_X1  g541(.A1(new_n723_), .A2(new_n740_), .A3(new_n496_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1334gat));
  INV_X1    g543(.A(G78gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n717_), .B2(new_n653_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT50), .Z(new_n747_));
  NAND3_X1  g546(.A1(new_n723_), .A2(new_n745_), .A3(new_n653_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1335gat));
  NAND3_X1  g548(.A1(new_n680_), .A2(new_n667_), .A3(new_n288_), .ZN(new_n750_));
  INV_X1    g549(.A(G85gat), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n750_), .A2(new_n751_), .A3(new_n486_), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n720_), .A2(new_n721_), .A3(new_n288_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(new_n693_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n619_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n752_), .B1(new_n756_), .B2(new_n751_), .ZN(G1336gat));
  AOI21_X1  g556(.A(G92gat), .B1(new_n755_), .B2(new_n635_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n750_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n635_), .A2(G92gat), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT110), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n758_), .B1(new_n759_), .B2(new_n761_), .ZN(G1337gat));
  OAI21_X1  g561(.A(G99gat), .B1(new_n750_), .B2(new_n495_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n496_), .A2(new_n226_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n754_), .B2(new_n764_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g565(.A1(new_n680_), .A2(new_n667_), .A3(new_n288_), .A4(new_n653_), .ZN(new_n767_));
  XOR2_X1   g566(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n767_), .A2(G106gat), .A3(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n767_), .B2(G106gat), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n653_), .A2(new_n227_), .ZN(new_n772_));
  OAI22_X1  g571(.A1(new_n770_), .A2(new_n771_), .B1(new_n754_), .B2(new_n772_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n773_), .B(new_n775_), .ZN(G1339gat));
  INV_X1    g575(.A(KEYINPUT117), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n601_), .A2(new_n604_), .A3(new_n605_), .A4(new_n612_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n602_), .A2(new_n596_), .A3(new_n599_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n591_), .A2(new_n595_), .A3(new_n597_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n780_), .B2(new_n599_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n778_), .B1(new_n781_), .B2(new_n612_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n279_), .B2(new_n285_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT114), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n787_), .A2(KEYINPUT113), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n283_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n788_), .ZN(new_n790_));
  AOI211_X1 g589(.A(new_n269_), .B(new_n790_), .C1(new_n282_), .C2(new_n261_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n282_), .A2(new_n269_), .A3(new_n261_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n787_), .A2(KEYINPUT113), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n789_), .A2(new_n791_), .A3(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT56), .B1(new_n795_), .B2(new_n280_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n284_), .A2(new_n272_), .A3(new_n280_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n263_), .A2(new_n790_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n283_), .A2(new_n788_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n798_), .A2(new_n799_), .A3(new_n793_), .A4(new_n792_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT56), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n800_), .A2(new_n801_), .A3(new_n278_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n796_), .A2(new_n615_), .A3(new_n797_), .A4(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(KEYINPUT114), .B(new_n783_), .C1(new_n279_), .C2(new_n285_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n786_), .A2(new_n803_), .A3(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n623_), .A2(new_n625_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(KEYINPUT57), .A3(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(KEYINPUT115), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n805_), .A2(new_n809_), .A3(KEYINPUT57), .A4(new_n806_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n795_), .A2(KEYINPUT56), .A3(new_n280_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n801_), .B1(new_n800_), .B2(new_n278_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n814_), .A2(KEYINPUT58), .A3(new_n797_), .A4(new_n783_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n796_), .A2(new_n797_), .A3(new_n802_), .A4(new_n783_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT58), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n815_), .A2(new_n567_), .A3(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT57), .B1(new_n805_), .B2(new_n806_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n811_), .A2(KEYINPUT116), .A3(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT116), .B1(new_n811_), .B2(new_n821_), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n822_), .A2(new_n823_), .A3(new_n628_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n287_), .A2(new_n589_), .A3(new_n616_), .ZN(new_n825_));
  XOR2_X1   g624(.A(new_n825_), .B(KEYINPUT54), .Z(new_n826_));
  OAI21_X1  g625(.A(new_n777_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n811_), .A2(new_n821_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n811_), .A2(new_n821_), .A3(KEYINPUT116), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n830_), .A2(new_n588_), .A3(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n826_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(KEYINPUT117), .A3(new_n833_), .ZN(new_n834_));
  NOR4_X1   g633(.A1(new_n635_), .A2(new_n653_), .A3(new_n486_), .A4(new_n495_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n827_), .A2(new_n834_), .A3(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT118), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT118), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n827_), .A2(new_n838_), .A3(new_n835_), .A4(new_n834_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(G113gat), .B1(new_n840_), .B2(new_n615_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n828_), .A2(new_n588_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n833_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n844_), .A3(new_n835_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT119), .B1(new_n836_), .B2(KEYINPUT59), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n836_), .A2(KEYINPUT119), .A3(KEYINPUT59), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n846_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n616_), .A2(new_n453_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n841_), .B1(new_n850_), .B2(new_n851_), .ZN(G1340gat));
  AND3_X1   g651(.A1(new_n836_), .A2(KEYINPUT119), .A3(KEYINPUT59), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n288_), .B(new_n845_), .C1(new_n853_), .C2(new_n847_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(G120gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n445_), .B1(new_n287_), .B2(KEYINPUT60), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n445_), .A2(KEYINPUT60), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(KEYINPUT120), .B2(new_n857_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n840_), .B(new_n858_), .C1(KEYINPUT120), .C2(new_n856_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n855_), .A2(new_n859_), .ZN(G1341gat));
  AOI21_X1  g659(.A(G127gat), .B1(new_n840_), .B2(new_n628_), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n628_), .A2(G127gat), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n861_), .B1(new_n850_), .B2(new_n862_), .ZN(G1342gat));
  AOI21_X1  g662(.A(G134gat), .B1(new_n840_), .B2(new_n626_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n567_), .A2(G134gat), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(KEYINPUT121), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n864_), .B1(new_n850_), .B2(new_n866_), .ZN(G1343gat));
  NAND4_X1  g666(.A1(new_n827_), .A2(new_n495_), .A3(new_n653_), .A4(new_n834_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n868_), .A2(new_n486_), .A3(new_n635_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n615_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n288_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g672(.A1(new_n869_), .A2(new_n628_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(KEYINPUT61), .B(G155gat), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1346gat));
  AOI21_X1  g675(.A(G162gat), .B1(new_n869_), .B2(new_n626_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n673_), .A2(new_n556_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n869_), .B2(new_n878_), .ZN(G1347gat));
  NOR2_X1   g678(.A1(new_n374_), .A2(new_n619_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n496_), .ZN(new_n881_));
  XOR2_X1   g680(.A(new_n881_), .B(KEYINPUT122), .Z(new_n882_));
  NAND3_X1  g681(.A1(new_n843_), .A2(new_n655_), .A3(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(G169gat), .B1(new_n883_), .B2(new_n667_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(KEYINPUT62), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n883_), .B(KEYINPUT123), .ZN(new_n886_));
  XNOR2_X1  g685(.A(KEYINPUT22), .B(G169gat), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n615_), .A2(new_n887_), .ZN(new_n888_));
  XOR2_X1   g687(.A(new_n888_), .B(KEYINPUT124), .Z(new_n889_));
  OAI21_X1  g688(.A(new_n885_), .B1(new_n886_), .B2(new_n889_), .ZN(G1348gat));
  INV_X1    g689(.A(new_n886_), .ZN(new_n891_));
  AOI21_X1  g690(.A(G176gat), .B1(new_n891_), .B2(new_n288_), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n827_), .A2(new_n655_), .A3(new_n834_), .ZN(new_n893_));
  AND3_X1   g692(.A1(new_n882_), .A2(G176gat), .A3(new_n288_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n892_), .B1(new_n893_), .B2(new_n894_), .ZN(G1349gat));
  NOR3_X1   g694(.A1(new_n886_), .A2(new_n588_), .A3(new_n330_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n893_), .A2(new_n628_), .A3(new_n882_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n897_), .B2(new_n314_), .ZN(G1350gat));
  OAI21_X1  g697(.A(G190gat), .B1(new_n886_), .B2(new_n673_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n626_), .A2(new_n329_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n886_), .B2(new_n900_), .ZN(G1351gat));
  INV_X1    g700(.A(new_n880_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n868_), .A2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n615_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n288_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g706(.A(KEYINPUT63), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n908_), .A2(new_n571_), .ZN(new_n909_));
  NOR4_X1   g708(.A1(new_n868_), .A2(new_n588_), .A3(new_n902_), .A4(new_n909_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n908_), .A2(new_n571_), .A3(KEYINPUT125), .ZN(new_n911_));
  XOR2_X1   g710(.A(new_n911_), .B(KEYINPUT126), .Z(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(KEYINPUT125), .B1(new_n908_), .B2(new_n571_), .ZN(new_n914_));
  OR3_X1    g713(.A1(new_n910_), .A2(new_n913_), .A3(new_n914_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n913_), .B1(new_n910_), .B2(new_n914_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1354gat));
  XOR2_X1   g716(.A(KEYINPUT127), .B(G218gat), .Z(new_n918_));
  AOI21_X1  g717(.A(new_n918_), .B1(new_n903_), .B2(new_n626_), .ZN(new_n919_));
  AND2_X1   g718(.A1(new_n567_), .A2(new_n918_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n919_), .B1(new_n903_), .B2(new_n920_), .ZN(G1355gat));
endmodule


