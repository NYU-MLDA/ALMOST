//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0 0 1 1 0 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n875_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_;
  XNOR2_X1  g000(.A(G85gat), .B(G92gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n205_), .A2(KEYINPUT7), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT67), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n205_), .A2(KEYINPUT7), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n203_), .B1(new_n208_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT8), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n216_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT10), .B(G99gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(G106gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT9), .ZN(new_n221_));
  OAI22_X1  g020(.A1(new_n219_), .A2(new_n220_), .B1(new_n202_), .B2(new_n221_), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n221_), .A2(G85gat), .A3(G92gat), .ZN(new_n223_));
  NOR3_X1   g022(.A1(new_n222_), .A2(new_n213_), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT66), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n224_), .A2(KEYINPUT66), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n217_), .A2(new_n218_), .A3(new_n225_), .A4(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT12), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G57gat), .B(G64gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT11), .ZN(new_n230_));
  XOR2_X1   g029(.A(G71gat), .B(G78gat), .Z(new_n231_));
  NOR2_X1   g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n230_), .A2(new_n231_), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n229_), .A2(KEYINPUT11), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n232_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n227_), .A2(new_n228_), .A3(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n228_), .B1(new_n227_), .B2(new_n235_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G230gat), .A2(G233gat), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n240_), .B(KEYINPUT64), .Z(new_n241_));
  OAI21_X1  g040(.A(new_n241_), .B1(new_n227_), .B2(new_n235_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  OAI211_X1 g043(.A(KEYINPUT68), .B(new_n241_), .C1(new_n227_), .C2(new_n235_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n239_), .A2(new_n244_), .A3(KEYINPUT69), .A4(new_n245_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n227_), .A2(new_n235_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n227_), .A2(new_n235_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n241_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n245_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n244_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n252_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n246_), .A2(new_n251_), .A3(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G120gat), .B(G148gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT5), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G176gat), .B(G204gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT70), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n256_), .A2(new_n262_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n246_), .A2(new_n255_), .A3(new_n251_), .A4(new_n260_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT13), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT13), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n263_), .A2(new_n267_), .A3(new_n264_), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT71), .B1(new_n266_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n266_), .A2(KEYINPUT71), .A3(new_n268_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT74), .B(KEYINPUT37), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G232gat), .A2(G233gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT35), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n278_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G29gat), .B(G36gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G43gat), .B(G50gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n280_), .B1(new_n227_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n279_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n283_), .B(KEYINPUT15), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n227_), .A2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n289_), .A2(new_n285_), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n287_), .A2(new_n290_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G190gat), .B(G218gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G134gat), .B(G162gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n296_), .B(KEYINPUT36), .Z(new_n297_));
  AND2_X1   g096(.A1(new_n293_), .A2(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n296_), .A2(KEYINPUT36), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n291_), .A2(new_n299_), .A3(new_n292_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n274_), .B1(new_n298_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n293_), .A2(new_n297_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n303_), .A2(new_n300_), .A3(new_n273_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G15gat), .B(G22gat), .ZN(new_n306_));
  INV_X1    g105(.A(G1gat), .ZN(new_n307_));
  INV_X1    g106(.A(G8gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT14), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n306_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G1gat), .B(G8gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(new_n235_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G231gat), .A2(G233gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT17), .ZN(new_n317_));
  XOR2_X1   g116(.A(G127gat), .B(G155gat), .Z(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT16), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G183gat), .B(G211gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  OR3_X1    g120(.A1(new_n316_), .A2(new_n317_), .A3(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(KEYINPUT17), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n316_), .A2(new_n323_), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n305_), .A2(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n272_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT107), .ZN(new_n328_));
  INV_X1    g127(.A(G141gat), .ZN(new_n329_));
  INV_X1    g128(.A(G148gat), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n329_), .A2(new_n330_), .A3(KEYINPUT3), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT3), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n332_), .B1(G141gat), .B2(G148gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  AND3_X1   g133(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n335_));
  AOI21_X1  g134(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n334_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT85), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n334_), .A2(new_n337_), .A3(KEYINPUT85), .ZN(new_n341_));
  NOR2_X1   g140(.A1(G155gat), .A2(G162gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT86), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n345_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT86), .B1(new_n347_), .B2(new_n342_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n340_), .A2(new_n341_), .A3(new_n346_), .A4(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n329_), .A2(new_n330_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G141gat), .A2(G148gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n345_), .A2(KEYINPUT1), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n345_), .B1(new_n342_), .B2(KEYINPUT1), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT83), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n353_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  OAI211_X1 g155(.A(KEYINPUT83), .B(new_n345_), .C1(new_n342_), .C2(KEYINPUT1), .ZN(new_n357_));
  AOI211_X1 g156(.A(KEYINPUT84), .B(new_n352_), .C1(new_n356_), .C2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT84), .ZN(new_n359_));
  INV_X1    g158(.A(G155gat), .ZN(new_n360_));
  INV_X1    g159(.A(G162gat), .ZN(new_n361_));
  AOI21_X1  g160(.A(KEYINPUT1), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n355_), .B1(new_n362_), .B2(new_n347_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n353_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n363_), .A2(new_n357_), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n352_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n359_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n349_), .B1(new_n358_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT87), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT87), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n370_), .B(new_n349_), .C1(new_n358_), .C2(new_n367_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G127gat), .B(G134gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G113gat), .B(G120gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n369_), .A2(new_n371_), .A3(new_n375_), .ZN(new_n376_));
  AND3_X1   g175(.A1(new_n334_), .A2(new_n337_), .A3(KEYINPUT85), .ZN(new_n377_));
  AOI21_X1  g176(.A(KEYINPUT85), .B1(new_n334_), .B2(new_n337_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n346_), .A2(new_n348_), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n377_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n365_), .A2(new_n366_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT84), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n365_), .A2(new_n359_), .A3(new_n366_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n380_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n375_), .A2(KEYINPUT101), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n375_), .A2(KEYINPUT101), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n384_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n376_), .A2(new_n387_), .A3(KEYINPUT4), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT4), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n369_), .A2(new_n389_), .A3(new_n371_), .A4(new_n375_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G225gat), .A2(G233gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT102), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n388_), .A2(new_n390_), .A3(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n376_), .A2(new_n387_), .A3(new_n391_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  XOR2_X1   g194(.A(G1gat), .B(G29gat), .Z(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT103), .B(KEYINPUT0), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G57gat), .B(G85gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n395_), .A2(new_n401_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n394_), .A2(new_n400_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(new_n393_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(G197gat), .A2(G204gat), .ZN(new_n406_));
  XOR2_X1   g205(.A(KEYINPUT90), .B(G204gat), .Z(new_n407_));
  AOI21_X1  g206(.A(new_n406_), .B1(new_n407_), .B2(G197gat), .ZN(new_n408_));
  XOR2_X1   g207(.A(G211gat), .B(G218gat), .Z(new_n409_));
  NAND4_X1  g208(.A1(new_n408_), .A2(KEYINPUT92), .A3(KEYINPUT21), .A4(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT92), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(KEYINPUT21), .ZN(new_n412_));
  INV_X1    g211(.A(new_n406_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT90), .B(G204gat), .ZN(new_n414_));
  INV_X1    g213(.A(G197gat), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n413_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n411_), .B1(new_n412_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n410_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(G204gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(G197gat), .ZN(new_n420_));
  OAI211_X1 g219(.A(KEYINPUT91), .B(new_n420_), .C1(new_n414_), .C2(G197gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n407_), .A2(new_n415_), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n421_), .B(KEYINPUT21), .C1(new_n422_), .C2(KEYINPUT91), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT21), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n409_), .B1(new_n416_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n418_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(G169gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT22), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT22), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(G169gat), .ZN(new_n431_));
  INV_X1    g230(.A(G176gat), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n429_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT78), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT22), .B(G169gat), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(KEYINPUT78), .A3(new_n432_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(G183gat), .ZN(new_n439_));
  INV_X1    g238(.A(G190gat), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT23), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT23), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n442_), .A2(G183gat), .A3(G190gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n441_), .A2(KEYINPUT79), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT79), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n445_), .B(KEYINPUT23), .C1(new_n439_), .C2(new_n440_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n439_), .A2(new_n440_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n444_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G169gat), .A2(G176gat), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n438_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  OR3_X1    g249(.A1(KEYINPUT77), .A2(G169gat), .A3(G176gat), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT77), .B1(G169gat), .B2(G176gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT24), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT25), .B(G183gat), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT26), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT76), .B1(new_n457_), .B2(G190gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT26), .B(G190gat), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n456_), .B(new_n458_), .C1(new_n459_), .C2(KEYINPUT76), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n451_), .A2(KEYINPUT24), .A3(new_n449_), .A4(new_n452_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n441_), .A2(new_n443_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n455_), .A2(new_n460_), .A3(new_n461_), .A4(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n450_), .A2(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT20), .B1(new_n427_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT97), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G226gat), .A2(G233gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT19), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n444_), .A2(new_n446_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n459_), .A2(new_n456_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n471_), .A2(new_n461_), .A3(new_n455_), .A4(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n462_), .A2(new_n447_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n433_), .A2(KEYINPUT98), .A3(new_n449_), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n433_), .A2(new_n449_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT98), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(KEYINPUT99), .B1(new_n476_), .B2(new_n479_), .ZN(new_n480_));
  AND4_X1   g279(.A1(KEYINPUT99), .A2(new_n479_), .A3(new_n474_), .A4(new_n475_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n473_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n427_), .ZN(new_n483_));
  OAI211_X1 g282(.A(KEYINPUT97), .B(KEYINPUT20), .C1(new_n427_), .C2(new_n464_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n467_), .A2(new_n470_), .A3(new_n483_), .A4(new_n484_), .ZN(new_n485_));
  AOI22_X1  g284(.A1(new_n417_), .A2(new_n410_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n476_), .A2(new_n479_), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n486_), .A2(new_n473_), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n464_), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT20), .B1(new_n486_), .B2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n469_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n485_), .A2(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(G8gat), .B(G36gat), .Z(new_n493_));
  XNOR2_X1  g292(.A(G64gat), .B(G92gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT32), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n492_), .A2(new_n500_), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n501_), .A2(KEYINPUT106), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n482_), .A2(new_n427_), .ZN(new_n503_));
  OAI211_X1 g302(.A(KEYINPUT20), .B(new_n470_), .C1(new_n486_), .C2(new_n489_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n467_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n505_), .B1(new_n506_), .B2(new_n469_), .ZN(new_n507_));
  AOI22_X1  g306(.A1(new_n501_), .A2(KEYINPUT106), .B1(new_n507_), .B2(new_n499_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n405_), .A2(new_n502_), .A3(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n403_), .A2(KEYINPUT33), .A3(new_n393_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT104), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT104), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n403_), .A2(new_n512_), .A3(new_n393_), .A4(KEYINPUT33), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n483_), .A2(new_n484_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n486_), .A2(new_n489_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT97), .B1(new_n516_), .B2(KEYINPUT20), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n469_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n505_), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n518_), .A2(new_n498_), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n498_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(KEYINPUT105), .B(KEYINPUT33), .Z(new_n523_));
  NAND2_X1  g322(.A1(new_n404_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n388_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n376_), .A2(new_n387_), .A3(new_n392_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n525_), .A2(new_n401_), .A3(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n522_), .A2(new_n524_), .A3(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n509_), .B1(new_n514_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT29), .ZN(new_n530_));
  OAI21_X1  g329(.A(KEYINPUT93), .B1(new_n384_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT93), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n368_), .A2(new_n532_), .A3(KEYINPUT29), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n531_), .A2(new_n533_), .A3(new_n427_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G228gat), .A2(G233gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT88), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n369_), .A2(KEYINPUT29), .A3(new_n371_), .ZN(new_n537_));
  XOR2_X1   g336(.A(new_n536_), .B(KEYINPUT89), .Z(new_n538_));
  NOR2_X1   g337(.A1(new_n486_), .A2(new_n538_), .ZN(new_n539_));
  AOI22_X1  g338(.A1(new_n534_), .A2(new_n536_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G78gat), .B(G106gat), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT95), .B1(new_n540_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT95), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n537_), .A2(new_n539_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n536_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n368_), .A2(KEYINPUT29), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n486_), .B1(new_n548_), .B2(KEYINPUT93), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n547_), .B1(new_n549_), .B2(new_n533_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n544_), .B(new_n541_), .C1(new_n546_), .C2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n540_), .A2(KEYINPUT96), .A3(new_n542_), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n543_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G22gat), .B(G50gat), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT28), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n369_), .A2(new_n371_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n556_), .B1(new_n557_), .B2(new_n530_), .ZN(new_n558_));
  AOI211_X1 g357(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n369_), .C2(new_n371_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n555_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n382_), .A2(new_n383_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n370_), .B1(new_n561_), .B2(new_n349_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n371_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n530_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT28), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n557_), .A2(new_n556_), .A3(new_n530_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n565_), .A2(new_n566_), .A3(new_n554_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n560_), .A2(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(KEYINPUT96), .B1(new_n540_), .B2(new_n542_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n553_), .A2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n541_), .B1(new_n546_), .B2(new_n550_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n540_), .A2(new_n542_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT94), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n574_), .A2(new_n575_), .A3(new_n568_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n575_), .B1(new_n574_), .B2(new_n568_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n571_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n529_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G71gat), .B(G99gat), .ZN(new_n581_));
  INV_X1    g380(.A(G43gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  AND2_X1   g382(.A1(G227gat), .A2(G233gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT30), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n464_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n450_), .A2(KEYINPUT30), .A3(new_n463_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT81), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n586_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n588_), .A2(KEYINPUT81), .A3(new_n589_), .A4(new_n585_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(KEYINPUT80), .B(G15gat), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n590_), .A2(new_n591_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n592_), .A2(new_n595_), .A3(new_n593_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n597_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT82), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT31), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT31), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n599_), .A2(new_n598_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n595_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n601_), .B(new_n604_), .C1(new_n605_), .C2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n603_), .A2(new_n375_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n607_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n604_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n374_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n608_), .A2(new_n611_), .ZN(new_n612_));
  AOI221_X4 g411(.A(new_n541_), .B1(new_n537_), .B2(new_n539_), .C1(new_n534_), .C2(new_n536_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n534_), .A2(new_n536_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n542_), .B1(new_n614_), .B2(new_n545_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n558_), .A2(new_n559_), .A3(new_n555_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n554_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n617_));
  OAI22_X1  g416(.A1(new_n613_), .A2(new_n615_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT94), .ZN(new_n619_));
  AOI22_X1  g418(.A1(new_n619_), .A2(new_n576_), .B1(new_n553_), .B2(new_n570_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT27), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n621_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n622_));
  AOI22_X1  g421(.A1(new_n395_), .A2(new_n401_), .B1(new_n393_), .B2(new_n403_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n507_), .A2(new_n498_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n492_), .A2(new_n497_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n624_), .A2(new_n625_), .A3(KEYINPUT27), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n622_), .A2(new_n623_), .A3(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n612_), .B1(new_n620_), .B2(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n328_), .B1(new_n580_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n627_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n579_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n511_), .A2(new_n513_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n632_), .A2(new_n524_), .A3(new_n522_), .A4(new_n527_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n620_), .A2(new_n633_), .A3(new_n509_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n631_), .A2(new_n634_), .A3(KEYINPUT107), .A4(new_n612_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n622_), .A2(new_n626_), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n636_), .A2(KEYINPUT108), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(KEYINPUT108), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n612_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n639_), .A2(new_n620_), .A3(new_n623_), .A4(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n629_), .A2(new_n635_), .A3(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n288_), .A2(new_n312_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT75), .ZN(new_n644_));
  NAND2_X1  g443(.A1(G229gat), .A2(G233gat), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n646_), .B1(new_n313_), .B2(new_n283_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n313_), .A2(new_n283_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n312_), .A2(new_n284_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  AOI22_X1  g449(.A1(new_n644_), .A2(new_n647_), .B1(new_n650_), .B2(new_n646_), .ZN(new_n651_));
  XOR2_X1   g450(.A(G113gat), .B(G141gat), .Z(new_n652_));
  XNOR2_X1  g451(.A(G169gat), .B(G197gat), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n651_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n651_), .A2(new_n654_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n642_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n327_), .A2(new_n658_), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n659_), .B(KEYINPUT109), .Z(new_n660_));
  NAND3_X1  g459(.A1(new_n660_), .A2(new_n307_), .A3(new_n405_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT38), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n657_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n325_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n272_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n298_), .A2(new_n301_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n642_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n666_), .A2(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G1gat), .B1(new_n670_), .B2(new_n623_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n661_), .A2(new_n662_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n663_), .A2(new_n671_), .A3(new_n672_), .ZN(G1324gat));
  INV_X1    g472(.A(new_n639_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n660_), .A2(new_n308_), .A3(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G8gat), .B1(new_n670_), .B2(new_n639_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n676_), .A2(KEYINPUT39), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(KEYINPUT39), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n675_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT40), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n675_), .B(KEYINPUT40), .C1(new_n677_), .C2(new_n678_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1325gat));
  OAI21_X1  g482(.A(G15gat), .B1(new_n670_), .B2(new_n612_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT41), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n659_), .A2(G15gat), .A3(new_n612_), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1326gat));
  OAI21_X1  g486(.A(G22gat), .B1(new_n670_), .B2(new_n620_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n688_), .A2(KEYINPUT42), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(KEYINPUT42), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n620_), .A2(G22gat), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT110), .ZN(new_n692_));
  OAI22_X1  g491(.A1(new_n689_), .A2(new_n690_), .B1(new_n659_), .B2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT111), .ZN(G1327gat));
  NAND2_X1  g493(.A1(new_n667_), .A2(new_n665_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n272_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(new_n658_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G29gat), .B1(new_n698_), .B2(new_n405_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n701_));
  INV_X1    g500(.A(new_n305_), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n642_), .A2(new_n701_), .A3(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n701_), .B1(new_n642_), .B2(new_n702_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n272_), .A2(new_n664_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(new_n665_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n700_), .B1(new_n705_), .B2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n642_), .A2(new_n702_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT43), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n642_), .A2(new_n701_), .A3(new_n702_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n712_), .A2(KEYINPUT44), .A3(new_n665_), .A4(new_n706_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n708_), .A2(new_n713_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n405_), .A2(G29gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n699_), .B1(new_n714_), .B2(new_n715_), .ZN(G1328gat));
  NOR3_X1   g515(.A1(new_n697_), .A2(G36gat), .A3(new_n639_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT45), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n717_), .B(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n708_), .A2(new_n713_), .A3(new_n674_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(G36gat), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT46), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n722_), .B(new_n723_), .ZN(G1329gat));
  NAND4_X1  g523(.A1(new_n708_), .A2(new_n713_), .A3(G43gat), .A4(new_n640_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n582_), .B1(new_n697_), .B2(new_n612_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g527(.A1(new_n697_), .A2(G50gat), .A3(new_n620_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n714_), .A2(new_n579_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n730_), .A2(KEYINPUT112), .ZN(new_n731_));
  OAI21_X1  g530(.A(G50gat), .B1(new_n730_), .B2(KEYINPUT112), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n729_), .B1(new_n731_), .B2(new_n732_), .ZN(G1331gat));
  NAND4_X1  g532(.A1(new_n669_), .A2(new_n664_), .A3(new_n272_), .A4(new_n325_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n405_), .A2(G57gat), .ZN(new_n735_));
  OR3_X1    g534(.A1(new_n734_), .A2(KEYINPUT113), .A3(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(KEYINPUT113), .B1(new_n734_), .B2(new_n735_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n642_), .A2(new_n664_), .ZN(new_n738_));
  AND4_X1   g537(.A1(new_n272_), .A2(new_n738_), .A3(new_n325_), .A4(new_n305_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n740_), .A2(new_n623_), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n736_), .B(new_n737_), .C1(new_n741_), .C2(G57gat), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT114), .Z(G1332gat));
  OAI21_X1  g542(.A(G64gat), .B1(new_n734_), .B2(new_n639_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT48), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n639_), .A2(G64gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n740_), .B2(new_n746_), .ZN(G1333gat));
  OAI21_X1  g546(.A(G71gat), .B1(new_n734_), .B2(new_n612_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT49), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n612_), .A2(G71gat), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n749_), .B1(new_n740_), .B2(new_n750_), .ZN(G1334gat));
  OAI21_X1  g550(.A(G78gat), .B1(new_n734_), .B2(new_n620_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT50), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n620_), .A2(G78gat), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n753_), .B1(new_n740_), .B2(new_n754_), .ZN(G1335gat));
  NOR2_X1   g554(.A1(new_n657_), .A2(new_n325_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n272_), .A2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n757_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(G85gat), .B1(new_n759_), .B2(new_n623_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n738_), .A2(new_n272_), .A3(new_n665_), .A4(new_n667_), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n623_), .A2(G85gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n760_), .B1(new_n761_), .B2(new_n762_), .ZN(G1336gat));
  OAI21_X1  g562(.A(G92gat), .B1(new_n759_), .B2(new_n639_), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n639_), .A2(G92gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n761_), .B2(new_n765_), .ZN(G1337gat));
  OR3_X1    g565(.A1(new_n761_), .A2(new_n612_), .A3(new_n219_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n758_), .A2(new_n640_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n768_), .A2(KEYINPUT115), .A3(G99gat), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT115), .B1(new_n768_), .B2(G99gat), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n767_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT51), .ZN(G1338gat));
  AOI211_X1 g571(.A(new_n657_), .B(new_n325_), .C1(new_n270_), .C2(new_n271_), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n773_), .B(new_n579_), .C1(new_n703_), .C2(new_n704_), .ZN(new_n774_));
  OAI21_X1  g573(.A(G106gat), .B1(new_n774_), .B2(KEYINPUT116), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n776_), .B1(new_n758_), .B2(new_n579_), .ZN(new_n777_));
  OAI21_X1  g576(.A(KEYINPUT52), .B1(new_n775_), .B2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n758_), .A2(new_n776_), .A3(new_n579_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n774_), .A2(KEYINPUT116), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n779_), .A2(new_n780_), .A3(new_n781_), .A4(G106gat), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n778_), .A2(new_n782_), .ZN(new_n783_));
  OR3_X1    g582(.A1(new_n761_), .A2(new_n620_), .A3(new_n220_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT53), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n783_), .A2(new_n787_), .A3(new_n784_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(G1339gat));
  NOR4_X1   g588(.A1(new_n674_), .A2(new_n579_), .A3(new_n623_), .A4(new_n612_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT118), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n644_), .A2(new_n648_), .A3(new_n646_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n654_), .B1(new_n650_), .B2(new_n645_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n656_), .A2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n265_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n246_), .A2(new_n799_), .A3(new_n255_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n253_), .A2(new_n254_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n247_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n802_));
  AOI22_X1  g601(.A1(new_n801_), .A2(KEYINPUT55), .B1(new_n250_), .B2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n261_), .B1(new_n800_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT56), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT117), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n657_), .B(new_n264_), .C1(new_n804_), .C2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n804_), .A2(KEYINPUT117), .A3(new_n805_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n798_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n792_), .B1(new_n811_), .B2(new_n667_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT58), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n804_), .A2(new_n805_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n264_), .A2(new_n796_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n804_), .A2(new_n805_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n813_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n817_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n819_), .A2(KEYINPUT58), .A3(new_n814_), .A4(new_n815_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n818_), .A2(new_n820_), .A3(new_n702_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n810_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n797_), .B1(new_n822_), .B2(new_n808_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n823_), .A2(KEYINPUT57), .A3(new_n668_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n812_), .A2(new_n821_), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n665_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n266_), .A2(new_n268_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n664_), .A2(new_n325_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n828_), .B1(new_n302_), .B2(new_n304_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n827_), .A2(new_n829_), .A3(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n830_), .B1(new_n827_), .B2(new_n829_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n791_), .B1(new_n826_), .B2(new_n835_), .ZN(new_n836_));
  AOI211_X1 g635(.A(KEYINPUT118), .B(new_n834_), .C1(new_n825_), .C2(new_n665_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n657_), .B(new_n790_), .C1(new_n836_), .C2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(G113gat), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT119), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n838_), .A2(KEYINPUT119), .A3(new_n839_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n790_), .A2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n845_), .B1(new_n826_), .B2(new_n835_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n790_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n847_), .B2(KEYINPUT59), .ZN(new_n848_));
  XOR2_X1   g647(.A(KEYINPUT121), .B(G113gat), .Z(new_n849_));
  NOR2_X1   g648(.A1(new_n664_), .A2(new_n849_), .ZN(new_n850_));
  AOI22_X1  g649(.A1(new_n842_), .A2(new_n843_), .B1(new_n848_), .B2(new_n850_), .ZN(G1340gat));
  INV_X1    g650(.A(new_n272_), .ZN(new_n852_));
  AOI211_X1 g651(.A(new_n852_), .B(new_n846_), .C1(new_n847_), .C2(KEYINPUT59), .ZN(new_n853_));
  INV_X1    g652(.A(G120gat), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT60), .ZN(new_n855_));
  AOI21_X1  g654(.A(G120gat), .B1(new_n272_), .B2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(KEYINPUT122), .B1(new_n855_), .B2(G120gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n856_), .B2(new_n859_), .ZN(new_n860_));
  OAI22_X1  g659(.A1(new_n853_), .A2(new_n854_), .B1(new_n847_), .B2(new_n860_), .ZN(G1341gat));
  AOI211_X1 g660(.A(new_n665_), .B(new_n846_), .C1(new_n847_), .C2(KEYINPUT59), .ZN(new_n862_));
  INV_X1    g661(.A(G127gat), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n325_), .A2(new_n863_), .ZN(new_n864_));
  OAI22_X1  g663(.A1(new_n862_), .A2(new_n863_), .B1(new_n847_), .B2(new_n864_), .ZN(G1342gat));
  AOI211_X1 g664(.A(new_n305_), .B(new_n846_), .C1(new_n847_), .C2(KEYINPUT59), .ZN(new_n866_));
  INV_X1    g665(.A(G134gat), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n667_), .A2(new_n867_), .ZN(new_n868_));
  OAI22_X1  g667(.A1(new_n866_), .A2(new_n867_), .B1(new_n847_), .B2(new_n868_), .ZN(G1343gat));
  OR2_X1    g668(.A1(new_n836_), .A2(new_n837_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n640_), .A2(new_n620_), .ZN(new_n871_));
  AND3_X1   g670(.A1(new_n871_), .A2(new_n405_), .A3(new_n639_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n870_), .A2(new_n657_), .A3(new_n872_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g673(.A1(new_n870_), .A2(new_n272_), .A3(new_n872_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g675(.A1(new_n870_), .A2(new_n325_), .A3(new_n872_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(KEYINPUT61), .B(G155gat), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1346gat));
  NOR2_X1   g678(.A1(new_n305_), .A2(new_n361_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n870_), .A2(new_n872_), .A3(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT123), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n667_), .B(new_n872_), .C1(new_n836_), .C2(new_n837_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n883_), .B1(new_n885_), .B2(G162gat), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n884_), .A2(KEYINPUT123), .A3(new_n361_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n882_), .B1(new_n886_), .B2(new_n887_), .ZN(G1347gat));
  NOR2_X1   g687(.A1(new_n639_), .A2(new_n405_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n640_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(KEYINPUT124), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n657_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(KEYINPUT125), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n579_), .B1(new_n826_), .B2(new_n835_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n428_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT62), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n895_), .A2(new_n896_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n894_), .A2(new_n891_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n657_), .A2(new_n436_), .ZN(new_n900_));
  OAI22_X1  g699(.A1(new_n897_), .A2(new_n898_), .B1(new_n899_), .B2(new_n900_), .ZN(G1348gat));
  AND2_X1   g700(.A1(new_n870_), .A2(new_n620_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n891_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n903_), .A2(new_n432_), .A3(new_n852_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n894_), .A2(new_n272_), .A3(new_n891_), .ZN(new_n905_));
  AOI22_X1  g704(.A1(new_n902_), .A2(new_n904_), .B1(new_n432_), .B2(new_n905_), .ZN(G1349gat));
  NAND4_X1  g705(.A1(new_n870_), .A2(new_n620_), .A3(new_n325_), .A4(new_n891_), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n903_), .A2(new_n456_), .A3(new_n665_), .ZN(new_n908_));
  AOI22_X1  g707(.A1(new_n907_), .A2(new_n439_), .B1(new_n894_), .B2(new_n908_), .ZN(G1350gat));
  OAI21_X1  g708(.A(G190gat), .B1(new_n899_), .B2(new_n305_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n667_), .A2(new_n459_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n899_), .B2(new_n911_), .ZN(G1351gat));
  AND2_X1   g711(.A1(new_n889_), .A2(new_n871_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n870_), .A2(new_n657_), .A3(new_n913_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G197gat), .ZN(G1352gat));
  OAI211_X1 g714(.A(new_n272_), .B(new_n913_), .C1(new_n836_), .C2(new_n837_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(new_n414_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n917_), .B1(new_n419_), .B2(new_n916_), .ZN(G1353gat));
  AOI21_X1  g717(.A(new_n665_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n870_), .A2(new_n913_), .A3(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(KEYINPUT126), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n920_), .B(new_n923_), .ZN(G1354gat));
  AND2_X1   g723(.A1(new_n702_), .A2(G218gat), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n870_), .A2(new_n913_), .A3(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  OAI211_X1 g726(.A(new_n667_), .B(new_n913_), .C1(new_n836_), .C2(new_n837_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(G218gat), .B1(new_n929_), .B2(KEYINPUT127), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n928_), .A2(new_n931_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n927_), .B1(new_n930_), .B2(new_n932_), .ZN(G1355gat));
endmodule


