//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n606_, new_n607_, new_n608_, new_n609_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n616_, new_n617_, new_n618_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n816_, new_n817_, new_n818_, new_n820_,
    new_n821_, new_n822_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n834_,
    new_n835_, new_n836_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n870_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n894_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(G15gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT30), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G169gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n207_), .A2(KEYINPUT22), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT86), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n207_), .A2(KEYINPUT22), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT85), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT87), .B(G176gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n210_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT88), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n218_), .B(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT89), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n219_), .A2(KEYINPUT89), .A3(G183gat), .A4(G190gat), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  OR2_X1    g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225_));
  AOI22_X1  g024(.A1(new_n224_), .A2(new_n225_), .B1(G169gat), .B2(G176gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n217_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(G176gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT24), .B1(new_n207_), .B2(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT25), .B(G183gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT26), .B(G190gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT24), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n230_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n220_), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n231_), .A2(new_n234_), .A3(new_n236_), .A4(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n227_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G71gat), .B(G99gat), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n240_), .B(G43gat), .Z(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n239_), .A2(new_n241_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n206_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n244_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n246_), .A2(new_n205_), .A3(new_n242_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(G127gat), .B(G134gat), .Z(new_n249_));
  XOR2_X1   g048(.A(G113gat), .B(G120gat), .Z(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT90), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT31), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT91), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n248_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT92), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n256_), .B1(new_n247_), .B2(new_n245_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT92), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n245_), .A2(new_n247_), .A3(new_n254_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n260_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT93), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT93), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n260_), .A2(new_n262_), .A3(new_n266_), .A4(new_n263_), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G225gat), .A2(G233gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT103), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n271_));
  NOR2_X1   g070(.A1(G155gat), .A2(G162gat), .ZN(new_n272_));
  INV_X1    g071(.A(G155gat), .ZN(new_n273_));
  INV_X1    g072(.A(G162gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(G141gat), .A2(G148gat), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT3), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G141gat), .A2(G148gat), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT2), .ZN(new_n279_));
  OAI22_X1  g078(.A1(new_n276_), .A2(new_n277_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n280_), .B1(new_n277_), .B2(new_n276_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n278_), .A2(new_n279_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT94), .ZN(new_n283_));
  AOI211_X1 g082(.A(new_n272_), .B(new_n275_), .C1(new_n281_), .C2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n278_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT1), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n272_), .B1(new_n275_), .B2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(KEYINPUT1), .B1(new_n273_), .B2(new_n274_), .ZN(new_n288_));
  AOI211_X1 g087(.A(new_n285_), .B(new_n276_), .C1(new_n287_), .C2(new_n288_), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n284_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(new_n253_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n251_), .ZN(new_n292_));
  OR3_X1    g091(.A1(new_n284_), .A2(new_n292_), .A3(new_n289_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n271_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT4), .B1(new_n290_), .B2(new_n253_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n270_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n291_), .A2(new_n293_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n269_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G1gat), .B(G29gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(G85gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT0), .B(G57gat), .ZN(new_n302_));
  XOR2_X1   g101(.A(new_n301_), .B(new_n302_), .Z(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n299_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n296_), .A2(new_n298_), .A3(new_n303_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(KEYINPUT95), .A2(G233gat), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(KEYINPUT95), .A2(G233gat), .ZN(new_n310_));
  OAI21_X1  g109(.A(G228gat), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n290_), .A2(KEYINPUT29), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT96), .B(G204gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(G197gat), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n315_), .B1(G197gat), .B2(G204gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G211gat), .B(G218gat), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT21), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT21), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n321_), .B1(G197gat), .B2(G204gat), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n322_), .B1(new_n314_), .B2(G197gat), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n323_), .B(KEYINPUT97), .Z(new_n324_));
  AOI21_X1  g123(.A(new_n318_), .B1(new_n316_), .B2(new_n321_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n320_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n312_), .B1(new_n313_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n290_), .A2(KEYINPUT29), .ZN(new_n328_));
  INV_X1    g127(.A(new_n326_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n328_), .A2(new_n329_), .A3(new_n311_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n327_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G78gat), .B(G106gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n332_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n327_), .A2(new_n330_), .A3(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n290_), .A2(KEYINPUT29), .ZN(new_n337_));
  XOR2_X1   g136(.A(G22gat), .B(G50gat), .Z(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT28), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n337_), .B(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n334_), .B1(new_n327_), .B2(new_n330_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n340_), .B1(new_n341_), .B2(KEYINPUT98), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n336_), .A2(new_n342_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n333_), .A2(KEYINPUT98), .A3(new_n335_), .A4(new_n340_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n307_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G226gat), .A2(G233gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT19), .ZN(new_n347_));
  AND4_X1   g146(.A1(new_n223_), .A2(new_n222_), .A3(new_n234_), .A4(new_n236_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n230_), .B1(new_n229_), .B2(KEYINPUT99), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n349_), .B1(KEYINPUT99), .B2(new_n229_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT22), .B(G169gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT100), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(new_n214_), .ZN(new_n353_));
  AOI22_X1  g152(.A1(new_n237_), .A2(new_n225_), .B1(G169gat), .B2(G176gat), .ZN(new_n354_));
  AOI22_X1  g153(.A1(new_n348_), .A2(new_n350_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n326_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT20), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n239_), .A2(new_n329_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n347_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n347_), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n326_), .A2(KEYINPUT101), .A3(new_n355_), .ZN(new_n361_));
  AOI21_X1  g160(.A(KEYINPUT101), .B1(new_n326_), .B2(new_n355_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n360_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n239_), .A2(new_n329_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT20), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n359_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  XOR2_X1   g165(.A(G8gat), .B(G36gat), .Z(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT102), .B(KEYINPUT18), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G64gat), .B(G92gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n366_), .A2(new_n371_), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n365_), .A2(new_n363_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n371_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(new_n359_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n372_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT27), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n326_), .A2(new_n355_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n347_), .B1(new_n365_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n358_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n381_), .A2(new_n356_), .A3(KEYINPUT20), .A4(new_n360_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(new_n371_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(KEYINPUT27), .A3(new_n375_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n345_), .A2(new_n378_), .A3(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n343_), .A2(new_n344_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n374_), .A2(KEYINPUT32), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n383_), .A2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n373_), .A2(new_n359_), .A3(new_n388_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n307_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT33), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n269_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n303_), .B1(new_n297_), .B2(new_n270_), .ZN(new_n395_));
  AOI22_X1  g194(.A1(new_n306_), .A2(new_n393_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n296_), .A2(new_n298_), .A3(KEYINPUT33), .A4(new_n303_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n396_), .A2(new_n372_), .A3(new_n375_), .A4(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n387_), .B1(new_n392_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT104), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n386_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  AOI211_X1 g200(.A(KEYINPUT104), .B(new_n387_), .C1(new_n398_), .C2(new_n392_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n268_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT105), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  OAI211_X1 g204(.A(KEYINPUT105), .B(new_n268_), .C1(new_n401_), .C2(new_n402_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n268_), .A2(new_n307_), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n378_), .A2(new_n385_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n409_), .A2(new_n387_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n407_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n405_), .A2(new_n406_), .A3(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT79), .B(G15gat), .ZN(new_n413_));
  INV_X1    g212(.A(G22gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT14), .ZN(new_n416_));
  XOR2_X1   g215(.A(KEYINPUT81), .B(G8gat), .Z(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT80), .B(G1gat), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n416_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n415_), .A2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G1gat), .B(G8gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G29gat), .B(G36gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G43gat), .B(G50gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(new_n425_), .B(KEYINPUT15), .Z(new_n426_));
  NOR2_X1   g225(.A1(new_n422_), .A2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT84), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n422_), .A2(new_n425_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G229gat), .A2(G233gat), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n422_), .B(new_n425_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n430_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n431_), .A2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G113gat), .B(G141gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G169gat), .B(G197gat), .ZN(new_n437_));
  XOR2_X1   g236(.A(new_n436_), .B(new_n437_), .Z(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n435_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n431_), .A2(new_n434_), .A3(new_n438_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n412_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT13), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G230gat), .A2(G233gat), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  AND3_X1   g245(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  XOR2_X1   g248(.A(KEYINPUT10), .B(G99gat), .Z(new_n450_));
  INV_X1    g249(.A(G106gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  XOR2_X1   g251(.A(G85gat), .B(G92gat), .Z(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT9), .ZN(new_n454_));
  INV_X1    g253(.A(G85gat), .ZN(new_n455_));
  INV_X1    g254(.A(G92gat), .ZN(new_n456_));
  OR3_X1    g255(.A1(new_n455_), .A2(new_n456_), .A3(KEYINPUT9), .ZN(new_n457_));
  AND4_X1   g256(.A1(new_n449_), .A2(new_n452_), .A3(new_n454_), .A4(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NOR3_X1   g259(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G99gat), .A2(G106gat), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT6), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT64), .ZN(new_n466_));
  NAND3_X1  g265(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT64), .B1(new_n447_), .B2(new_n448_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n462_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n453_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT65), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n470_), .A2(KEYINPUT65), .A3(new_n453_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(KEYINPUT8), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n462_), .A2(new_n449_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT8), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n476_), .A2(new_n477_), .A3(new_n453_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n458_), .B1(new_n475_), .B2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G57gat), .B(G64gat), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n480_), .A2(KEYINPUT11), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G71gat), .B(G78gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n481_), .A2(new_n482_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n480_), .A2(KEYINPUT11), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n483_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n479_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT66), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n479_), .A2(new_n486_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n446_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT67), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT67), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n492_), .B(new_n446_), .C1(new_n488_), .C2(new_n489_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  OAI211_X1 g293(.A(KEYINPUT12), .B(new_n483_), .C1(new_n484_), .C2(new_n485_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT69), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT68), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n470_), .A2(KEYINPUT65), .A3(new_n453_), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT65), .B1(new_n470_), .B2(new_n453_), .ZN(new_n500_));
  NOR3_X1   g299(.A1(new_n499_), .A2(new_n500_), .A3(new_n477_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n478_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n498_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n475_), .A2(KEYINPUT68), .A3(new_n478_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n458_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n497_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  AOI211_X1 g306(.A(KEYINPUT69), .B(new_n458_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n496_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(KEYINPUT70), .B(KEYINPUT12), .Z(new_n510_));
  OAI21_X1  g309(.A(new_n510_), .B1(new_n479_), .B2(new_n486_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT71), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  OAI211_X1 g312(.A(KEYINPUT71), .B(new_n510_), .C1(new_n479_), .C2(new_n486_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n446_), .B1(new_n479_), .B2(new_n486_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n509_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  XOR2_X1   g316(.A(G120gat), .B(G148gat), .Z(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G176gat), .B(G204gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n494_), .A2(new_n517_), .A3(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n523_), .B1(new_n494_), .B2(new_n517_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n444_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n494_), .A2(new_n517_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n522_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n494_), .A2(new_n517_), .A3(new_n523_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n528_), .A2(KEYINPUT13), .A3(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G231gat), .A2(G233gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT82), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n422_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(new_n486_), .ZN(new_n534_));
  XOR2_X1   g333(.A(G127gat), .B(G155gat), .Z(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT16), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G183gat), .B(G211gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT17), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n538_), .A2(new_n539_), .ZN(new_n541_));
  NOR3_X1   g340(.A1(new_n534_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(KEYINPUT83), .B1(new_n534_), .B2(new_n541_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NOR4_X1   g343(.A1(new_n534_), .A2(KEYINPUT83), .A3(new_n540_), .A4(new_n541_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n526_), .A2(new_n530_), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT78), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT37), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(KEYINPUT78), .A2(KEYINPUT37), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT36), .ZN(new_n552_));
  INV_X1    g351(.A(new_n426_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n553_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT74), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n479_), .A2(new_n425_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT73), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n479_), .A2(KEYINPUT73), .A3(new_n425_), .ZN(new_n559_));
  AOI21_X1  g358(.A(KEYINPUT77), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n554_), .A2(new_n555_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G232gat), .A2(G233gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT34), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT35), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n561_), .A2(new_n565_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n554_), .A2(new_n555_), .A3(new_n560_), .A4(new_n564_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n554_), .A2(new_n560_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT35), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n566_), .A2(new_n567_), .A3(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G190gat), .B(G218gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT75), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G134gat), .B(G162gat), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n573_), .B(new_n574_), .Z(new_n575_));
  NAND2_X1  g374(.A1(new_n571_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT76), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n571_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n575_), .ZN(new_n579_));
  AOI22_X1  g378(.A1(new_n552_), .A2(new_n576_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  AOI211_X1 g379(.A(KEYINPUT36), .B(new_n575_), .C1(new_n571_), .C2(new_n577_), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n550_), .B(new_n551_), .C1(new_n580_), .C2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n578_), .A2(new_n579_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n576_), .A2(new_n552_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n578_), .A2(new_n552_), .A3(new_n579_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n585_), .A2(new_n548_), .A3(new_n549_), .A4(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n582_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n443_), .A2(new_n547_), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n307_), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n590_), .A2(new_n591_), .A3(new_n418_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n592_), .A2(KEYINPUT38), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(KEYINPUT38), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n585_), .A2(new_n586_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n526_), .A2(new_n530_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n442_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n546_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n597_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n412_), .A2(new_n596_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(G1gat), .B1(new_n602_), .B2(new_n591_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n593_), .A2(new_n594_), .A3(new_n603_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT106), .Z(G1324gat));
  OAI21_X1  g404(.A(G8gat), .B1(new_n602_), .B2(new_n408_), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n606_), .B(KEYINPUT39), .Z(new_n607_));
  NOR3_X1   g406(.A1(new_n590_), .A2(new_n408_), .A3(new_n417_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT40), .ZN(G1325gat));
  INV_X1    g409(.A(new_n268_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n203_), .B1(new_n601_), .B2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT41), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n203_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n613_), .B1(new_n590_), .B2(new_n614_), .ZN(G1326gat));
  AOI21_X1  g414(.A(new_n414_), .B1(new_n601_), .B2(new_n387_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT42), .Z(new_n617_));
  NAND2_X1  g416(.A1(new_n387_), .A2(new_n414_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n617_), .B1(new_n590_), .B2(new_n618_), .ZN(G1327gat));
  INV_X1    g418(.A(new_n597_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n596_), .A2(new_n546_), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n443_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(G29gat), .B1(new_n622_), .B2(new_n307_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT43), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n412_), .A2(new_n624_), .A3(new_n588_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n624_), .B1(new_n412_), .B2(new_n588_), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n597_), .A2(new_n598_), .A3(new_n546_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(KEYINPUT44), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n630_), .A2(G29gat), .A3(new_n307_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n629_), .A2(KEYINPUT44), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n623_), .B1(new_n631_), .B2(new_n633_), .ZN(G1328gat));
  NAND2_X1  g433(.A1(new_n630_), .A2(new_n409_), .ZN(new_n635_));
  OAI21_X1  g434(.A(G36gat), .B1(new_n635_), .B2(new_n632_), .ZN(new_n636_));
  INV_X1    g435(.A(G36gat), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n622_), .A2(new_n637_), .A3(new_n409_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT45), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n636_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT46), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n636_), .A2(KEYINPUT46), .A3(new_n639_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(G1329gat));
  AOI21_X1  g443(.A(G43gat), .B1(new_n622_), .B2(new_n611_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT107), .Z(new_n646_));
  NAND3_X1  g445(.A1(new_n630_), .A2(G43gat), .A3(new_n611_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n646_), .B1(new_n647_), .B2(new_n632_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g448(.A(G50gat), .B1(new_n622_), .B2(new_n387_), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n630_), .A2(G50gat), .A3(new_n387_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n651_), .B2(new_n633_), .ZN(G1331gat));
  INV_X1    g451(.A(G57gat), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n412_), .A2(new_n598_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n654_), .A2(new_n597_), .A3(new_n546_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(new_n589_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n653_), .B1(new_n656_), .B2(new_n591_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n596_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n658_), .A2(new_n653_), .A3(new_n591_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n657_), .B1(new_n659_), .B2(KEYINPUT108), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n660_), .B1(KEYINPUT108), .B2(new_n659_), .ZN(G1332gat));
  OAI21_X1  g460(.A(G64gat), .B1(new_n658_), .B2(new_n408_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT48), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n408_), .A2(G64gat), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n663_), .B1(new_n656_), .B2(new_n664_), .ZN(G1333gat));
  OAI21_X1  g464(.A(G71gat), .B1(new_n658_), .B2(new_n268_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT49), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n268_), .A2(G71gat), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT109), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n667_), .B1(new_n656_), .B2(new_n669_), .ZN(G1334gat));
  INV_X1    g469(.A(new_n387_), .ZN(new_n671_));
  OAI21_X1  g470(.A(G78gat), .B1(new_n658_), .B2(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT50), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n671_), .A2(G78gat), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n673_), .B1(new_n656_), .B2(new_n674_), .ZN(G1335gat));
  NAND3_X1  g474(.A1(new_n654_), .A2(new_n597_), .A3(new_n621_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n455_), .B1(new_n676_), .B2(new_n591_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT110), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n620_), .A2(new_n442_), .A3(new_n546_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n627_), .A2(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n591_), .A2(new_n455_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n678_), .B1(new_n680_), .B2(new_n681_), .ZN(G1336gat));
  NOR3_X1   g481(.A1(new_n676_), .A2(G92gat), .A3(new_n408_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n680_), .A2(new_n409_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n684_), .B2(G92gat), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT111), .ZN(G1337gat));
  NAND2_X1  g485(.A1(new_n611_), .A2(new_n450_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n676_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n680_), .A2(new_n611_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(G99gat), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT51), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n691_), .A2(KEYINPUT112), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n690_), .B(new_n692_), .Z(G1338gat));
  OAI211_X1 g492(.A(new_n387_), .B(new_n679_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT113), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n451_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT114), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n696_), .A2(KEYINPUT114), .A3(new_n697_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n700_), .A2(KEYINPUT52), .A3(new_n701_), .ZN(new_n702_));
  OR3_X1    g501(.A1(new_n676_), .A2(G106gat), .A3(new_n671_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT52), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n698_), .A2(new_n699_), .A3(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n702_), .A2(new_n703_), .A3(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT53), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT53), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n702_), .A2(new_n708_), .A3(new_n703_), .A4(new_n705_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(G1339gat));
  NAND3_X1  g509(.A1(new_n428_), .A2(new_n429_), .A3(new_n433_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n438_), .B1(new_n432_), .B2(new_n430_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n441_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n524_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n488_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n509_), .A2(new_n718_), .A3(new_n515_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n517_), .A2(KEYINPUT55), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT55), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n509_), .A2(new_n515_), .A3(new_n721_), .A4(new_n516_), .ZN(new_n722_));
  AOI221_X4 g521(.A(KEYINPUT116), .B1(new_n719_), .B2(new_n446_), .C1(new_n720_), .C2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT116), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n720_), .A2(new_n722_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n719_), .A2(new_n446_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n724_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n522_), .B1(new_n723_), .B2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT56), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n477_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n731_));
  AOI211_X1 g530(.A(new_n498_), .B(new_n502_), .C1(new_n731_), .C2(new_n474_), .ZN(new_n732_));
  AOI21_X1  g531(.A(KEYINPUT68), .B1(new_n475_), .B2(new_n478_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n506_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT69), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n505_), .A2(new_n497_), .A3(new_n506_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  AOI22_X1  g536(.A1(new_n737_), .A2(new_n496_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n721_), .B1(new_n738_), .B2(new_n516_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n722_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n726_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT116), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n725_), .A2(new_n724_), .A3(new_n726_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n744_), .A2(KEYINPUT56), .A3(new_n522_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n717_), .B1(new_n730_), .B2(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(KEYINPUT58), .B1(new_n746_), .B2(KEYINPUT117), .ZN(new_n747_));
  AOI21_X1  g546(.A(KEYINPUT56), .B1(new_n744_), .B2(new_n522_), .ZN(new_n748_));
  AOI211_X1 g547(.A(new_n729_), .B(new_n523_), .C1(new_n742_), .C2(new_n743_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n716_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT117), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT58), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n750_), .A2(new_n751_), .A3(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n747_), .A2(new_n753_), .A3(new_n588_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT115), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n755_), .B1(new_n524_), .B2(new_n598_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n529_), .A2(KEYINPUT115), .A3(new_n442_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n730_), .B2(new_n745_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n715_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n596_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT57), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n756_), .A2(new_n757_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n764_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n760_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n767_), .A2(KEYINPUT57), .A3(new_n596_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n754_), .A2(new_n763_), .A3(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n599_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n582_), .A2(new_n587_), .A3(new_n598_), .A4(new_n547_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT54), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n771_), .B(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n770_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n611_), .A2(new_n410_), .A3(new_n307_), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n776_), .A2(KEYINPUT121), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT59), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(KEYINPUT121), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n777_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n775_), .A2(KEYINPUT122), .A3(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT122), .B1(new_n775_), .B2(new_n781_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT120), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT57), .B1(new_n767_), .B2(new_n596_), .ZN(new_n786_));
  AOI211_X1 g585(.A(new_n762_), .B(new_n595_), .C1(new_n765_), .C2(new_n766_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n546_), .B1(new_n788_), .B2(new_n754_), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT118), .B1(new_n789_), .B2(new_n773_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT118), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n770_), .A2(new_n791_), .A3(new_n774_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n776_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n785_), .B1(new_n793_), .B2(new_n778_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n776_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n791_), .B1(new_n770_), .B2(new_n774_), .ZN(new_n796_));
  AOI211_X1 g595(.A(KEYINPUT118), .B(new_n773_), .C1(new_n769_), .C2(new_n599_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n795_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(KEYINPUT120), .A3(KEYINPUT59), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n784_), .B1(new_n794_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(G113gat), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n598_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n793_), .A2(KEYINPUT119), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n798_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n803_), .A2(new_n442_), .A3(new_n805_), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n800_), .A2(new_n802_), .B1(new_n806_), .B2(new_n801_), .ZN(G1340gat));
  INV_X1    g606(.A(KEYINPUT60), .ZN(new_n808_));
  AOI21_X1  g607(.A(G120gat), .B1(new_n597_), .B2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n809_), .B1(new_n808_), .B2(G120gat), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n803_), .A2(new_n805_), .A3(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n597_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(new_n794_), .B2(new_n799_), .ZN(new_n813_));
  INV_X1    g612(.A(G120gat), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n811_), .B1(new_n813_), .B2(new_n814_), .ZN(G1341gat));
  INV_X1    g614(.A(G127gat), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n599_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n803_), .A2(new_n546_), .A3(new_n805_), .ZN(new_n818_));
  AOI22_X1  g617(.A1(new_n800_), .A2(new_n817_), .B1(new_n818_), .B2(new_n816_), .ZN(G1342gat));
  INV_X1    g618(.A(G134gat), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n589_), .A2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n803_), .A2(new_n595_), .A3(new_n805_), .ZN(new_n822_));
  AOI22_X1  g621(.A1(new_n800_), .A2(new_n821_), .B1(new_n822_), .B2(new_n820_), .ZN(G1343gat));
  NAND2_X1  g622(.A1(new_n790_), .A2(new_n792_), .ZN(new_n824_));
  NOR4_X1   g623(.A1(new_n611_), .A2(new_n671_), .A3(new_n591_), .A4(new_n409_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT123), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  OAI211_X1 g625(.A(KEYINPUT123), .B(new_n825_), .C1(new_n796_), .C2(new_n797_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(G141gat), .B1(new_n829_), .B2(new_n598_), .ZN(new_n830_));
  INV_X1    g629(.A(G141gat), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n831_), .B(new_n442_), .C1(new_n826_), .C2(new_n828_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1344gat));
  OAI21_X1  g632(.A(G148gat), .B1(new_n829_), .B2(new_n620_), .ZN(new_n834_));
  INV_X1    g633(.A(G148gat), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n835_), .B(new_n597_), .C1(new_n826_), .C2(new_n828_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(G1345gat));
  XNOR2_X1  g636(.A(KEYINPUT61), .B(G155gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n829_), .B2(new_n599_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n838_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n546_), .B(new_n840_), .C1(new_n826_), .C2(new_n828_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n841_), .ZN(G1346gat));
  OAI21_X1  g641(.A(G162gat), .B1(new_n829_), .B2(new_n589_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n274_), .B(new_n595_), .C1(new_n826_), .C2(new_n828_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(G1347gat));
  AOI21_X1  g644(.A(new_n387_), .B1(new_n770_), .B2(new_n774_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n407_), .A2(new_n409_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n207_), .B1(new_n850_), .B2(new_n442_), .ZN(new_n851_));
  OR2_X1    g650(.A1(new_n851_), .A2(KEYINPUT62), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n442_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n853_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n854_));
  INV_X1    g653(.A(new_n352_), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n852_), .B(new_n854_), .C1(new_n855_), .C2(new_n853_), .ZN(G1348gat));
  NAND2_X1  g655(.A1(new_n850_), .A2(new_n597_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n387_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n847_), .A2(new_n228_), .A3(new_n620_), .ZN(new_n859_));
  AOI22_X1  g658(.A1(new_n857_), .A2(new_n214_), .B1(new_n858_), .B2(new_n859_), .ZN(G1349gat));
  NOR2_X1   g659(.A1(new_n847_), .A2(new_n599_), .ZN(new_n861_));
  AOI21_X1  g660(.A(G183gat), .B1(new_n858_), .B2(new_n861_), .ZN(new_n862_));
  NOR3_X1   g661(.A1(new_n847_), .A2(new_n232_), .A3(new_n599_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n862_), .B1(new_n846_), .B2(new_n863_), .ZN(G1350gat));
  OAI21_X1  g663(.A(G190gat), .B1(new_n849_), .B2(new_n589_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n595_), .A2(new_n233_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n849_), .B2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT124), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(G1351gat));
  NAND3_X1  g668(.A1(new_n268_), .A2(new_n409_), .A3(new_n345_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n442_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g672(.A(new_n870_), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n597_), .B(new_n874_), .C1(new_n796_), .C2(new_n797_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(G204gat), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n620_), .A2(new_n314_), .ZN(new_n877_));
  AOI21_X1  g676(.A(KEYINPUT125), .B1(new_n871_), .B2(new_n877_), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n874_), .B(new_n877_), .C1(new_n796_), .C2(new_n797_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT125), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n876_), .B1(new_n878_), .B2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(KEYINPUT126), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT126), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n884_), .B(new_n876_), .C1(new_n878_), .C2(new_n881_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(G1353gat));
  NAND2_X1  g685(.A1(new_n871_), .A2(new_n546_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n887_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n888_));
  XOR2_X1   g687(.A(KEYINPUT63), .B(G211gat), .Z(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n887_), .B2(new_n889_), .ZN(G1354gat));
  AOI21_X1  g689(.A(KEYINPUT127), .B1(new_n871_), .B2(new_n595_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(G218gat), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n871_), .A2(KEYINPUT127), .A3(new_n595_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n588_), .A2(G218gat), .ZN(new_n894_));
  AOI22_X1  g693(.A1(new_n892_), .A2(new_n893_), .B1(new_n871_), .B2(new_n894_), .ZN(G1355gat));
endmodule


