//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 1 1 0 0 0 1 0 0 1 0 0 0 1 0 1 0 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n816_, new_n817_, new_n818_, new_n820_,
    new_n821_, new_n822_, new_n824_, new_n825_, new_n826_, new_n828_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n857_,
    new_n859_, new_n860_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_;
  XOR2_X1   g000(.A(G71gat), .B(G99gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G43gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT30), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT31), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT25), .B(G183gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT24), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n209_), .B1(G169gat), .B2(G176gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n210_), .B1(G169gat), .B2(G176gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT23), .ZN(new_n213_));
  OR3_X1    g012(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n208_), .A2(new_n211_), .A3(new_n213_), .A4(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n213_), .B1(G183gat), .B2(G190gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT81), .ZN(new_n217_));
  AND2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(G169gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n220_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n215_), .B1(new_n218_), .B2(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(KEYINPUT82), .B(G15gat), .Z(new_n223_));
  NAND2_X1  g022(.A1(G227gat), .A2(G233gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n223_), .B(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n222_), .B(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n205_), .B(new_n226_), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n227_), .A2(KEYINPUT83), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(KEYINPUT83), .ZN(new_n229_));
  XOR2_X1   g028(.A(G127gat), .B(G134gat), .Z(new_n230_));
  XOR2_X1   g029(.A(G113gat), .B(G120gat), .Z(new_n231_));
  XOR2_X1   g030(.A(new_n230_), .B(new_n231_), .Z(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  OR3_X1    g032(.A1(new_n228_), .A2(new_n229_), .A3(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n233_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(G1gat), .B(G29gat), .Z(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G57gat), .B(G85gat), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n239_), .B(new_n240_), .Z(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G225gat), .A2(G233gat), .ZN(new_n243_));
  NOR2_X1   g042(.A1(G141gat), .A2(G148gat), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G141gat), .A2(G148gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT1), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(G155gat), .A3(G162gat), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT85), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G155gat), .A2(G162gat), .ZN(new_n252_));
  NOR2_X1   g051(.A1(G155gat), .A2(G162gat), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n252_), .B1(new_n253_), .B2(KEYINPUT1), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n251_), .B1(KEYINPUT84), .B2(new_n254_), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n254_), .A2(KEYINPUT84), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n247_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n244_), .B(KEYINPUT3), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n246_), .B(KEYINPUT2), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT86), .ZN(new_n262_));
  INV_X1    g061(.A(new_n252_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n263_), .A2(new_n253_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n233_), .B1(new_n258_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n243_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT93), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n258_), .A2(new_n265_), .A3(new_n233_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n264_), .ZN(new_n271_));
  OR2_X1    g070(.A1(new_n261_), .A2(KEYINPUT86), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n261_), .A2(KEYINPUT86), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n271_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n232_), .B1(new_n274_), .B2(new_n257_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n270_), .A2(KEYINPUT4), .A3(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n268_), .A2(new_n269_), .A3(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n270_), .A2(new_n275_), .A3(new_n243_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n269_), .B1(new_n268_), .B2(new_n276_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n242_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n276_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n243_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n283_), .B1(new_n275_), .B2(KEYINPUT4), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT93), .B1(new_n282_), .B2(new_n284_), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n285_), .A2(new_n241_), .A3(new_n277_), .A4(new_n278_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n281_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT96), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT20), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT89), .ZN(new_n290_));
  INV_X1    g089(.A(G197gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n290_), .B1(new_n291_), .B2(G204gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT88), .B(G197gat), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n292_), .B1(new_n293_), .B2(G204gat), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(KEYINPUT89), .A3(G204gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G211gat), .B(G218gat), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT21), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n295_), .A2(new_n296_), .A3(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(KEYINPUT21), .B1(new_n295_), .B2(new_n296_), .ZN(new_n301_));
  INV_X1    g100(.A(G204gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n293_), .A2(new_n302_), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n303_), .B(KEYINPUT21), .C1(new_n291_), .C2(new_n302_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n297_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n300_), .B1(new_n301_), .B2(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n289_), .B1(new_n222_), .B2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G226gat), .A2(G233gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n216_), .A2(new_n220_), .ZN(new_n311_));
  OAI22_X1  g110(.A1(new_n210_), .A2(KEYINPUT91), .B1(G169gat), .B2(G176gat), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n312_), .B1(KEYINPUT91), .B2(new_n210_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n208_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n311_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n307_), .B(new_n310_), .C1(new_n306_), .C2(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT20), .B1(new_n222_), .B2(new_n306_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n306_), .A2(new_n315_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT92), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n306_), .A2(KEYINPUT92), .A3(new_n315_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n317_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n316_), .B1(new_n322_), .B2(new_n310_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G8gat), .B(G36gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT18), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G64gat), .B(G92gat), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n325_), .B(new_n326_), .Z(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n323_), .A2(new_n328_), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n327_), .B(new_n316_), .C1(new_n322_), .C2(new_n310_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  XOR2_X1   g130(.A(KEYINPUT97), .B(KEYINPUT27), .Z(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n330_), .A2(KEYINPUT27), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n322_), .A2(new_n310_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n310_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT95), .ZN(new_n337_));
  OR2_X1    g136(.A1(new_n315_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n306_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n315_), .A2(new_n337_), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n338_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n307_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n336_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n335_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(new_n328_), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n331_), .A2(new_n333_), .B1(new_n334_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT96), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n281_), .A2(new_n347_), .A3(new_n286_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n258_), .A2(new_n265_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n339_), .B1(new_n349_), .B2(KEYINPUT29), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(G22gat), .B(G50gat), .Z(new_n354_));
  OR3_X1    g153(.A1(new_n349_), .A2(KEYINPUT29), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G228gat), .A2(G233gat), .ZN(new_n356_));
  INV_X1    g155(.A(G78gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(G106gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n354_), .B1(new_n349_), .B2(KEYINPUT29), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n355_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n361_), .B1(new_n355_), .B2(new_n362_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n353_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n365_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n367_), .A2(new_n352_), .A3(new_n363_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  AND4_X1   g168(.A1(new_n288_), .A2(new_n346_), .A3(new_n348_), .A4(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n279_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n371_), .A2(KEYINPUT33), .A3(new_n241_), .A4(new_n285_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT33), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n286_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n331_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n270_), .A2(new_n275_), .A3(new_n283_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n243_), .B1(new_n275_), .B2(KEYINPUT4), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n242_), .B(new_n376_), .C1(new_n282_), .C2(new_n377_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n372_), .A2(new_n374_), .A3(new_n375_), .A4(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n323_), .B1(KEYINPUT32), .B2(new_n327_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n327_), .A2(KEYINPUT32), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n381_), .B1(new_n335_), .B2(new_n343_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n287_), .A2(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n369_), .B1(new_n379_), .B2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n236_), .B1(new_n370_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n236_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n288_), .A2(new_n348_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n346_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n389_), .A2(new_n369_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n387_), .A2(new_n388_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n386_), .A2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G57gat), .B(G64gat), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n393_), .A2(KEYINPUT11), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(KEYINPUT11), .ZN(new_n395_));
  XOR2_X1   g194(.A(G71gat), .B(G78gat), .Z(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n395_), .A2(new_n396_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G99gat), .A2(G106gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT6), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT6), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(G99gat), .A3(G106gat), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT7), .ZN(new_n405_));
  INV_X1    g204(.A(G99gat), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n405_), .A2(new_n406_), .A3(new_n359_), .A4(KEYINPUT64), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT64), .ZN(new_n408_));
  OAI22_X1  g207(.A1(new_n408_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT65), .B1(new_n404_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n401_), .A2(new_n403_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT65), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n412_), .A2(new_n413_), .A3(new_n409_), .A4(new_n407_), .ZN(new_n414_));
  INV_X1    g213(.A(G85gat), .ZN(new_n415_));
  INV_X1    g214(.A(G92gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G85gat), .A2(G92gat), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT8), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n419_), .A2(KEYINPUT66), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(KEYINPUT66), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n417_), .B(new_n418_), .C1(new_n420_), .C2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n411_), .A2(new_n414_), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n417_), .A2(new_n418_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n426_), .B1(new_n404_), .B2(new_n410_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT8), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n424_), .A2(new_n428_), .ZN(new_n429_));
  OR2_X1    g228(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n430_), .A2(new_n359_), .A3(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n417_), .A2(KEYINPUT9), .A3(new_n418_), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n418_), .A2(KEYINPUT9), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n412_), .A2(new_n432_), .A3(new_n433_), .A4(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT67), .B1(new_n429_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT67), .ZN(new_n437_));
  INV_X1    g236(.A(new_n435_), .ZN(new_n438_));
  AOI211_X1 g237(.A(new_n437_), .B(new_n438_), .C1(new_n424_), .C2(new_n428_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n399_), .B1(new_n436_), .B2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n402_), .B1(G99gat), .B2(G106gat), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n400_), .A2(KEYINPUT6), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n409_), .B(new_n407_), .C1(new_n441_), .C2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n422_), .B1(new_n443_), .B2(KEYINPUT65), .ZN(new_n444_));
  AOI22_X1  g243(.A1(new_n444_), .A2(new_n414_), .B1(KEYINPUT8), .B2(new_n427_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n437_), .B1(new_n445_), .B2(new_n438_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n429_), .A2(KEYINPUT67), .A3(new_n435_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n399_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n446_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n440_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G230gat), .A2(G233gat), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT68), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT12), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n449_), .A2(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(new_n435_), .B(KEYINPUT69), .Z(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n429_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(KEYINPUT12), .A3(new_n448_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n456_), .A2(new_n451_), .A3(new_n440_), .A4(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT68), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n450_), .A2(new_n461_), .A3(new_n452_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n454_), .A2(new_n460_), .A3(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G120gat), .B(G148gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT5), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G176gat), .B(G204gat), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n465_), .B(new_n466_), .Z(new_n467_));
  NAND2_X1  g266(.A1(new_n463_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n467_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n454_), .A2(new_n460_), .A3(new_n462_), .A4(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT13), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n468_), .A2(KEYINPUT13), .A3(new_n470_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G229gat), .A2(G233gat), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G29gat), .B(G36gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G43gat), .B(G50gat), .ZN(new_n479_));
  XOR2_X1   g278(.A(new_n478_), .B(new_n479_), .Z(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n478_), .B(new_n479_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n481_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n482_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G15gat), .B(G22gat), .ZN(new_n487_));
  INV_X1    g286(.A(G1gat), .ZN(new_n488_));
  INV_X1    g287(.A(G8gat), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT14), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n487_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G1gat), .B(G8gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n486_), .A2(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n493_), .B1(new_n482_), .B2(new_n485_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n477_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT80), .ZN(new_n498_));
  INV_X1    g297(.A(new_n496_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT15), .ZN(new_n500_));
  INV_X1    g299(.A(new_n485_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n483_), .A2(new_n484_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n500_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n482_), .A2(KEYINPUT15), .A3(new_n485_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n476_), .B(new_n499_), .C1(new_n505_), .C2(new_n494_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT80), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n507_), .B(new_n477_), .C1(new_n495_), .C2(new_n496_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n498_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G113gat), .B(G141gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G169gat), .B(G197gat), .ZN(new_n511_));
  XOR2_X1   g310(.A(new_n510_), .B(new_n511_), .Z(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n509_), .A2(new_n513_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n498_), .A2(new_n506_), .A3(new_n508_), .A4(new_n512_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n475_), .A2(new_n517_), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n392_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G232gat), .A2(G233gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT35), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n458_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n524_), .B1(new_n505_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n522_), .A2(new_n523_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n486_), .B1(new_n436_), .B2(new_n439_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n527_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n530_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n528_), .B1(new_n526_), .B2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G190gat), .B(G218gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT73), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G134gat), .B(G162gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT36), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n539_), .B(KEYINPUT74), .Z(new_n540_));
  AND3_X1   g339(.A1(new_n531_), .A2(new_n533_), .A3(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n537_), .B(new_n538_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT75), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n544_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT37), .B1(new_n541_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n542_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n533_), .ZN(new_n548_));
  NOR3_X1   g347(.A1(new_n526_), .A2(new_n532_), .A3(new_n528_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n547_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT37), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n531_), .A2(new_n533_), .A3(new_n540_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n550_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n546_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G231gat), .A2(G233gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n493_), .B(new_n556_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n557_), .A2(new_n448_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n448_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT76), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G127gat), .B(G155gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT16), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G183gat), .B(G211gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(KEYINPUT17), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT77), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n562_), .A2(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n566_), .B(KEYINPUT17), .Z(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT78), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n571_), .A2(new_n559_), .A3(new_n558_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n555_), .A2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT79), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n519_), .A2(new_n575_), .ZN(new_n576_));
  NOR3_X1   g375(.A1(new_n576_), .A2(G1gat), .A3(new_n388_), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n577_), .B(KEYINPUT38), .Z(new_n578_));
  NAND2_X1  g377(.A1(new_n550_), .A2(new_n552_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n580_), .A2(new_n573_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n519_), .A2(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(G1gat), .B1(new_n582_), .B2(new_n388_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n578_), .A2(new_n583_), .ZN(G1324gat));
  NOR3_X1   g383(.A1(new_n576_), .A2(G8gat), .A3(new_n346_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT98), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n586_), .B1(new_n582_), .B2(new_n346_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n519_), .A2(KEYINPUT98), .A3(new_n389_), .A4(new_n581_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n489_), .B1(KEYINPUT99), .B2(KEYINPUT39), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n587_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(KEYINPUT99), .A2(KEYINPUT39), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n585_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n591_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n587_), .A2(new_n588_), .A3(new_n589_), .A4(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n592_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n595_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(G1325gat));
  OAI21_X1  g397(.A(G15gat), .B1(new_n582_), .B2(new_n236_), .ZN(new_n599_));
  XOR2_X1   g398(.A(KEYINPUT101), .B(KEYINPUT41), .Z(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n236_), .A2(G15gat), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n601_), .B1(new_n576_), .B2(new_n602_), .ZN(G1326gat));
  INV_X1    g402(.A(new_n369_), .ZN(new_n604_));
  OAI21_X1  g403(.A(G22gat), .B1(new_n582_), .B2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT42), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n604_), .A2(G22gat), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n606_), .B1(new_n576_), .B2(new_n607_), .ZN(G1327gat));
  INV_X1    g407(.A(new_n573_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n609_), .A2(new_n579_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n392_), .A2(new_n518_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT103), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n392_), .A2(KEYINPUT103), .A3(new_n518_), .A4(new_n610_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n388_), .ZN(new_n616_));
  AOI21_X1  g415(.A(G29gat), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n518_), .A2(new_n573_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT102), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT43), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n620_), .B1(new_n392_), .B2(new_n555_), .ZN(new_n621_));
  AOI211_X1 g420(.A(KEYINPUT43), .B(new_n554_), .C1(new_n386_), .C2(new_n391_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n619_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT44), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  OAI211_X1 g424(.A(KEYINPUT44), .B(new_n619_), .C1(new_n621_), .C2(new_n622_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n616_), .A2(G29gat), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n617_), .B1(new_n627_), .B2(new_n628_), .ZN(G1328gat));
  XNOR2_X1  g428(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n625_), .A2(new_n389_), .A3(new_n626_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(G36gat), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n346_), .A2(G36gat), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n613_), .A2(new_n614_), .A3(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT45), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n632_), .A2(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n630_), .B1(new_n636_), .B2(KEYINPUT104), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT104), .ZN(new_n638_));
  INV_X1    g437(.A(new_n630_), .ZN(new_n639_));
  AOI211_X1 g438(.A(new_n638_), .B(new_n639_), .C1(new_n632_), .C2(new_n635_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n637_), .A2(new_n640_), .ZN(G1329gat));
  NAND4_X1  g440(.A1(new_n625_), .A2(G43gat), .A3(new_n387_), .A4(new_n626_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n615_), .A2(new_n387_), .ZN(new_n643_));
  XOR2_X1   g442(.A(KEYINPUT106), .B(G43gat), .Z(new_n644_));
  OAI21_X1  g443(.A(new_n642_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(G1330gat));
  AOI21_X1  g446(.A(G50gat), .B1(new_n615_), .B2(new_n369_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n369_), .A2(G50gat), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n627_), .B2(new_n649_), .ZN(G1331gat));
  INV_X1    g449(.A(G57gat), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n473_), .A2(new_n474_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n652_), .A2(new_n516_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n392_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(new_n575_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n651_), .B1(new_n655_), .B2(new_n388_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT108), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n654_), .A2(new_n581_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n658_), .A2(new_n651_), .A3(new_n388_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n657_), .A2(new_n659_), .ZN(G1332gat));
  INV_X1    g459(.A(new_n655_), .ZN(new_n661_));
  INV_X1    g460(.A(G64gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n661_), .A2(new_n662_), .A3(new_n389_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n658_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n662_), .B1(new_n664_), .B2(new_n389_), .ZN(new_n665_));
  XOR2_X1   g464(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n665_), .A2(new_n666_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n663_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT110), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OAI211_X1 g471(.A(KEYINPUT110), .B(new_n663_), .C1(new_n668_), .C2(new_n669_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1333gat));
  OAI21_X1  g473(.A(G71gat), .B1(new_n658_), .B2(new_n236_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT49), .ZN(new_n676_));
  OR3_X1    g475(.A1(new_n655_), .A2(G71gat), .A3(new_n236_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT111), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n676_), .A2(KEYINPUT111), .A3(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1334gat));
  OAI21_X1  g481(.A(G78gat), .B1(new_n658_), .B2(new_n604_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT50), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n661_), .A2(new_n357_), .A3(new_n369_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1335gat));
  NAND2_X1  g485(.A1(new_n654_), .A2(new_n610_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n688_), .A2(new_n415_), .A3(new_n616_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n621_), .A2(new_n622_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n653_), .A2(new_n573_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n690_), .A2(new_n388_), .A3(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n689_), .B1(new_n692_), .B2(new_n415_), .ZN(G1336gat));
  OAI21_X1  g492(.A(new_n416_), .B1(new_n687_), .B2(new_n346_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT112), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n695_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n690_), .A2(new_n691_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n698_), .A2(G92gat), .A3(new_n389_), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n696_), .A2(new_n697_), .A3(new_n699_), .ZN(G1337gat));
  AND4_X1   g499(.A1(new_n430_), .A2(new_n688_), .A3(new_n431_), .A4(new_n387_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n406_), .B1(new_n698_), .B2(new_n387_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT113), .ZN(new_n703_));
  OAI22_X1  g502(.A1(new_n701_), .A2(new_n702_), .B1(new_n703_), .B2(KEYINPUT51), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(KEYINPUT51), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(G1338gat));
  XNOR2_X1  g505(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT114), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT52), .ZN(new_n710_));
  OAI21_X1  g509(.A(G106gat), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n711_), .B1(new_n698_), .B2(new_n369_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n709_), .A2(new_n710_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n688_), .A2(new_n359_), .A3(new_n369_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n716_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n708_), .B1(new_n715_), .B2(new_n717_), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n712_), .A2(new_n713_), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n719_), .A2(new_n714_), .A3(new_n716_), .A4(new_n707_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1339gat));
  INV_X1    g520(.A(KEYINPUT122), .ZN(new_n722_));
  INV_X1    g521(.A(G113gat), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n517_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n470_), .A2(new_n516_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n436_), .A2(new_n439_), .ZN(new_n727_));
  AOI21_X1  g526(.A(KEYINPUT12), .B1(new_n727_), .B2(new_n448_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n440_), .A2(new_n459_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n452_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT118), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT117), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT55), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n460_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  OAI211_X1 g534(.A(KEYINPUT118), .B(new_n452_), .C1(new_n728_), .C2(new_n729_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n732_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n734_), .B1(new_n460_), .B2(new_n733_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n467_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT56), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n460_), .A2(new_n733_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT55), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n743_), .A2(new_n735_), .A3(new_n732_), .A4(new_n736_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n744_), .A2(KEYINPUT56), .A3(new_n467_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n726_), .B1(new_n741_), .B2(new_n745_), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n477_), .B(new_n499_), .C1(new_n505_), .C2(new_n494_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n476_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n747_), .A2(new_n513_), .A3(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n515_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT119), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT119), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n515_), .A2(new_n749_), .A3(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n471_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  OAI211_X1 g555(.A(KEYINPUT57), .B(new_n579_), .C1(new_n746_), .C2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT121), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n754_), .A2(new_n470_), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n744_), .A2(KEYINPUT56), .A3(new_n467_), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT56), .B1(new_n744_), .B2(new_n467_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n759_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT58), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n554_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n741_), .A2(new_n745_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n765_), .A2(KEYINPUT120), .A3(KEYINPUT58), .A4(new_n759_), .ZN(new_n766_));
  OAI211_X1 g565(.A(KEYINPUT58), .B(new_n759_), .C1(new_n760_), .C2(new_n761_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT120), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n764_), .A2(new_n766_), .A3(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n579_), .B1(new_n746_), .B2(new_n756_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT57), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n726_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n774_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n755_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT121), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n776_), .A2(new_n777_), .A3(KEYINPUT57), .A4(new_n579_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n758_), .A2(new_n770_), .A3(new_n773_), .A4(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n573_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT54), .ZN(new_n781_));
  AOI211_X1 g580(.A(new_n516_), .B(new_n573_), .C1(new_n546_), .C2(new_n553_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n652_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n783_), .B1(new_n652_), .B2(new_n782_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n781_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n786_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n788_), .A2(new_n784_), .A3(KEYINPUT54), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n780_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n387_), .A2(new_n390_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n791_), .A2(new_n616_), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT59), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n388_), .B1(new_n780_), .B2(new_n790_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n797_), .A2(KEYINPUT59), .A3(new_n793_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n725_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n794_), .ZN(new_n800_));
  AOI21_X1  g599(.A(G113gat), .B1(new_n800_), .B2(new_n516_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n722_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n787_), .A2(new_n789_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n803_), .B1(new_n573_), .B2(new_n779_), .ZN(new_n804_));
  NOR4_X1   g603(.A1(new_n804_), .A2(new_n795_), .A3(new_n388_), .A4(new_n792_), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT59), .B1(new_n797_), .B2(new_n793_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n724_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n723_), .B1(new_n794_), .B2(new_n517_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(KEYINPUT122), .A3(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n802_), .A2(new_n809_), .ZN(G1340gat));
  INV_X1    g609(.A(G120gat), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n652_), .B2(KEYINPUT60), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n800_), .B(new_n812_), .C1(KEYINPUT60), .C2(new_n811_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n652_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(new_n811_), .ZN(G1341gat));
  INV_X1    g614(.A(G127gat), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n800_), .A2(new_n816_), .A3(new_n609_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n573_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n818_), .B2(new_n816_), .ZN(G1342gat));
  INV_X1    g618(.A(G134gat), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n800_), .A2(new_n820_), .A3(new_n580_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n554_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n822_), .B2(new_n820_), .ZN(G1343gat));
  NOR3_X1   g622(.A1(new_n387_), .A2(new_n604_), .A3(new_n389_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n797_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n516_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n475_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g628(.A1(new_n797_), .A2(new_n609_), .A3(new_n824_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT123), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n797_), .A2(KEYINPUT123), .A3(new_n609_), .A4(new_n824_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(KEYINPUT61), .B(G155gat), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n832_), .A2(new_n833_), .A3(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n835_), .A2(new_n836_), .ZN(G1346gat));
  INV_X1    g636(.A(G162gat), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n825_), .A2(new_n838_), .A3(new_n580_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n825_), .A2(new_n555_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(new_n838_), .ZN(G1347gat));
  NOR2_X1   g640(.A1(new_n804_), .A2(new_n346_), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n616_), .A2(new_n369_), .A3(new_n236_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n516_), .A3(new_n843_), .ZN(new_n844_));
  OAI211_X1 g643(.A(KEYINPUT62), .B(G169gat), .C1(new_n844_), .C2(KEYINPUT22), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT62), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n842_), .A2(new_n516_), .A3(new_n843_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT22), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n846_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(G169gat), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n850_), .B1(new_n847_), .B2(new_n846_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n845_), .B1(new_n849_), .B2(new_n851_), .ZN(G1348gat));
  NAND2_X1  g651(.A1(new_n842_), .A2(new_n843_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(new_n652_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(KEYINPUT124), .B(G176gat), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n854_), .B(new_n855_), .ZN(G1349gat));
  NAND3_X1  g655(.A1(new_n842_), .A2(new_n609_), .A3(new_n843_), .ZN(new_n857_));
  MUX2_X1   g656(.A(new_n206_), .B(G183gat), .S(new_n857_), .Z(G1350gat));
  OAI21_X1  g657(.A(G190gat), .B1(new_n853_), .B2(new_n554_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n580_), .A2(new_n207_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n853_), .B2(new_n860_), .ZN(G1351gat));
  NOR2_X1   g660(.A1(new_n616_), .A2(new_n604_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n842_), .A2(new_n862_), .A3(new_n236_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(new_n517_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT125), .B(G197gat), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1352gat));
  NAND2_X1  g665(.A1(new_n791_), .A2(new_n389_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n862_), .A2(new_n236_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n475_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g670(.A(new_n573_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n872_));
  XOR2_X1   g671(.A(new_n872_), .B(KEYINPUT126), .Z(new_n873_));
  NOR2_X1   g672(.A1(new_n863_), .A2(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1354gat));
  NOR3_X1   g675(.A1(new_n867_), .A2(new_n579_), .A3(new_n868_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT127), .ZN(new_n878_));
  AOI21_X1  g677(.A(G218gat), .B1(new_n877_), .B2(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(KEYINPUT127), .B1(new_n863_), .B2(new_n579_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n555_), .A2(G218gat), .ZN(new_n881_));
  AOI22_X1  g680(.A1(new_n879_), .A2(new_n880_), .B1(new_n869_), .B2(new_n881_), .ZN(G1355gat));
endmodule


