//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 1 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n763_, new_n764_,
    new_n765_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n935_,
    new_n936_, new_n937_, new_n939_, new_n940_, new_n942_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n962_, new_n963_, new_n964_;
  OR4_X1    g000(.A1(KEYINPUT92), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT2), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G141gat), .ZN(new_n206_));
  INV_X1    g005(.A(G148gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n208_), .B1(KEYINPUT92), .B2(KEYINPUT3), .ZN(new_n209_));
  NAND3_X1  g008(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n202_), .A2(new_n205_), .A3(new_n209_), .A4(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(KEYINPUT1), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(new_n212_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n213_), .A2(KEYINPUT1), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n208_), .B(new_n203_), .C1(new_n216_), .C2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT29), .ZN(new_n220_));
  XOR2_X1   g019(.A(G197gat), .B(G204gat), .Z(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT21), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G211gat), .B(G218gat), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n221_), .A2(KEYINPUT21), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT93), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n227_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NOR3_X1   g028(.A1(new_n222_), .A2(new_n227_), .A3(new_n223_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n226_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n220_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G228gat), .ZN(new_n233_));
  INV_X1    g032(.A(G233gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n232_), .A2(new_n235_), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n231_), .B(new_n220_), .C1(new_n233_), .C2(new_n234_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G78gat), .B(G106gat), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n236_), .A2(new_n237_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT94), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n219_), .A2(KEYINPUT29), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G22gat), .B(G50gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT28), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n242_), .B(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n241_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n236_), .A2(new_n237_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(new_n238_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(new_n240_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n241_), .A2(new_n248_), .A3(new_n240_), .A4(new_n245_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G127gat), .B(G134gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G113gat), .B(G120gat), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT90), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n253_), .A2(new_n254_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT89), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  OR3_X1    g059(.A1(new_n257_), .A2(new_n260_), .A3(KEYINPUT91), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT91), .B1(new_n257_), .B2(new_n260_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  XOR2_X1   g062(.A(new_n263_), .B(KEYINPUT31), .Z(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G227gat), .A2(G233gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(G15gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT87), .B(G43gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  XOR2_X1   g068(.A(G71gat), .B(G99gat), .Z(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT23), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n272_), .A2(G183gat), .A3(G190gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT84), .ZN(new_n274_));
  INV_X1    g073(.A(G183gat), .ZN(new_n275_));
  INV_X1    g074(.A(G190gat), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT23), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n274_), .A2(new_n277_), .ZN(new_n278_));
  OR2_X1    g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n279_), .A2(KEYINPUT24), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT85), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n278_), .A2(KEYINPUT85), .A3(new_n280_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT25), .B(G183gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT83), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n286_), .B1(new_n276_), .B2(KEYINPUT26), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT26), .B(G190gat), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n285_), .B(new_n287_), .C1(new_n288_), .C2(new_n286_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n279_), .A2(KEYINPUT24), .A3(new_n290_), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n283_), .A2(new_n284_), .A3(new_n289_), .A4(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(KEYINPUT86), .B(G176gat), .Z(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT22), .B(G169gat), .ZN(new_n294_));
  AOI22_X1  g093(.A1(new_n293_), .A2(new_n294_), .B1(G169gat), .B2(G176gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n277_), .A2(new_n273_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n295_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n292_), .A2(KEYINPUT30), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(KEYINPUT30), .B1(new_n292_), .B2(new_n300_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT88), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n292_), .A2(new_n300_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT30), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT88), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n307_), .A2(new_n308_), .A3(new_n301_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n271_), .B1(new_n304_), .B2(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n308_), .B1(new_n307_), .B2(new_n301_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n271_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n265_), .B1(new_n310_), .B2(new_n313_), .ZN(new_n314_));
  NOR3_X1   g113(.A1(new_n302_), .A2(new_n303_), .A3(KEYINPUT88), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n312_), .B1(new_n315_), .B2(new_n311_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n304_), .A2(new_n271_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n316_), .A2(new_n317_), .A3(new_n264_), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n252_), .A2(new_n314_), .A3(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n252_), .B1(new_n318_), .B2(new_n314_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(G8gat), .B(G36gat), .Z(new_n322_));
  XNOR2_X1  g121(.A(G64gat), .B(G92gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n288_), .A2(new_n285_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(new_n291_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT95), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n330_), .A2(new_n296_), .A3(new_n280_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n230_), .ZN(new_n332_));
  AOI22_X1  g131(.A1(new_n332_), .A2(new_n228_), .B1(new_n225_), .B2(new_n224_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n278_), .A2(new_n298_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n295_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n331_), .A2(new_n333_), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G226gat), .A2(G233gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT19), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n336_), .A2(KEYINPUT20), .A3(new_n339_), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n284_), .A2(new_n289_), .A3(new_n291_), .ZN(new_n341_));
  AOI22_X1  g140(.A1(new_n341_), .A2(new_n283_), .B1(new_n295_), .B2(new_n299_), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT96), .B1(new_n342_), .B2(new_n333_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT96), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n305_), .A2(new_n344_), .A3(new_n231_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n340_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n342_), .A2(new_n333_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT20), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n331_), .A2(new_n335_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n348_), .B1(new_n349_), .B2(new_n231_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n339_), .B1(new_n347_), .B2(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n327_), .B1(new_n346_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n340_), .ZN(new_n353_));
  NOR3_X1   g152(.A1(new_n342_), .A2(KEYINPUT96), .A3(new_n333_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n344_), .B1(new_n305_), .B2(new_n231_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n353_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n347_), .A2(new_n350_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(new_n338_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n356_), .A2(new_n358_), .A3(new_n326_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n352_), .A2(new_n359_), .A3(KEYINPUT98), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT27), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n356_), .A2(new_n358_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT98), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(new_n363_), .A3(new_n327_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n360_), .A2(new_n361_), .A3(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n357_), .A2(new_n338_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n336_), .A2(KEYINPUT20), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT102), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT102), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n336_), .A2(new_n369_), .A3(KEYINPUT20), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n368_), .B(new_n370_), .C1(new_n354_), .C2(new_n355_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n366_), .B1(new_n371_), .B2(new_n338_), .ZN(new_n372_));
  OAI211_X1 g171(.A(KEYINPUT27), .B(new_n359_), .C1(new_n372_), .C2(new_n326_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n365_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G225gat), .A2(G233gat), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n263_), .A2(new_n219_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n258_), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n380_), .A2(new_n255_), .ZN(new_n381_));
  OR2_X1    g180(.A1(new_n381_), .A2(KEYINPUT100), .ZN(new_n382_));
  INV_X1    g181(.A(new_n219_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n381_), .A2(KEYINPUT100), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT99), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n377_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n263_), .A2(KEYINPUT99), .A3(new_n219_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n386_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n376_), .B(new_n379_), .C1(new_n390_), .C2(new_n378_), .ZN(new_n391_));
  AOI21_X1  g190(.A(KEYINPUT99), .B1(new_n263_), .B2(new_n219_), .ZN(new_n392_));
  AOI211_X1 g191(.A(new_n387_), .B(new_n383_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n385_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n375_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n391_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G1gat), .B(G29gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(G85gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT0), .B(G57gat), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n398_), .B(new_n399_), .Z(new_n400_));
  NAND2_X1  g199(.A1(new_n396_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n400_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n391_), .A2(new_n402_), .A3(new_n395_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  NOR3_X1   g203(.A1(new_n321_), .A2(new_n374_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n326_), .A2(KEYINPUT32), .ZN(new_n406_));
  MUX2_X1   g205(.A(new_n372_), .B(new_n362_), .S(new_n406_), .Z(new_n407_));
  NAND2_X1  g206(.A1(new_n404_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT101), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n402_), .B1(new_n391_), .B2(new_n395_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n409_), .B1(new_n410_), .B2(KEYINPUT33), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT33), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n394_), .A2(new_n375_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n379_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n414_), .B1(new_n394_), .B2(KEYINPUT4), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n413_), .B1(new_n376_), .B2(new_n415_), .ZN(new_n416_));
  OAI211_X1 g215(.A(KEYINPUT101), .B(new_n412_), .C1(new_n416_), .C2(new_n402_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n411_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n410_), .A2(KEYINPUT33), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n415_), .A2(new_n376_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n402_), .B1(new_n394_), .B2(new_n375_), .ZN(new_n421_));
  OR2_X1    g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n360_), .A2(new_n364_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n419_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n408_), .B1(new_n418_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n314_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n318_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n252_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n405_), .B1(new_n425_), .B2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G15gat), .B(G22gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G1gat), .B(G8gat), .ZN(new_n433_));
  INV_X1    g232(.A(G8gat), .ZN(new_n434_));
  INV_X1    g233(.A(G1gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT74), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT74), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(G1gat), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n434_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT14), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n432_), .B(new_n433_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT74), .B(G1gat), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT14), .B1(new_n443_), .B2(new_n434_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n433_), .B1(new_n444_), .B2(new_n432_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n442_), .A2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G43gat), .B(G50gat), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(G36gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(G29gat), .ZN(new_n450_));
  INV_X1    g249(.A(G29gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(G36gat), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT71), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n450_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n453_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n448_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n450_), .A2(new_n452_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT71), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n450_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(new_n459_), .A3(new_n447_), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n456_), .A2(new_n460_), .A3(KEYINPUT15), .ZN(new_n461_));
  AOI21_X1  g260(.A(KEYINPUT15), .B1(new_n456_), .B2(new_n460_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n446_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n456_), .A2(new_n460_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n465_), .B1(new_n442_), .B2(new_n445_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G229gat), .A2(G233gat), .ZN(new_n467_));
  XOR2_X1   g266(.A(new_n467_), .B(KEYINPUT80), .Z(new_n468_));
  NAND3_X1  g267(.A1(new_n463_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT81), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n444_), .A2(new_n432_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n433_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n473_), .A2(new_n464_), .A3(new_n441_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n464_), .B1(new_n473_), .B2(new_n441_), .ZN(new_n475_));
  OAI211_X1 g274(.A(G229gat), .B(G233gat), .C1(new_n474_), .C2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT81), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n463_), .A2(new_n466_), .A3(new_n477_), .A4(new_n468_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G113gat), .B(G141gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G169gat), .B(G197gat), .ZN(new_n480_));
  XOR2_X1   g279(.A(new_n479_), .B(new_n480_), .Z(new_n481_));
  NAND4_X1  g280(.A1(new_n470_), .A2(new_n476_), .A3(new_n478_), .A4(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT82), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n478_), .A2(new_n476_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n485_), .A2(KEYINPUT82), .A3(new_n470_), .A4(new_n481_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n470_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n481_), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n484_), .A2(new_n486_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n431_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G127gat), .B(G155gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT16), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G183gat), .B(G211gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT17), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n495_), .B(KEYINPUT77), .Z(new_n496_));
  XNOR2_X1  g295(.A(G57gat), .B(G64gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G71gat), .B(G78gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n497_), .A2(new_n498_), .A3(KEYINPUT11), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(KEYINPUT11), .ZN(new_n500_));
  INV_X1    g299(.A(new_n498_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n497_), .A2(KEYINPUT11), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n499_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(KEYINPUT75), .B(KEYINPUT76), .Z(new_n505_));
  NAND2_X1  g304(.A1(G231gat), .A2(G233gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n504_), .B(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(new_n446_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n496_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT78), .ZN(new_n511_));
  INV_X1    g310(.A(new_n509_), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n494_), .A2(KEYINPUT17), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(new_n495_), .A3(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n511_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT37), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G190gat), .B(G218gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G134gat), .B(G162gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n520_), .A2(KEYINPUT36), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G232gat), .A2(G233gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT34), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT35), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT72), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n524_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n527_), .A2(KEYINPUT72), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT7), .ZN(new_n529_));
  INV_X1    g328(.A(G99gat), .ZN(new_n530_));
  INV_X1    g329(.A(G106gat), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n529_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  AND2_X1   g331(.A1(G99gat), .A2(G106gat), .ZN(new_n533_));
  AND2_X1   g332(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n534_));
  NOR2_X1   g333(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n533_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT67), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT6), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G99gat), .A2(G106gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n543_));
  AND4_X1   g342(.A1(new_n532_), .A2(new_n536_), .A3(new_n542_), .A4(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G85gat), .B(G92gat), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT8), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(new_n531_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n538_), .A2(KEYINPUT66), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT66), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT6), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n553_), .A2(new_n555_), .A3(new_n533_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n533_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n552_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  AND2_X1   g357(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n559_));
  NOR2_X1   g358(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n560_));
  OAI21_X1  g359(.A(G92gat), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT9), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(G92gat), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n561_), .A2(new_n562_), .B1(new_n545_), .B2(new_n564_), .ZN(new_n565_));
  OAI22_X1  g364(.A1(new_n544_), .A2(new_n548_), .B1(new_n558_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n532_), .A2(new_n543_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n568_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n545_), .ZN(new_n570_));
  AOI21_X1  g369(.A(KEYINPUT8), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT68), .B1(new_n566_), .B2(new_n571_), .ZN(new_n572_));
  AND2_X1   g371(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n573_));
  NOR3_X1   g372(.A1(new_n573_), .A2(new_n549_), .A3(G106gat), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n554_), .A2(KEYINPUT6), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n538_), .A2(KEYINPUT66), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n540_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n553_), .A2(new_n555_), .A3(new_n533_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n574_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  AND2_X1   g378(.A1(G85gat), .A2(G92gat), .ZN(new_n580_));
  NOR2_X1   g379(.A1(G85gat), .A2(G92gat), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n564_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(G92gat), .ZN(new_n583_));
  OR2_X1    g382(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n584_));
  NAND2_X1  g383(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n583_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(KEYINPUT64), .B(KEYINPUT9), .Z(new_n587_));
  OAI21_X1  g386(.A(new_n582_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n536_), .A2(new_n542_), .A3(new_n532_), .A4(new_n543_), .ZN(new_n589_));
  AOI22_X1  g388(.A1(new_n579_), .A2(new_n588_), .B1(new_n589_), .B2(new_n547_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n567_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n546_), .B1(new_n591_), .B2(new_n545_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT68), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n590_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n572_), .B(new_n594_), .C1(new_n461_), .C2(new_n462_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n523_), .A2(KEYINPUT35), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n566_), .A2(new_n571_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n596_), .B1(new_n597_), .B2(new_n465_), .ZN(new_n598_));
  AOI211_X1 g397(.A(new_n526_), .B(new_n528_), .C1(new_n595_), .C2(new_n598_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n595_), .A2(new_n598_), .A3(KEYINPUT72), .A4(new_n527_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n521_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n528_), .B1(new_n595_), .B2(new_n598_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n526_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n520_), .B(KEYINPUT36), .Z(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT73), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n605_), .A2(new_n600_), .A3(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n517_), .B1(new_n602_), .B2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n605_), .A2(new_n600_), .A3(new_n606_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n602_), .A2(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n609_), .B1(new_n517_), .B2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n516_), .A2(new_n612_), .ZN(new_n613_));
  OAI211_X1 g412(.A(KEYINPUT12), .B(new_n499_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n572_), .A2(new_n594_), .A3(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n590_), .A2(new_n592_), .A3(new_n504_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G230gat), .A2(G233gat), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n504_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n620_), .B1(new_n566_), .B2(new_n571_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT12), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n616_), .A2(new_n619_), .A3(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n621_), .A2(new_n617_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n618_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n624_), .A2(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(G120gat), .B(G148gat), .Z(new_n629_));
  XNOR2_X1  g428(.A(G176gat), .B(G204gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT69), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n628_), .B(new_n635_), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n636_), .A2(KEYINPUT13), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(KEYINPUT13), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n613_), .A2(new_n639_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT79), .Z(new_n641_));
  AND2_X1   g440(.A1(new_n490_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n642_), .A2(new_n404_), .A3(new_n443_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT38), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n431_), .A2(new_n611_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n639_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n647_), .A2(new_n489_), .A3(new_n516_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n404_), .ZN(new_n650_));
  OAI21_X1  g449(.A(G1gat), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n643_), .A2(new_n644_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n645_), .A2(new_n651_), .A3(new_n652_), .ZN(G1324gat));
  NAND3_X1  g452(.A1(new_n642_), .A2(new_n434_), .A3(new_n374_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n646_), .A2(new_n374_), .A3(new_n648_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT39), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(new_n656_), .A3(G8gat), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n656_), .B1(new_n655_), .B2(G8gat), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n654_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g460(.A(new_n428_), .ZN(new_n662_));
  OAI21_X1  g461(.A(G15gat), .B1(new_n649_), .B2(new_n662_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT41), .Z(new_n664_));
  INV_X1    g463(.A(G15gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n642_), .A2(new_n665_), .A3(new_n428_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(G1326gat));
  OAI21_X1  g466(.A(G22gat), .B1(new_n649_), .B2(new_n252_), .ZN(new_n668_));
  XOR2_X1   g467(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n669_));
  XNOR2_X1  g468(.A(new_n668_), .B(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(G22gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n642_), .A2(new_n671_), .A3(new_n429_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(G1327gat));
  INV_X1    g472(.A(new_n611_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n647_), .A2(new_n515_), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n490_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n677_), .A2(new_n451_), .A3(new_n404_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n647_), .A2(new_n489_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(new_n516_), .ZN(new_n680_));
  XOR2_X1   g479(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n681_));
  XNOR2_X1  g480(.A(new_n612_), .B(KEYINPUT105), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n681_), .B1(new_n431_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n612_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n684_), .A2(KEYINPUT43), .ZN(new_n685_));
  INV_X1    g484(.A(new_n430_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n420_), .A2(new_n421_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n410_), .B2(KEYINPUT33), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n688_), .A2(new_n411_), .A3(new_n417_), .A4(new_n423_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n686_), .B1(new_n689_), .B2(new_n408_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n685_), .B1(new_n690_), .B2(new_n405_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n680_), .B1(new_n683_), .B2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT106), .B1(new_n692_), .B2(KEYINPUT44), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695_));
  INV_X1    g494(.A(new_n682_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n696_), .B1(new_n690_), .B2(new_n405_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n425_), .A2(new_n430_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n405_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  AOI22_X1  g499(.A1(new_n697_), .A2(new_n681_), .B1(new_n700_), .B2(new_n685_), .ZN(new_n701_));
  OAI211_X1 g500(.A(new_n694_), .B(new_n695_), .C1(new_n701_), .C2(new_n680_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n693_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT107), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n650_), .B1(new_n692_), .B2(KEYINPUT44), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n703_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(G29gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n704_), .B1(new_n703_), .B2(new_n705_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n678_), .B1(new_n707_), .B2(new_n708_), .ZN(G1328gat));
  NOR2_X1   g508(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n710_));
  INV_X1    g509(.A(new_n374_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n711_), .B1(new_n692_), .B2(KEYINPUT44), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n449_), .B1(new_n703_), .B2(new_n712_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n711_), .A2(G36gat), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  OR3_X1    g514(.A1(new_n676_), .A2(KEYINPUT45), .A3(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(KEYINPUT45), .B1(new_n676_), .B2(new_n715_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n710_), .B1(new_n713_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n710_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n683_), .A2(new_n691_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n680_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n722_), .A2(KEYINPUT44), .A3(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(new_n374_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n693_), .B2(new_n702_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n721_), .B(new_n718_), .C1(new_n726_), .C2(new_n449_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n720_), .A2(new_n727_), .ZN(G1329gat));
  NAND3_X1  g527(.A1(new_n724_), .A2(G43gat), .A3(new_n428_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n729_), .B1(new_n693_), .B2(new_n702_), .ZN(new_n730_));
  AOI21_X1  g529(.A(G43gat), .B1(new_n677_), .B2(new_n428_), .ZN(new_n731_));
  OAI21_X1  g530(.A(KEYINPUT47), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n729_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n731_), .B1(new_n733_), .B2(new_n703_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT47), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n732_), .A2(new_n736_), .ZN(G1330gat));
  OR3_X1    g536(.A1(new_n676_), .A2(G50gat), .A3(new_n252_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n252_), .B1(new_n692_), .B2(KEYINPUT44), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n703_), .A2(KEYINPUT109), .A3(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(G50gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT109), .B1(new_n703_), .B2(new_n739_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n738_), .B1(new_n741_), .B2(new_n742_), .ZN(G1331gat));
  NAND2_X1  g542(.A1(new_n484_), .A2(new_n486_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n487_), .A2(new_n488_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n639_), .A2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n646_), .A2(new_n515_), .A3(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G57gat), .B1(new_n748_), .B2(new_n650_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n431_), .A2(new_n746_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n750_), .A2(new_n647_), .A3(new_n613_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n650_), .A2(G57gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n749_), .B1(new_n751_), .B2(new_n752_), .ZN(G1332gat));
  OAI21_X1  g552(.A(G64gat), .B1(new_n748_), .B2(new_n711_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT48), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n711_), .A2(G64gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n755_), .B1(new_n751_), .B2(new_n756_), .ZN(G1333gat));
  OAI21_X1  g556(.A(G71gat), .B1(new_n748_), .B2(new_n662_), .ZN(new_n758_));
  XOR2_X1   g557(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n759_));
  XNOR2_X1  g558(.A(new_n758_), .B(new_n759_), .ZN(new_n760_));
  OR2_X1    g559(.A1(new_n662_), .A2(G71gat), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n751_), .B2(new_n761_), .ZN(G1334gat));
  OAI21_X1  g561(.A(G78gat), .B1(new_n748_), .B2(new_n252_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT50), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n252_), .A2(G78gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n751_), .B2(new_n765_), .ZN(G1335gat));
  NAND4_X1  g565(.A1(new_n750_), .A2(new_n647_), .A3(new_n516_), .A4(new_n611_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(G85gat), .B1(new_n768_), .B2(new_n404_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n747_), .A2(new_n516_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n770_), .B1(new_n683_), .B2(new_n691_), .ZN(new_n771_));
  XOR2_X1   g570(.A(new_n771_), .B(KEYINPUT111), .Z(new_n772_));
  AOI21_X1  g571(.A(new_n650_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(G1336gat));
  NAND3_X1  g573(.A1(new_n768_), .A2(new_n583_), .A3(new_n374_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n772_), .A2(new_n374_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(new_n583_), .ZN(G1337gat));
  NAND4_X1  g576(.A1(new_n768_), .A2(new_n428_), .A3(new_n550_), .A4(new_n551_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n701_), .A2(new_n662_), .A3(new_n770_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(new_n530_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT113), .B1(KEYINPUT112), .B2(KEYINPUT51), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n778_), .B(new_n781_), .C1(new_n530_), .C2(new_n779_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n783_), .A2(new_n784_), .A3(new_n785_), .ZN(G1338gat));
  NAND3_X1  g585(.A1(new_n768_), .A2(new_n531_), .A3(new_n429_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n771_), .A2(new_n429_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n790_), .B2(G106gat), .ZN(new_n791_));
  AOI211_X1 g590(.A(new_n531_), .B(new_n788_), .C1(new_n771_), .C2(new_n429_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n787_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT53), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n795_), .B(new_n787_), .C1(new_n791_), .C2(new_n792_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(G1339gat));
  NAND2_X1  g596(.A1(new_n711_), .A2(new_n404_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n319_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT57), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n628_), .A2(new_n634_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n746_), .A2(new_n802_), .A3(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n616_), .A2(new_n617_), .A3(new_n623_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n626_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n624_), .A2(new_n808_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n616_), .A2(new_n619_), .A3(new_n623_), .A4(KEYINPUT55), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n807_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n634_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT56), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n811_), .A2(KEYINPUT56), .A3(new_n634_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(KEYINPUT115), .B1(new_n489_), .B2(new_n803_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n805_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n468_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n463_), .A2(new_n466_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n819_), .B(new_n488_), .C1(new_n820_), .C2(new_n468_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n744_), .A2(new_n821_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n822_), .A2(new_n636_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n611_), .B1(new_n818_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n801_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n803_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n828_), .A2(new_n802_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n823_), .B1(new_n829_), .B2(new_n817_), .ZN(new_n830_));
  OAI211_X1 g629(.A(KEYINPUT116), .B(KEYINPUT57), .C1(new_n830_), .C2(new_n611_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n827_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT58), .ZN(new_n833_));
  INV_X1    g632(.A(new_n815_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT56), .B1(new_n811_), .B2(new_n634_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n744_), .A2(new_n804_), .A3(new_n821_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n833_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n612_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n837_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT58), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n612_), .B(KEYINPUT117), .C1(new_n842_), .C2(KEYINPUT58), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n841_), .A2(KEYINPUT118), .A3(new_n843_), .A4(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n843_), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT117), .B1(new_n838_), .B2(new_n612_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n846_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n832_), .A2(new_n845_), .A3(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT119), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n832_), .A2(new_n845_), .A3(new_n849_), .A4(KEYINPUT119), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(new_n516_), .A3(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n613_), .A2(new_n489_), .A3(new_n639_), .ZN(new_n855_));
  XOR2_X1   g654(.A(new_n855_), .B(KEYINPUT54), .Z(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n800_), .B1(new_n854_), .B2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(G113gat), .B1(new_n858_), .B2(new_n746_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n858_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n841_), .A2(new_n843_), .A3(new_n844_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n515_), .B1(new_n832_), .B2(new_n861_), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n856_), .A2(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n800_), .A2(KEYINPUT59), .ZN(new_n864_));
  AOI22_X1  g663(.A1(new_n860_), .A2(KEYINPUT59), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n746_), .A2(G113gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(KEYINPUT120), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n859_), .B1(new_n865_), .B2(new_n867_), .ZN(G1340gat));
  INV_X1    g667(.A(G120gat), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(new_n639_), .B2(KEYINPUT60), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n858_), .B(new_n870_), .C1(KEYINPUT60), .C2(new_n869_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n863_), .A2(new_n864_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n647_), .B(new_n872_), .C1(new_n858_), .C2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n871_), .B1(new_n875_), .B2(new_n869_), .ZN(G1341gat));
  NAND2_X1  g675(.A1(new_n854_), .A2(new_n857_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n800_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n877_), .A2(new_n515_), .A3(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(G127gat), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n515_), .A2(G127gat), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n872_), .B(new_n883_), .C1(new_n858_), .C2(new_n873_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n881_), .A2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(KEYINPUT121), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n881_), .A2(new_n884_), .A3(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n888_), .ZN(G1342gat));
  NAND3_X1  g688(.A1(new_n877_), .A2(new_n611_), .A3(new_n878_), .ZN(new_n890_));
  INV_X1    g689(.A(G134gat), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  XOR2_X1   g691(.A(KEYINPUT122), .B(G134gat), .Z(new_n893_));
  NOR2_X1   g692(.A1(new_n684_), .A2(new_n893_), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n872_), .B(new_n894_), .C1(new_n858_), .C2(new_n873_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n892_), .A2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT123), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n892_), .A2(new_n895_), .A3(KEYINPUT123), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1343gat));
  AND3_X1   g699(.A1(new_n877_), .A2(new_n320_), .A3(new_n799_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(G141gat), .B1(new_n902_), .B2(new_n489_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n901_), .A2(new_n206_), .A3(new_n746_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1344gat));
  OAI21_X1  g704(.A(G148gat), .B1(new_n902_), .B2(new_n639_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n901_), .A2(new_n207_), .A3(new_n647_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(G1345gat));
  XNOR2_X1  g707(.A(KEYINPUT61), .B(G155gat), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n909_), .B1(new_n902_), .B2(new_n516_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n909_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n901_), .A2(new_n515_), .A3(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n910_), .A2(new_n912_), .ZN(G1346gat));
  AOI21_X1  g712(.A(G162gat), .B1(new_n901_), .B2(new_n611_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n696_), .A2(G162gat), .ZN(new_n915_));
  XOR2_X1   g714(.A(new_n915_), .B(KEYINPUT124), .Z(new_n916_));
  AOI21_X1  g715(.A(new_n914_), .B1(new_n901_), .B2(new_n916_), .ZN(G1347gat));
  INV_X1    g716(.A(G169gat), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n711_), .A2(new_n404_), .ZN(new_n919_));
  AND2_X1   g718(.A1(new_n919_), .A2(new_n319_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n863_), .A2(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n918_), .B1(new_n922_), .B2(new_n746_), .ZN(new_n923_));
  OR2_X1    g722(.A1(new_n923_), .A2(KEYINPUT62), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n922_), .A2(new_n294_), .A3(new_n746_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n923_), .A2(KEYINPUT62), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n924_), .A2(new_n925_), .A3(new_n926_), .ZN(G1348gat));
  NAND3_X1  g726(.A1(new_n863_), .A2(new_n647_), .A3(new_n920_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n293_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n877_), .A2(new_n252_), .ZN(new_n930_));
  NAND4_X1  g729(.A1(new_n919_), .A2(G176gat), .A3(new_n428_), .A4(new_n647_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n929_), .B1(new_n930_), .B2(new_n931_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT125), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n932_), .B(new_n933_), .ZN(G1349gat));
  NOR3_X1   g733(.A1(new_n921_), .A2(new_n285_), .A3(new_n516_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n919_), .A2(new_n428_), .A3(new_n515_), .ZN(new_n936_));
  OR2_X1    g735(.A1(new_n930_), .A2(new_n936_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n935_), .B1(new_n937_), .B2(new_n275_), .ZN(G1350gat));
  OAI21_X1  g737(.A(G190gat), .B1(new_n921_), .B2(new_n684_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n611_), .A2(new_n288_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n921_), .B2(new_n940_), .ZN(G1351gat));
  NAND4_X1  g740(.A1(new_n877_), .A2(new_n320_), .A3(new_n746_), .A4(new_n919_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g742(.A(G204gat), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n944_), .A2(KEYINPUT126), .ZN(new_n945_));
  AND2_X1   g744(.A1(new_n877_), .A2(new_n320_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(new_n919_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n945_), .B1(new_n947_), .B2(new_n639_), .ZN(new_n948_));
  INV_X1    g747(.A(new_n945_), .ZN(new_n949_));
  NAND4_X1  g748(.A1(new_n946_), .A2(new_n647_), .A3(new_n919_), .A4(new_n949_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n948_), .A2(new_n950_), .ZN(G1353gat));
  NOR2_X1   g750(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n952_), .B(KEYINPUT127), .ZN(new_n953_));
  INV_X1    g752(.A(new_n953_), .ZN(new_n954_));
  INV_X1    g753(.A(KEYINPUT63), .ZN(new_n955_));
  INV_X1    g754(.A(G211gat), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n515_), .B1(new_n955_), .B2(new_n956_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n954_), .B1(new_n947_), .B2(new_n957_), .ZN(new_n958_));
  INV_X1    g757(.A(new_n957_), .ZN(new_n959_));
  NAND4_X1  g758(.A1(new_n946_), .A2(new_n919_), .A3(new_n953_), .A4(new_n959_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n958_), .A2(new_n960_), .ZN(G1354gat));
  OAI21_X1  g760(.A(G218gat), .B1(new_n947_), .B2(new_n684_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n674_), .A2(G218gat), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n946_), .A2(new_n919_), .A3(new_n963_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n962_), .A2(new_n964_), .ZN(G1355gat));
endmodule


