//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 0 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 1 0 1 0 0 1 1 0 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n685_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n796_,
    new_n797_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n963_, new_n964_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n972_, new_n973_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT23), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND3_X1  g003(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n205_));
  AND2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G169gat), .ZN(new_n207_));
  INV_X1    g006(.A(G176gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n209_), .A2(KEYINPUT24), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n209_), .A2(KEYINPUT24), .A3(new_n211_), .ZN(new_n212_));
  AND3_X1   g011(.A1(new_n206_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT26), .B(G190gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT76), .ZN(new_n215_));
  INV_X1    g014(.A(G183gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT25), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n216_), .A2(KEYINPUT25), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n214_), .B(new_n217_), .C1(new_n218_), .C2(new_n215_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n213_), .A2(new_n219_), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n204_), .B(new_n205_), .C1(G183gat), .C2(G190gat), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n221_), .A2(new_n211_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT77), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n223_), .B1(new_n207_), .B2(KEYINPUT22), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT22), .B(G169gat), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n208_), .B(new_n224_), .C1(new_n225_), .C2(new_n223_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n222_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n220_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G227gat), .A2(G233gat), .ZN(new_n229_));
  INV_X1    g028(.A(G15gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n228_), .A2(new_n231_), .ZN(new_n232_));
  AOI22_X1  g031(.A1(new_n219_), .A2(new_n213_), .B1(new_n222_), .B2(new_n226_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n231_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G71gat), .B(G99gat), .ZN(new_n236_));
  INV_X1    g035(.A(G43gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT78), .B(KEYINPUT30), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  OR3_X1    g039(.A1(new_n232_), .A2(new_n235_), .A3(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n240_), .B1(new_n232_), .B2(new_n235_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G127gat), .B(G134gat), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(G113gat), .B(G120gat), .Z(new_n245_));
  INV_X1    g044(.A(KEYINPUT80), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n244_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G113gat), .B(G120gat), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT80), .B1(new_n243_), .B2(new_n248_), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n243_), .A2(new_n248_), .A3(KEYINPUT79), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT79), .B1(new_n243_), .B2(new_n248_), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n247_), .B(new_n249_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n241_), .A2(new_n242_), .A3(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n254_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT96), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G1gat), .B(G29gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(G85gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT0), .B(G57gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(G155gat), .A2(G162gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G155gat), .A2(G162gat), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n263_), .B1(KEYINPUT1), .B2(new_n264_), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n264_), .A2(KEYINPUT1), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G141gat), .A2(G148gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(G141gat), .A2(G148gat), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n267_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n243_), .B(new_n248_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT3), .ZN(new_n274_));
  INV_X1    g073(.A(G141gat), .ZN(new_n275_));
  INV_X1    g074(.A(G148gat), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT2), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n268_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n277_), .A2(new_n279_), .A3(new_n280_), .A4(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT82), .ZN(new_n283_));
  XOR2_X1   g082(.A(G155gat), .B(G162gat), .Z(new_n284_));
  AND3_X1   g083(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n283_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n272_), .B(new_n273_), .C1(new_n285_), .C2(new_n286_), .ZN(new_n287_));
  AOI211_X1 g086(.A(new_n269_), .B(new_n270_), .C1(new_n265_), .C2(new_n266_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n282_), .A2(new_n284_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT82), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n288_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n287_), .B1(new_n292_), .B2(new_n252_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT4), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G225gat), .A2(G233gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n252_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n272_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT4), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n294_), .A2(new_n296_), .A3(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n293_), .A2(new_n295_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n262_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT93), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n304_), .A2(KEYINPUT33), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  AOI211_X1 g106(.A(new_n262_), .B(new_n305_), .C1(new_n301_), .C2(new_n302_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G8gat), .B(G36gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT18), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G64gat), .B(G92gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G226gat), .A2(G233gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT19), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT91), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT20), .ZN(new_n318_));
  INV_X1    g117(.A(G204gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(G197gat), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT85), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n319_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(KEYINPUT85), .A2(G204gat), .ZN(new_n323_));
  AOI21_X1  g122(.A(G197gat), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT86), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n320_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(G197gat), .ZN(new_n327_));
  AND2_X1   g126(.A1(KEYINPUT85), .A2(G204gat), .ZN(new_n328_));
  NOR2_X1   g127(.A1(KEYINPUT85), .A2(G204gat), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n325_), .B(new_n327_), .C1(new_n328_), .C2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT21), .B1(new_n326_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(G218gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(G211gat), .ZN(new_n334_));
  INV_X1    g133(.A(G211gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(G218gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n322_), .A2(KEYINPUT87), .A3(G197gat), .A4(new_n323_), .ZN(new_n338_));
  NOR3_X1   g137(.A1(new_n328_), .A2(new_n329_), .A3(new_n327_), .ZN(new_n339_));
  AOI21_X1  g138(.A(KEYINPUT87), .B1(new_n327_), .B2(G204gat), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n338_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT21), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n337_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n343_), .B1(new_n334_), .B2(new_n336_), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n338_), .B(new_n345_), .C1(new_n339_), .C2(new_n341_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT88), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n322_), .A2(new_n323_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n340_), .B1(new_n349_), .B2(new_n327_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n350_), .A2(KEYINPUT88), .A3(new_n338_), .A4(new_n345_), .ZN(new_n351_));
  AOI22_X1  g150(.A1(new_n332_), .A2(new_n344_), .B1(new_n348_), .B2(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n318_), .B1(new_n352_), .B2(new_n233_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n344_), .A2(new_n332_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n348_), .A2(new_n351_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n225_), .A2(new_n208_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n357_), .A2(new_n221_), .A3(new_n211_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT25), .B(G183gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n214_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n360_), .A2(new_n206_), .A3(new_n210_), .ZN(new_n361_));
  AND3_X1   g160(.A1(new_n211_), .A2(KEYINPUT92), .A3(KEYINPUT24), .ZN(new_n362_));
  INV_X1    g161(.A(new_n209_), .ZN(new_n363_));
  AOI21_X1  g162(.A(KEYINPUT92), .B1(new_n211_), .B2(KEYINPUT24), .ZN(new_n364_));
  NOR3_X1   g163(.A1(new_n362_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n358_), .B1(new_n361_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n356_), .A2(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n317_), .B1(new_n353_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n315_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n369_), .B1(new_n356_), .B2(new_n366_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT20), .B1(new_n352_), .B2(new_n233_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n313_), .B1(new_n368_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT4), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n297_), .A2(new_n298_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n374_), .B1(new_n375_), .B2(new_n287_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n295_), .B1(new_n376_), .B2(new_n299_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT94), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n293_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n375_), .A2(KEYINPUT94), .A3(new_n287_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(new_n296_), .A3(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n377_), .A2(new_n381_), .A3(new_n262_), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT20), .B1(new_n356_), .B2(new_n228_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n366_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n352_), .A2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n316_), .B1(new_n383_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n313_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n318_), .B1(new_n356_), .B2(new_n228_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n315_), .B1(new_n352_), .B2(new_n384_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n386_), .A2(new_n387_), .A3(new_n390_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n373_), .A2(new_n382_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n262_), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n376_), .A2(new_n295_), .A3(new_n299_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n302_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n393_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n301_), .A2(new_n262_), .A3(new_n302_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n353_), .A2(new_n367_), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n398_), .A2(new_n316_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n387_), .A2(KEYINPUT32), .ZN(new_n400_));
  AOI22_X1  g199(.A1(new_n396_), .A2(new_n397_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n400_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT90), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n356_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT95), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n366_), .A2(new_n405_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n358_), .B(KEYINPUT95), .C1(new_n361_), .C2(new_n365_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n352_), .A2(KEYINPUT90), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n404_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n369_), .B1(new_n411_), .B2(new_n388_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n353_), .A2(new_n317_), .A3(new_n367_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n402_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n415_));
  AOI22_X1  g214(.A1(new_n309_), .A2(new_n392_), .B1(new_n401_), .B2(new_n415_), .ZN(new_n416_));
  XOR2_X1   g215(.A(KEYINPUT83), .B(KEYINPUT28), .Z(new_n417_));
  OR3_X1    g216(.A1(new_n298_), .A2(KEYINPUT29), .A3(new_n417_), .ZN(new_n418_));
  XOR2_X1   g217(.A(G22gat), .B(G50gat), .Z(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n417_), .B1(new_n298_), .B2(KEYINPUT29), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n418_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n420_), .B1(new_n418_), .B2(new_n421_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(G78gat), .B(G106gat), .Z(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT89), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT29), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n428_), .B1(new_n292_), .B2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n298_), .A2(KEYINPUT89), .A3(KEYINPUT29), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n354_), .A2(KEYINPUT90), .A3(new_n355_), .ZN(new_n432_));
  AOI21_X1  g231(.A(KEYINPUT90), .B1(new_n354_), .B2(new_n355_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n430_), .B(new_n431_), .C1(new_n432_), .C2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(G233gat), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n435_), .A2(KEYINPUT84), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n435_), .A2(KEYINPUT84), .ZN(new_n437_));
  OAI21_X1  g236(.A(G228gat), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n434_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n298_), .A2(KEYINPUT29), .ZN(new_n441_));
  AND3_X1   g240(.A1(new_n356_), .A2(new_n438_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n427_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n444_));
  AOI211_X1 g243(.A(new_n426_), .B(new_n442_), .C1(new_n434_), .C2(new_n439_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n425_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n404_), .A2(new_n410_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n430_), .A2(new_n431_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n438_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n426_), .B1(new_n449_), .B2(new_n442_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n440_), .A2(new_n427_), .A3(new_n443_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n450_), .A2(new_n451_), .A3(new_n424_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n446_), .A2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n258_), .B1(new_n416_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT98), .ZN(new_n455_));
  NOR3_X1   g254(.A1(new_n432_), .A2(new_n433_), .A3(new_n408_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n315_), .B1(new_n456_), .B2(new_n371_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n387_), .B1(new_n457_), .B2(new_n413_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n391_), .A2(KEYINPUT27), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n455_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n313_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n461_), .A2(KEYINPUT98), .A3(KEYINPUT27), .A4(new_n391_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT97), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n301_), .A2(new_n262_), .A3(new_n302_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n464_), .B1(new_n465_), .B2(new_n303_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n396_), .A2(KEYINPUT97), .A3(new_n397_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n373_), .A2(new_n391_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT99), .B(KEYINPUT27), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n463_), .A2(new_n468_), .A3(new_n453_), .A4(new_n471_), .ZN(new_n472_));
  NOR3_X1   g271(.A1(new_n444_), .A2(new_n445_), .A3(new_n425_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n424_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n396_), .A2(new_n305_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n303_), .A2(new_n306_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n373_), .A2(new_n391_), .A3(new_n382_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n386_), .A2(new_n390_), .ZN(new_n480_));
  OAI22_X1  g279(.A1(new_n465_), .A2(new_n303_), .B1(new_n480_), .B2(new_n402_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n400_), .B1(new_n457_), .B2(new_n413_), .ZN(new_n482_));
  OAI22_X1  g281(.A1(new_n478_), .A2(new_n479_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n475_), .A2(new_n483_), .A3(KEYINPUT96), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n454_), .A2(new_n472_), .A3(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n257_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n475_), .A2(new_n463_), .A3(new_n471_), .A4(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT100), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n460_), .A2(new_n462_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT100), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n489_), .A2(new_n490_), .A3(new_n475_), .A4(new_n486_), .ZN(new_n491_));
  AOI22_X1  g290(.A1(new_n257_), .A2(new_n485_), .B1(new_n488_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT13), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G99gat), .A2(G106gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT6), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT6), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n496_), .A2(G99gat), .A3(G106gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT65), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(G99gat), .A2(G106gat), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT7), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n495_), .A2(new_n497_), .A3(KEYINPUT65), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n500_), .A2(new_n503_), .A3(new_n504_), .A4(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(G85gat), .ZN(new_n507_));
  INV_X1    g306(.A(G92gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G85gat), .A2(G92gat), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT8), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n506_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n498_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n511_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT8), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n509_), .A2(KEYINPUT9), .A3(new_n510_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n519_), .B1(KEYINPUT9), .B2(new_n510_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT10), .B(G99gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT64), .B(G106gat), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT67), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n524_), .A2(new_n525_), .A3(new_n505_), .A4(new_n500_), .ZN(new_n526_));
  OAI221_X1 g325(.A(new_n519_), .B1(KEYINPUT9), .B2(new_n510_), .C1(new_n521_), .C2(new_n522_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n500_), .A2(new_n505_), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT67), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  AOI22_X1  g328(.A1(new_n518_), .A2(KEYINPUT66), .B1(new_n526_), .B2(new_n529_), .ZN(new_n530_));
  AOI22_X1  g329(.A1(new_n506_), .A2(new_n513_), .B1(new_n516_), .B2(KEYINPUT8), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT66), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n530_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G57gat), .B(G64gat), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n535_), .A2(KEYINPUT11), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(KEYINPUT11), .ZN(new_n537_));
  XOR2_X1   g336(.A(G71gat), .B(G78gat), .Z(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  OR2_X1    g338(.A1(new_n537_), .A2(new_n538_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT12), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n527_), .A2(new_n528_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n518_), .A2(new_n546_), .A3(new_n541_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT12), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n518_), .A2(new_n546_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(new_n542_), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n534_), .A2(new_n544_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G230gat), .A2(G233gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n550_), .A2(new_n547_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n552_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G120gat), .B(G148gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G176gat), .B(G204gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n558_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n557_), .A2(new_n563_), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n565_), .A2(KEYINPUT69), .A3(new_n566_), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n558_), .A2(KEYINPUT69), .A3(new_n564_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n493_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n568_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n565_), .A2(KEYINPUT69), .A3(new_n566_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n570_), .A2(new_n571_), .A3(KEYINPUT13), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G29gat), .B(G36gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G43gat), .B(G50gat), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n575_), .B(new_n576_), .Z(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT15), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G15gat), .B(G22gat), .ZN(new_n580_));
  INV_X1    g379(.A(G1gat), .ZN(new_n581_));
  INV_X1    g380(.A(G8gat), .ZN(new_n582_));
  OAI21_X1  g381(.A(KEYINPUT14), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n580_), .A2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G1gat), .B(G8gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n579_), .A2(new_n586_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n586_), .A2(new_n577_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G229gat), .A2(G233gat), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n586_), .B(new_n577_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n589_), .ZN(new_n592_));
  AOI22_X1  g391(.A1(new_n587_), .A2(new_n590_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G113gat), .B(G141gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT74), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G169gat), .B(G197gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n593_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n593_), .A2(new_n597_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n600_), .B(KEYINPUT75), .Z(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n492_), .A2(new_n574_), .A3(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G232gat), .A2(G233gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n545_), .B1(new_n517_), .B2(new_n514_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n577_), .ZN(new_n608_));
  AOI21_X1  g407(.A(KEYINPUT71), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT71), .ZN(new_n610_));
  NOR4_X1   g409(.A1(new_n531_), .A2(new_n545_), .A3(new_n577_), .A4(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n578_), .B1(new_n530_), .B2(new_n533_), .ZN(new_n613_));
  OAI211_X1 g412(.A(KEYINPUT35), .B(new_n606_), .C1(new_n612_), .C2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n534_), .A2(new_n579_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n610_), .B1(new_n549_), .B2(new_n577_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n607_), .A2(KEYINPUT71), .A3(new_n608_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n606_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT35), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n619_), .A2(new_n620_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n615_), .A2(new_n618_), .A3(new_n622_), .A4(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n614_), .A2(new_n624_), .A3(KEYINPUT73), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G190gat), .B(G218gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT72), .ZN(new_n627_));
  XOR2_X1   g426(.A(G134gat), .B(G162gat), .Z(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n630_), .A2(KEYINPUT36), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n625_), .A2(new_n632_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n614_), .A2(new_n624_), .A3(KEYINPUT73), .A4(new_n631_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n614_), .A2(new_n624_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n636_), .A2(KEYINPUT36), .A3(new_n630_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT37), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT37), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n635_), .A2(new_n640_), .A3(new_n637_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n541_), .B(new_n586_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(G231gat), .A2(G233gat), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT17), .ZN(new_n646_));
  XOR2_X1   g445(.A(G127gat), .B(G155gat), .Z(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT16), .ZN(new_n648_));
  XNOR2_X1  g447(.A(G183gat), .B(G211gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(new_n650_));
  OR3_X1    g449(.A1(new_n645_), .A2(new_n646_), .A3(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(KEYINPUT17), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n645_), .A2(new_n652_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n642_), .A2(new_n655_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n603_), .A2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n468_), .B(KEYINPUT101), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT38), .ZN(new_n659_));
  AOI21_X1  g458(.A(G1gat), .B1(new_n659_), .B2(KEYINPUT102), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n657_), .A2(new_n658_), .A3(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n659_), .A2(KEYINPUT102), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n492_), .A2(new_n638_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n573_), .A2(new_n600_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n665_), .A2(new_n655_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n468_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n581_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT103), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n663_), .A2(new_n670_), .ZN(G1324gat));
  INV_X1    g470(.A(new_n489_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n657_), .A2(new_n582_), .A3(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n664_), .A2(new_n672_), .A3(new_n666_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n582_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT39), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n674_), .A2(KEYINPUT104), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n677_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n678_), .B1(new_n677_), .B2(new_n679_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n673_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT40), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n682_), .B(new_n683_), .ZN(G1325gat));
  INV_X1    g483(.A(new_n257_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n230_), .B1(new_n667_), .B2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT41), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n657_), .A2(new_n230_), .A3(new_n685_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1326gat));
  INV_X1    g488(.A(G22gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n690_), .B1(new_n667_), .B2(new_n453_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n691_), .B(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n657_), .A2(new_n690_), .A3(new_n453_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1327gat));
  INV_X1    g494(.A(new_n638_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n696_), .A2(new_n654_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n603_), .A2(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G29gat), .B1(new_n698_), .B2(new_n668_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT107), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n573_), .A2(new_n655_), .A3(new_n600_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n702_), .B1(new_n642_), .B2(KEYINPUT106), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n639_), .A2(new_n641_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n492_), .B2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n485_), .A2(new_n257_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n488_), .A2(new_n491_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT106), .ZN(new_n709_));
  OAI21_X1  g508(.A(KEYINPUT43), .B1(new_n704_), .B2(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n708_), .A2(new_n710_), .A3(new_n642_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n701_), .B1(new_n705_), .B2(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n700_), .B1(new_n712_), .B2(KEYINPUT44), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n710_), .B1(new_n708_), .B2(new_n642_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n492_), .A2(new_n704_), .A3(new_n703_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  OAI211_X1 g516(.A(KEYINPUT107), .B(new_n714_), .C1(new_n717_), .C2(new_n701_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n701_), .ZN(new_n719_));
  OAI211_X1 g518(.A(KEYINPUT44), .B(new_n719_), .C1(new_n715_), .C2(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT108), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT108), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n712_), .A2(new_n722_), .A3(KEYINPUT44), .ZN(new_n723_));
  AOI22_X1  g522(.A1(new_n713_), .A2(new_n718_), .B1(new_n721_), .B2(new_n723_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n658_), .A2(G29gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n699_), .B1(new_n724_), .B2(new_n725_), .ZN(G1328gat));
  INV_X1    g525(.A(KEYINPUT46), .ZN(new_n727_));
  INV_X1    g526(.A(G36gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n724_), .B2(new_n672_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n698_), .A2(new_n728_), .A3(new_n672_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT45), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n727_), .B1(new_n729_), .B2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n718_), .A2(new_n713_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n721_), .A2(new_n723_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n734_), .A2(new_n735_), .A3(new_n672_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(G36gat), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(KEYINPUT46), .A3(new_n731_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n733_), .A2(new_n738_), .ZN(G1329gat));
  NAND4_X1  g538(.A1(new_n734_), .A2(new_n735_), .A3(G43gat), .A4(new_n685_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n698_), .A2(new_n685_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(new_n237_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT47), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT47), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n740_), .A2(new_n745_), .A3(new_n742_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(G1330gat));
  INV_X1    g546(.A(G50gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n698_), .A2(new_n748_), .A3(new_n453_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT109), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n724_), .A2(new_n750_), .A3(new_n453_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(G50gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n750_), .B1(new_n724_), .B2(new_n453_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n749_), .B1(new_n752_), .B2(new_n753_), .ZN(G1331gat));
  NOR3_X1   g553(.A1(new_n492_), .A2(new_n600_), .A3(new_n573_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n656_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT110), .Z(new_n757_));
  INV_X1    g556(.A(G57gat), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n757_), .A2(new_n758_), .A3(new_n658_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n601_), .A2(new_n655_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NOR4_X1   g560(.A1(new_n492_), .A2(new_n638_), .A3(new_n573_), .A4(new_n761_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n762_), .A2(new_n668_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n759_), .B1(new_n758_), .B2(new_n763_), .ZN(G1332gat));
  INV_X1    g563(.A(G64gat), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n757_), .A2(new_n765_), .A3(new_n672_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n762_), .A2(new_n672_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(G64gat), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT48), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n766_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT111), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n770_), .B(new_n771_), .ZN(G1333gat));
  INV_X1    g571(.A(G71gat), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n757_), .A2(new_n773_), .A3(new_n685_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n773_), .B1(new_n762_), .B2(new_n685_), .ZN(new_n775_));
  XOR2_X1   g574(.A(new_n775_), .B(KEYINPUT49), .Z(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1334gat));
  INV_X1    g576(.A(G78gat), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n757_), .A2(new_n778_), .A3(new_n453_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n762_), .B2(new_n453_), .ZN(new_n780_));
  XOR2_X1   g579(.A(new_n780_), .B(KEYINPUT50), .Z(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1335gat));
  NOR3_X1   g581(.A1(new_n573_), .A2(new_n654_), .A3(new_n600_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n717_), .A2(KEYINPUT112), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n705_), .A2(new_n711_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n784_), .B1(new_n785_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(G85gat), .B1(new_n790_), .B2(new_n468_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n755_), .A2(new_n697_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n793_), .A2(new_n507_), .A3(new_n658_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n791_), .A2(new_n794_), .ZN(G1336gat));
  OAI21_X1  g594(.A(G92gat), .B1(new_n790_), .B2(new_n489_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n793_), .A2(new_n508_), .A3(new_n672_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(G1337gat));
  INV_X1    g597(.A(G99gat), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n799_), .B1(new_n789_), .B2(new_n685_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n792_), .A2(new_n521_), .A3(new_n257_), .ZN(new_n801_));
  OR3_X1    g600(.A1(new_n800_), .A2(KEYINPUT51), .A3(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(KEYINPUT51), .B1(new_n800_), .B2(new_n801_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(G1338gat));
  OR3_X1    g603(.A1(new_n792_), .A2(new_n522_), .A3(new_n475_), .ZN(new_n805_));
  INV_X1    g604(.A(G106gat), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n784_), .A2(new_n475_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n786_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n808_), .A2(new_n809_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n805_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(KEYINPUT53), .ZN(G1339gat));
  AND3_X1   g612(.A1(new_n573_), .A2(KEYINPUT113), .A3(new_n760_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT113), .B1(new_n573_), .B2(new_n760_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n704_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT54), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n818_), .B(new_n704_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n587_), .A2(new_n588_), .A3(new_n592_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n597_), .B1(new_n591_), .B2(new_n589_), .ZN(new_n822_));
  AOI22_X1  g621(.A1(new_n593_), .A2(new_n597_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n565_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n551_), .A2(KEYINPUT55), .A3(new_n552_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT115), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n551_), .A2(KEYINPUT115), .A3(KEYINPUT55), .A4(new_n552_), .ZN(new_n828_));
  XOR2_X1   g627(.A(KEYINPUT114), .B(KEYINPUT55), .Z(new_n829_));
  INV_X1    g628(.A(new_n551_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n555_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n553_), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n827_), .B(new_n828_), .C1(new_n831_), .C2(new_n832_), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n833_), .A2(KEYINPUT56), .A3(new_n563_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT56), .B1(new_n833_), .B2(new_n563_), .ZN(new_n835_));
  OAI211_X1 g634(.A(KEYINPUT58), .B(new_n824_), .C1(new_n834_), .C2(new_n835_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n836_), .A2(new_n642_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n824_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT58), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n565_), .A2(new_n600_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n570_), .A2(new_n571_), .A3(new_n823_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n638_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n837_), .A2(new_n840_), .B1(new_n845_), .B2(KEYINPUT57), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(KEYINPUT57), .B2(new_n845_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n655_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n820_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n658_), .A2(new_n685_), .A3(new_n475_), .A4(new_n489_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(KEYINPUT118), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n849_), .A2(new_n850_), .A3(new_n853_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n845_), .A2(KEYINPUT116), .A3(KEYINPUT57), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n833_), .A2(new_n563_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT56), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n833_), .A2(KEYINPUT56), .A3(new_n563_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n841_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n844_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n696_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n856_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n846_), .B1(new_n855_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n846_), .B(KEYINPUT117), .C1(new_n865_), .C2(new_n855_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n868_), .A2(new_n655_), .A3(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n852_), .B1(new_n870_), .B2(new_n820_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n854_), .B1(new_n871_), .B2(new_n850_), .ZN(new_n872_));
  OAI21_X1  g671(.A(G113gat), .B1(new_n872_), .B2(new_n602_), .ZN(new_n873_));
  INV_X1    g672(.A(G113gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n871_), .A2(new_n874_), .A3(new_n600_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n875_), .ZN(G1340gat));
  XOR2_X1   g675(.A(KEYINPUT119), .B(G120gat), .Z(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n878_), .B1(new_n872_), .B2(new_n573_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n877_), .B1(new_n573_), .B2(KEYINPUT60), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n871_), .B(new_n880_), .C1(KEYINPUT60), .C2(new_n877_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n881_), .ZN(G1341gat));
  NOR3_X1   g681(.A1(new_n820_), .A2(new_n655_), .A3(new_n852_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n884_));
  OR3_X1    g683(.A1(new_n883_), .A2(new_n884_), .A3(G127gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n883_), .B2(G127gat), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n654_), .A2(G127gat), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n854_), .B(new_n888_), .C1(new_n871_), .C2(new_n850_), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n887_), .A2(new_n889_), .ZN(G1342gat));
  NAND2_X1  g689(.A1(new_n642_), .A2(G134gat), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(KEYINPUT121), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n854_), .B(new_n892_), .C1(new_n871_), .C2(new_n850_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(G134gat), .B1(new_n871_), .B2(new_n638_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1343gat));
  NAND2_X1  g695(.A1(new_n870_), .A2(new_n820_), .ZN(new_n897_));
  AND4_X1   g696(.A1(new_n257_), .A2(new_n658_), .A3(new_n453_), .A4(new_n489_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n897_), .A2(new_n600_), .A3(new_n898_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G141gat), .ZN(G1344gat));
  XNOR2_X1  g699(.A(KEYINPUT122), .B(G148gat), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n897_), .A2(new_n898_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n901_), .B1(new_n902_), .B2(new_n574_), .ZN(new_n903_));
  AND4_X1   g702(.A1(new_n574_), .A2(new_n897_), .A3(new_n898_), .A4(new_n901_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1345gat));
  NAND3_X1  g704(.A1(new_n897_), .A2(new_n654_), .A3(new_n898_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT61), .B(G155gat), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n906_), .B(new_n907_), .ZN(G1346gat));
  NAND2_X1  g707(.A1(new_n902_), .A2(new_n638_), .ZN(new_n909_));
  INV_X1    g708(.A(G162gat), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n642_), .A2(G162gat), .ZN(new_n911_));
  XOR2_X1   g710(.A(new_n911_), .B(KEYINPUT123), .Z(new_n912_));
  AOI22_X1  g711(.A1(new_n909_), .A2(new_n910_), .B1(new_n902_), .B2(new_n912_), .ZN(G1347gat));
  AOI21_X1  g712(.A(new_n453_), .B1(new_n820_), .B2(new_n848_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n658_), .A2(new_n257_), .A3(new_n489_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n914_), .A2(new_n600_), .A3(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(G169gat), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n916_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n920_));
  INV_X1    g719(.A(new_n225_), .ZN(new_n921_));
  OAI211_X1 g720(.A(new_n919_), .B(new_n920_), .C1(new_n921_), .C2(new_n916_), .ZN(G1348gat));
  INV_X1    g721(.A(new_n915_), .ZN(new_n923_));
  AOI211_X1 g722(.A(new_n453_), .B(new_n923_), .C1(new_n820_), .C2(new_n848_), .ZN(new_n924_));
  AOI21_X1  g723(.A(G176gat), .B1(new_n924_), .B2(new_n574_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n453_), .B1(new_n870_), .B2(new_n820_), .ZN(new_n926_));
  NOR3_X1   g725(.A1(new_n923_), .A2(new_n573_), .A3(new_n208_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n925_), .B1(new_n926_), .B2(new_n927_), .ZN(G1349gat));
  NOR2_X1   g727(.A1(new_n923_), .A2(new_n655_), .ZN(new_n929_));
  AOI21_X1  g728(.A(G183gat), .B1(new_n926_), .B2(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n929_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n931_), .A2(new_n359_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n914_), .A2(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n933_), .ZN(new_n934_));
  OAI21_X1  g733(.A(KEYINPUT124), .B1(new_n930_), .B2(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT124), .ZN(new_n936_));
  AOI211_X1 g735(.A(new_n453_), .B(new_n931_), .C1(new_n870_), .C2(new_n820_), .ZN(new_n937_));
  OAI211_X1 g736(.A(new_n933_), .B(new_n936_), .C1(new_n937_), .C2(G183gat), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n935_), .A2(new_n938_), .ZN(G1350gat));
  INV_X1    g738(.A(KEYINPUT125), .ZN(new_n940_));
  INV_X1    g739(.A(G190gat), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n941_), .B1(new_n924_), .B2(new_n642_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n914_), .A2(new_n915_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n638_), .A2(new_n214_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n943_), .A2(new_n944_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n940_), .B1(new_n942_), .B2(new_n945_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n914_), .A2(new_n642_), .A3(new_n915_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(G190gat), .ZN(new_n948_));
  OAI211_X1 g747(.A(new_n948_), .B(KEYINPUT125), .C1(new_n943_), .C2(new_n944_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n946_), .A2(new_n949_), .ZN(G1351gat));
  NOR3_X1   g749(.A1(new_n475_), .A2(new_n668_), .A3(new_n685_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n951_), .A2(new_n672_), .ZN(new_n952_));
  INV_X1    g751(.A(new_n952_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n897_), .A2(new_n953_), .ZN(new_n954_));
  INV_X1    g753(.A(new_n600_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n327_), .B1(new_n954_), .B2(new_n955_), .ZN(new_n956_));
  NAND4_X1  g755(.A1(new_n897_), .A2(G197gat), .A3(new_n600_), .A4(new_n953_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n957_), .A2(KEYINPUT126), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n952_), .B1(new_n870_), .B2(new_n820_), .ZN(new_n959_));
  INV_X1    g758(.A(KEYINPUT126), .ZN(new_n960_));
  NAND4_X1  g759(.A1(new_n959_), .A2(new_n960_), .A3(G197gat), .A4(new_n600_), .ZN(new_n961_));
  AND3_X1   g760(.A1(new_n956_), .A2(new_n958_), .A3(new_n961_), .ZN(G1352gat));
  AOI21_X1  g761(.A(G204gat), .B1(new_n959_), .B2(new_n574_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n954_), .A2(new_n573_), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n963_), .B1(new_n964_), .B2(new_n349_), .ZN(G1353gat));
  NOR3_X1   g764(.A1(KEYINPUT127), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n966_));
  AOI21_X1  g765(.A(new_n966_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n959_), .A2(new_n654_), .A3(new_n967_), .ZN(new_n968_));
  OAI21_X1  g767(.A(KEYINPUT127), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n969_));
  INV_X1    g768(.A(new_n969_), .ZN(new_n970_));
  XNOR2_X1  g769(.A(new_n968_), .B(new_n970_), .ZN(G1354gat));
  OAI21_X1  g770(.A(G218gat), .B1(new_n954_), .B2(new_n704_), .ZN(new_n972_));
  NAND3_X1  g771(.A1(new_n959_), .A2(new_n333_), .A3(new_n638_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n972_), .A2(new_n973_), .ZN(G1355gat));
endmodule


