//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0' ..
//Module:
 module locked_c1355( 
    G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, G57gat,
    G64gat, G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, G113gat,
    G120gat, G127gat, G134gat, G141gat, G148gat, G155gat, G162gat, G169gat,
    G176gat, G183gat, G190gat, G197gat, G204gat, G211gat, G218gat, G225gat,
    G226gat, G227gat, G228gat, G229gat, G230gat, G231gat, G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  , KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0);
input KEYINPUT0;
input KEYINPUT1;
input KEYINPUT2;
input KEYINPUT3;
input KEYINPUT4;
input KEYINPUT5;
input KEYINPUT6;
input KEYINPUT7;
input KEYINPUT8;
input KEYINPUT9;
input KEYINPUT10;
input KEYINPUT11;
input KEYINPUT12;
input KEYINPUT13;
input KEYINPUT14;
input KEYINPUT15;
input KEYINPUT16;
input KEYINPUT17;
input KEYINPUT18;
input KEYINPUT19;
input KEYINPUT20;
input KEYINPUT21;
input KEYINPUT22;
input KEYINPUT23;
input KEYINPUT24;
input KEYINPUT25;
input KEYINPUT26;
input KEYINPUT27;
input KEYINPUT28;
input KEYINPUT29;
input KEYINPUT30;
input KEYINPUT31;
input KEYINPUT32;
input KEYINPUT33;
input KEYINPUT34;
input KEYINPUT35;
input KEYINPUT36;
input KEYINPUT37;
input KEYINPUT38;
input KEYINPUT39;
input KEYINPUT40;
input KEYINPUT41;
input KEYINPUT42;
input KEYINPUT43;
input KEYINPUT44;
input KEYINPUT45;
input KEYINPUT46;
input KEYINPUT47;
input KEYINPUT48;
input KEYINPUT49;
input KEYINPUT50;
input KEYINPUT51;
input KEYINPUT52;
input KEYINPUT53;
input KEYINPUT54;
input KEYINPUT55;
input KEYINPUT56;
input KEYINPUT57;
input KEYINPUT58;
input KEYINPUT59;
input KEYINPUT60;
input KEYINPUT61;
input KEYINPUT62;
input KEYINPUT63;
//Header:
   input  G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat,
    G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat, G106gat,
    G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat, G162gat,
    G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat, G218gat,
    G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat, G232gat,
    G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_, new_n80_,
    new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_, new_n87_,
    new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_,
    new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_, new_n101_,
    new_n102_, new_n103_, new_n104_, new_n105_, new_n106_, new_n107_,
    new_n108_, new_n109_, new_n110_, new_n111_, new_n112_, new_n113_,
    new_n114_, new_n115_, new_n116_, new_n117_, new_n118_, new_n119_,
    new_n120_, new_n121_, new_n122_, new_n123_, new_n124_, new_n125_,
    new_n126_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_,
    new_n132_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_,
    new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n325_, new_n326_, new_n327_, new_n329_, new_n330_, new_n332_,
    new_n333_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n342_, new_n343_, new_n344_, new_n346_, new_n347_,
    new_n349_, new_n350_, new_n352_, new_n353_, new_n354_, new_n355_,
    new_n356_, new_n358_, new_n359_, new_n361_, new_n362_, new_n364_,
    new_n365_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n373_, new_n374_, new_n375_, new_n377_, new_n378_, new_n380_,
    new_n381_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n406_,
    new_n407_, new_n408_, new_n410_, new_n411_, new_n413_, new_n414_,
    new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n422_,
    new_n423_, new_n425_, new_n426_, new_n428_, new_n429_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n436_, new_n437_, new_n439_,
    new_n440_, new_n442_, new_n443_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n450_, new_n451_, new_n453_, new_n454_, new_n456_,
    new_n457_;
wire RLL_wire_A_0;
wire RLL_wire_A_1;
wire RLL_wire_A_2;
wire RLL_wire_A_3;
wire RLL_wire_A_4;
wire RLL_wire_A_5;
wire RLL_wire_A_6;
wire RLL_wire_A_7;
wire RLL_wire_A_8;
wire RLL_wire_A_9;
wire RLL_wire_A_10;
wire RLL_wire_A_11;
wire RLL_wire_A_12;
wire RLL_wire_A_13;
wire RLL_wire_A_14;
wire RLL_wire_A_15;
wire RLL_wire_A_16;
wire RLL_wire_A_17;
wire RLL_wire_A_18;
wire RLL_wire_A_19;
wire RLL_wire_A_20;
wire RLL_wire_A_21;
wire RLL_wire_A_22;
wire RLL_wire_A_23;
wire RLL_wire_A_24;
wire RLL_wire_A_25;
wire RLL_wire_A_26;
wire RLL_wire_A_27;
wire RLL_wire_A_28;
wire RLL_wire_A_29;
wire RLL_wire_A_30;
wire RLL_wire_A_31;
wire RLL_wire_A_32;
wire RLL_wire_A_33;
wire RLL_wire_A_34;
wire RLL_wire_A_35;
wire RLL_wire_A_36;
wire RLL_wire_A_37;
wire RLL_wire_A_38;
wire RLL_wire_A_39;
wire RLL_wire_A_40;
wire RLL_wire_A_41;
wire RLL_wire_A_42;
wire RLL_wire_A_43;
wire RLL_wire_A_44;
wire RLL_wire_A_45;
wire RLL_wire_A_46;
wire RLL_wire_A_47;
wire RLL_wire_A_48;
wire RLL_wire_A_49;
wire RLL_wire_A_50;
wire RLL_wire_A_51;
wire RLL_wire_A_52;
wire RLL_wire_A_53;
wire RLL_wire_A_54;
wire RLL_wire_A_55;
wire RLL_wire_A_56;
wire RLL_wire_A_57;
wire RLL_wire_A_58;
wire RLL_wire_A_59;
wire RLL_wire_A_60;
wire RLL_wire_A_61;
wire RLL_wire_A_62;
wire RLL_wire_A_63;

//Body:
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(RLL_wire_A_0));
  XNOR2_X1 RLL_XNOR_0 (.A(RLL_wire_A_0), .B(KEYINPUT0), .ZN(new_n74_) );
  XNOR2_X1  g001(.A(G57gat), .B(G85gat), .ZN(new_n75_));
  XNOR2_X1  g002(.A(new_n74_), .B(new_n75_), .ZN(new_n76_));
  INV_X1    g003(.A(new_n76_), .ZN(new_n77_));
  NAND2_X1  g004(.A1(G225gat), .A2(G233gat), .ZN(new_n78_));
  INV_X1    g005(.A(new_n78_), .ZN(new_n79_));
  AND2_X1   g006(.A1(G113gat), .A2(G120gat), .ZN(new_n80_));
  NOR2_X1   g007(.A1(G113gat), .A2(G120gat), .ZN(new_n81_));
  NOR2_X1   g008(.A1(new_n80_), .A2(new_n81_), .ZN(new_n82_));
  NAND2_X1  g009(.A1(G127gat), .A2(G134gat), .ZN(new_n83_));
  INV_X1    g010(.A(G127gat), .ZN(new_n84_));
  INV_X1    g011(.A(G134gat), .ZN(new_n85_));
  NAND2_X1  g012(.A1(new_n84_), .A2(new_n85_), .ZN(new_n86_));
  NAND2_X1  g013(.A1(new_n86_), .A2(new_n83_), .ZN(new_n87_));
  NAND2_X1  g014(.A1(new_n87_), .A2(new_n82_), .ZN(new_n88_));
  OAI211_X1 g015(.A(new_n86_), .B(new_n83_), .C1(new_n80_), .C2(new_n81_), .ZN(new_n89_));
  NAND2_X1  g016(.A1(G141gat), .A2(G148gat), .ZN(new_n90_));
  INV_X1    g017(.A(G141gat), .ZN(new_n91_));
  INV_X1    g018(.A(G148gat), .ZN(new_n92_));
  NAND2_X1  g019(.A1(new_n91_), .A2(new_n92_), .ZN(new_n93_));
  NAND2_X1  g020(.A1(G155gat), .A2(G162gat), .ZN(new_n94_));
  INV_X1    g021(.A(new_n94_), .ZN(RLL_wire_A_1));
  XOR2_X1 RLL_XOR_1 (.A(RLL_wire_A_1), .B(KEYINPUT1), .Z(new_n95_) );
  NOR2_X1   g022(.A1(G155gat), .A2(G162gat), .ZN(new_n96_));
  OAI211_X1 g023(.A(new_n93_), .B(new_n90_), .C1(new_n95_), .C2(new_n96_), .ZN(new_n97_));
  AND2_X1   g024(.A1(G141gat), .A2(G148gat), .ZN(RLL_wire_A_2));
  XNOR2_X1 RLL_XNOR_2 (.A(RLL_wire_A_2), .B(KEYINPUT2), .ZN(new_n98_) );
  NOR2_X1   g025(.A1(G141gat), .A2(G148gat), .ZN(RLL_wire_A_3));
  XOR2_X1 RLL_XOR_3 (.A(RLL_wire_A_3), .B(KEYINPUT3), .Z(new_n99_) );
  INV_X1    g026(.A(G155gat), .ZN(new_n100_));
  INV_X1    g027(.A(G162gat), .ZN(new_n101_));
  NAND2_X1  g028(.A1(new_n100_), .A2(new_n101_), .ZN(new_n102_));
  OAI211_X1 g029(.A(new_n102_), .B(new_n94_), .C1(new_n98_), .C2(new_n99_), .ZN(new_n103_));
  AOI22_X1  g030(.A1(new_n88_), .A2(new_n89_), .B1(new_n97_), .B2(new_n103_), .ZN(RLL_wire_A_4));
  XNOR2_X1 RLL_XNOR_4 (.A(RLL_wire_A_4), .B(KEYINPUT4), .ZN(new_n104_) );
  AND4_X1   g031(.A1(new_n88_), .A2(new_n89_), .A3(new_n97_), .A4(new_n103_), .ZN(new_n105_));
  OAI21_X1  g032(.A(new_n79_), .B1(new_n105_), .B2(new_n104_), .ZN(new_n106_));
  NAND2_X1  g033(.A1(new_n88_), .A2(new_n89_), .ZN(new_n107_));
  NAND2_X1  g034(.A1(new_n97_), .A2(new_n103_), .ZN(new_n108_));
  NAND2_X1  g035(.A1(new_n107_), .A2(new_n108_), .ZN(new_n109_));
  NAND4_X1  g036(.A1(new_n88_), .A2(new_n89_), .A3(new_n97_), .A4(new_n103_), .ZN(new_n110_));
  NAND3_X1  g037(.A1(new_n109_), .A2(new_n78_), .A3(new_n110_), .ZN(new_n111_));
  AND3_X1   g038(.A1(new_n106_), .A2(new_n77_), .A3(new_n111_), .ZN(new_n112_));
  AOI21_X1  g039(.A(new_n77_), .B1(new_n106_), .B2(new_n111_), .ZN(new_n113_));
  NOR2_X1   g040(.A1(new_n112_), .A2(new_n113_), .ZN(new_n114_));
  XNOR2_X1  g041(.A(G120gat), .B(G148gat), .ZN(new_n115_));
  XNOR2_X1  g042(.A(G176gat), .B(G204gat), .ZN(RLL_wire_A_5));
  XOR2_X1 RLL_XOR_5 (.A(RLL_wire_A_5), .B(KEYINPUT5), .Z(new_n116_) );
  XNOR2_X1  g043(.A(new_n115_), .B(new_n116_), .ZN(new_n117_));
  INV_X1    g044(.A(new_n117_), .ZN(new_n118_));
  NAND2_X1  g045(.A1(G230gat), .A2(G233gat), .ZN(new_n119_));
  INV_X1    g046(.A(new_n119_), .ZN(new_n120_));
  NAND2_X1  g047(.A1(G85gat), .A2(G92gat), .ZN(new_n121_));
  NOR2_X1   g048(.A1(G85gat), .A2(G92gat), .ZN(new_n122_));
  INV_X1    g049(.A(new_n122_), .ZN(new_n123_));
  NAND2_X1  g050(.A1(G99gat), .A2(G106gat), .ZN(RLL_wire_A_6));
  XNOR2_X1 RLL_XNOR_6 (.A(RLL_wire_A_6), .B(KEYINPUT6), .ZN(new_n124_) );
  INV_X1    g051(.A(new_n124_), .ZN(new_n125_));
  NOR2_X1   g052(.A1(G99gat), .A2(G106gat), .ZN(RLL_wire_A_7));
  XOR2_X1 RLL_XOR_7 (.A(RLL_wire_A_7), .B(KEYINPUT7), .Z(new_n126_) );
  OAI211_X1 g053(.A(new_n123_), .B(new_n121_), .C1(new_n125_), .C2(new_n126_), .ZN(RLL_wire_A_8));
  XNOR2_X1 RLL_XNOR_8 (.A(RLL_wire_A_8), .B(KEYINPUT8), .ZN(new_n127_) );
  INV_X1    g054(.A(new_n121_), .ZN(RLL_wire_A_9));
  XNOR2_X1 RLL_XNOR_9 (.A(RLL_wire_A_9), .B(KEYINPUT9), .ZN(new_n128_) );
  INV_X1    g055(.A(G99gat), .ZN(RLL_wire_A_10));
  XNOR2_X1 RLL_XNOR_10 (.A(RLL_wire_A_10), .B(KEYINPUT10), .ZN(new_n129_) );
  INV_X1    g056(.A(G106gat), .ZN(new_n130_));
  NAND2_X1  g057(.A1(new_n129_), .A2(new_n130_), .ZN(new_n131_));
  OAI211_X1 g058(.A(new_n131_), .B(new_n124_), .C1(new_n128_), .C2(new_n122_), .ZN(new_n132_));
  NAND2_X1  g059(.A1(G57gat), .A2(G64gat), .ZN(new_n133_));
  INV_X1    g060(.A(G57gat), .ZN(new_n134_));
  INV_X1    g061(.A(G64gat), .ZN(new_n135_));
  NAND2_X1  g062(.A1(new_n134_), .A2(new_n135_), .ZN(new_n136_));
  NAND2_X1  g063(.A1(G71gat), .A2(G78gat), .ZN(new_n137_));
  INV_X1    g064(.A(new_n137_), .ZN(new_n138_));
  NOR2_X1   g065(.A1(G71gat), .A2(G78gat), .ZN(new_n139_));
  OAI211_X1 g066(.A(new_n136_), .B(new_n133_), .C1(new_n138_), .C2(new_n139_), .ZN(new_n140_));
  AND2_X1   g067(.A1(G57gat), .A2(G64gat), .ZN(new_n141_));
  NOR2_X1   g068(.A1(G57gat), .A2(G64gat), .ZN(new_n142_));
  INV_X1    g069(.A(G71gat), .ZN(new_n143_));
  INV_X1    g070(.A(G78gat), .ZN(new_n144_));
  NAND2_X1  g071(.A1(new_n143_), .A2(new_n144_), .ZN(new_n145_));
  OAI211_X1 g072(.A(new_n145_), .B(new_n137_), .C1(new_n141_), .C2(new_n142_), .ZN(RLL_wire_A_11));
  XNOR2_X1 RLL_XNOR_11 (.A(RLL_wire_A_11), .B(KEYINPUT11), .ZN(new_n146_) );
  AOI22_X1  g073(.A1(new_n127_), .A2(new_n132_), .B1(new_n140_), .B2(new_n146_), .ZN(new_n147_));
  AND4_X1   g074(.A1(new_n127_), .A2(new_n132_), .A3(new_n140_), .A4(new_n146_), .ZN(new_n148_));
  OAI21_X1  g075(.A(new_n120_), .B1(new_n148_), .B2(new_n147_), .ZN(new_n149_));
  NAND2_X1  g076(.A1(new_n127_), .A2(new_n132_), .ZN(new_n150_));
  NAND2_X1  g077(.A1(new_n140_), .A2(new_n146_), .ZN(new_n151_));
  NAND2_X1  g078(.A1(new_n150_), .A2(new_n151_), .ZN(RLL_wire_A_12));
  XNOR2_X1 RLL_XNOR_12 (.A(RLL_wire_A_12), .B(KEYINPUT12), .ZN(new_n152_) );
  NAND4_X1  g079(.A1(new_n127_), .A2(new_n132_), .A3(new_n140_), .A4(new_n146_), .ZN(new_n153_));
  NAND3_X1  g080(.A1(new_n152_), .A2(new_n119_), .A3(new_n153_), .ZN(new_n154_));
  AND3_X1   g081(.A1(new_n149_), .A2(new_n118_), .A3(new_n154_), .ZN(new_n155_));
  AOI21_X1  g082(.A(new_n118_), .B1(new_n149_), .B2(new_n154_), .ZN(new_n156_));
  NOR2_X1   g083(.A1(new_n155_), .A2(new_n156_), .ZN(RLL_wire_A_13));
  XOR2_X1 RLL_XOR_13 (.A(RLL_wire_A_13), .B(KEYINPUT13), .Z(new_n157_) );
  XNOR2_X1  g084(.A(G113gat), .B(G141gat), .ZN(new_n158_));
  XNOR2_X1  g085(.A(G169gat), .B(G197gat), .ZN(new_n159_));
  XNOR2_X1  g086(.A(new_n158_), .B(new_n159_), .ZN(new_n160_));
  INV_X1    g087(.A(new_n160_), .ZN(new_n161_));
  NAND2_X1  g088(.A1(G229gat), .A2(G233gat), .ZN(new_n162_));
  INV_X1    g089(.A(new_n162_), .ZN(new_n163_));
  AND2_X1   g090(.A1(G29gat), .A2(G36gat), .ZN(new_n164_));
  NOR2_X1   g091(.A1(G29gat), .A2(G36gat), .ZN(new_n165_));
  NOR2_X1   g092(.A1(new_n164_), .A2(new_n165_), .ZN(new_n166_));
  NAND2_X1  g093(.A1(G43gat), .A2(G50gat), .ZN(new_n167_));
  INV_X1    g094(.A(G43gat), .ZN(new_n168_));
  INV_X1    g095(.A(G50gat), .ZN(new_n169_));
  NAND2_X1  g096(.A1(new_n168_), .A2(new_n169_), .ZN(new_n170_));
  NAND2_X1  g097(.A1(new_n170_), .A2(new_n167_), .ZN(new_n171_));
  NAND2_X1  g098(.A1(new_n171_), .A2(new_n166_), .ZN(new_n172_));
  OAI211_X1 g099(.A(new_n170_), .B(new_n167_), .C1(new_n164_), .C2(new_n165_), .ZN(new_n173_));
  NAND2_X1  g100(.A1(G1gat), .A2(G8gat), .ZN(new_n174_));
  INV_X1    g101(.A(G1gat), .ZN(new_n175_));
  INV_X1    g102(.A(G8gat), .ZN(new_n176_));
  NAND2_X1  g103(.A1(new_n175_), .A2(new_n176_), .ZN(RLL_wire_A_14));
  XOR2_X1 RLL_XOR_14 (.A(RLL_wire_A_14), .B(KEYINPUT14), .Z(new_n177_) );
  NAND2_X1  g104(.A1(G15gat), .A2(G22gat), .ZN(new_n178_));
  INV_X1    g105(.A(new_n178_), .ZN(new_n179_));
  NOR2_X1   g106(.A1(G15gat), .A2(G22gat), .ZN(new_n180_));
  OAI211_X1 g107(.A(new_n177_), .B(new_n174_), .C1(new_n179_), .C2(new_n180_), .ZN(new_n181_));
  AND2_X1   g108(.A1(G1gat), .A2(G8gat), .ZN(new_n182_));
  NOR2_X1   g109(.A1(G1gat), .A2(G8gat), .ZN(new_n183_));
  INV_X1    g110(.A(G15gat), .ZN(new_n184_));
  INV_X1    g111(.A(G22gat), .ZN(new_n185_));
  NAND2_X1  g112(.A1(new_n184_), .A2(new_n185_), .ZN(new_n186_));
  OAI211_X1 g113(.A(new_n186_), .B(new_n178_), .C1(new_n182_), .C2(new_n183_), .ZN(new_n187_));
  AOI22_X1  g114(.A1(new_n172_), .A2(new_n173_), .B1(new_n181_), .B2(new_n187_), .ZN(new_n188_));
  AND4_X1   g115(.A1(new_n172_), .A2(new_n173_), .A3(new_n181_), .A4(new_n187_), .ZN(new_n189_));
  OAI21_X1  g116(.A(new_n163_), .B1(new_n189_), .B2(new_n188_), .ZN(new_n190_));
  NAND2_X1  g117(.A1(new_n172_), .A2(new_n173_), .ZN(RLL_wire_A_15));
  XOR2_X1 RLL_XOR_15 (.A(RLL_wire_A_15), .B(KEYINPUT15), .Z(new_n191_) );
  NAND2_X1  g118(.A1(new_n181_), .A2(new_n187_), .ZN(new_n192_));
  NAND2_X1  g119(.A1(new_n191_), .A2(new_n192_), .ZN(new_n193_));
  NAND4_X1  g120(.A1(new_n172_), .A2(new_n173_), .A3(new_n181_), .A4(new_n187_), .ZN(new_n194_));
  NAND3_X1  g121(.A1(new_n193_), .A2(new_n162_), .A3(new_n194_), .ZN(new_n195_));
  AND3_X1   g122(.A1(new_n190_), .A2(new_n161_), .A3(new_n195_), .ZN(new_n196_));
  AOI21_X1  g123(.A(new_n161_), .B1(new_n190_), .B2(new_n195_), .ZN(new_n197_));
  NOR2_X1   g124(.A1(new_n196_), .A2(new_n197_), .ZN(new_n198_));
  INV_X1    g125(.A(new_n198_), .ZN(new_n199_));
  XOR2_X1   g126(.A(G127gat), .B(G155gat), .Z(new_n200_));
  XNOR2_X1  g127(.A(G183gat), .B(G211gat), .ZN(new_n201_));
  XOR2_X1   g128(.A(new_n200_), .B(new_n201_), .Z(new_n202_));
  INV_X1    g129(.A(new_n202_), .ZN(RLL_wire_A_16));
  XNOR2_X1 RLL_XNOR_16 (.A(RLL_wire_A_16), .B(KEYINPUT16), .ZN(new_n203_) );
  AND2_X1   g130(.A1(G231gat), .A2(G233gat), .ZN(new_n204_));
  NAND2_X1  g131(.A1(new_n151_), .A2(new_n192_), .ZN(new_n205_));
  NAND4_X1  g132(.A1(new_n140_), .A2(new_n146_), .A3(new_n181_), .A4(new_n187_), .ZN(new_n206_));
  NAND2_X1  g133(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g134(.A1(new_n207_), .A2(new_n204_), .ZN(new_n208_));
  NOR2_X1   g135(.A1(new_n207_), .A2(new_n204_), .ZN(new_n209_));
  INV_X1    g136(.A(new_n209_), .ZN(new_n210_));
  AND3_X1   g137(.A1(new_n210_), .A2(new_n203_), .A3(new_n208_), .ZN(new_n211_));
  AOI21_X1  g138(.A(new_n203_), .B1(new_n210_), .B2(new_n208_), .ZN(RLL_wire_A_17));
  XNOR2_X1 RLL_XNOR_17 (.A(RLL_wire_A_17), .B(KEYINPUT17), .ZN(new_n212_) );
  NOR2_X1   g139(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g140(.A(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g141(.A(G8gat), .B(G36gat), .ZN(RLL_wire_A_18));
  XOR2_X1 RLL_XOR_18 (.A(RLL_wire_A_18), .B(KEYINPUT18), .Z(new_n215_) );
  XNOR2_X1  g142(.A(G64gat), .B(G92gat), .ZN(new_n216_));
  XNOR2_X1  g143(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  INV_X1    g144(.A(new_n217_), .ZN(new_n218_));
  NAND2_X1  g145(.A1(G226gat), .A2(G233gat), .ZN(RLL_wire_A_19));
  XNOR2_X1 RLL_XNOR_19 (.A(RLL_wire_A_19), .B(KEYINPUT19), .ZN(new_n219_) );
  INV_X1    g146(.A(new_n219_), .ZN(RLL_wire_A_20));
  XNOR2_X1 RLL_XNOR_20 (.A(RLL_wire_A_20), .B(KEYINPUT20), .ZN(new_n220_) );
  NAND2_X1  g147(.A1(G197gat), .A2(G204gat), .ZN(new_n221_));
  INV_X1    g148(.A(G197gat), .ZN(new_n222_));
  INV_X1    g149(.A(G204gat), .ZN(new_n223_));
  NAND2_X1  g150(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g151(.A1(G211gat), .A2(G218gat), .ZN(new_n225_));
  INV_X1    g152(.A(new_n225_), .ZN(new_n226_));
  NOR2_X1   g153(.A1(G211gat), .A2(G218gat), .ZN(new_n227_));
  OAI211_X1 g154(.A(new_n224_), .B(new_n221_), .C1(new_n226_), .C2(new_n227_), .ZN(RLL_wire_A_21));
  XNOR2_X1 RLL_XNOR_21 (.A(RLL_wire_A_21), .B(KEYINPUT21), .ZN(new_n228_) );
  INV_X1    g155(.A(new_n221_), .ZN(new_n229_));
  NOR2_X1   g156(.A1(G197gat), .A2(G204gat), .ZN(new_n230_));
  INV_X1    g157(.A(G211gat), .ZN(new_n231_));
  INV_X1    g158(.A(G218gat), .ZN(new_n232_));
  NAND2_X1  g159(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  OAI211_X1 g160(.A(new_n233_), .B(new_n225_), .C1(new_n229_), .C2(new_n230_), .ZN(new_n234_));
  NAND2_X1  g161(.A1(G169gat), .A2(G176gat), .ZN(new_n235_));
  INV_X1    g162(.A(G169gat), .ZN(RLL_wire_A_22));
  XOR2_X1 RLL_XOR_22 (.A(RLL_wire_A_22), .B(KEYINPUT22), .Z(new_n236_) );
  INV_X1    g163(.A(G176gat), .ZN(new_n237_));
  NAND2_X1  g164(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g165(.A1(G183gat), .A2(G190gat), .ZN(RLL_wire_A_23));
  XNOR2_X1 RLL_XNOR_23 (.A(RLL_wire_A_23), .B(KEYINPUT23), .ZN(new_n239_) );
  INV_X1    g166(.A(new_n239_), .ZN(new_n240_));
  NOR2_X1   g167(.A1(G183gat), .A2(G190gat), .ZN(new_n241_));
  OAI211_X1 g168(.A(new_n238_), .B(new_n235_), .C1(new_n240_), .C2(new_n241_), .ZN(new_n242_));
  AND2_X1   g169(.A1(G169gat), .A2(G176gat), .ZN(new_n243_));
  NOR2_X1   g170(.A1(G169gat), .A2(G176gat), .ZN(RLL_wire_A_24));
  XNOR2_X1 RLL_XNOR_24 (.A(RLL_wire_A_24), .B(KEYINPUT24), .ZN(new_n244_) );
  INV_X1    g171(.A(G183gat), .ZN(RLL_wire_A_25));
  XOR2_X1 RLL_XOR_25 (.A(RLL_wire_A_25), .B(KEYINPUT25), .Z(new_n245_) );
  INV_X1    g172(.A(G190gat), .ZN(RLL_wire_A_26));
  XOR2_X1 RLL_XOR_26 (.A(RLL_wire_A_26), .B(KEYINPUT26), .Z(new_n246_) );
  NAND2_X1  g173(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  OAI211_X1 g174(.A(new_n247_), .B(new_n239_), .C1(new_n243_), .C2(new_n244_), .ZN(new_n248_));
  AOI22_X1  g175(.A1(new_n228_), .A2(new_n234_), .B1(new_n242_), .B2(new_n248_), .ZN(new_n249_));
  AND4_X1   g176(.A1(new_n228_), .A2(new_n234_), .A3(new_n242_), .A4(new_n248_), .ZN(new_n250_));
  OAI21_X1  g177(.A(new_n220_), .B1(new_n250_), .B2(new_n249_), .ZN(new_n251_));
  NAND2_X1  g178(.A1(new_n228_), .A2(new_n234_), .ZN(new_n252_));
  NAND2_X1  g179(.A1(new_n242_), .A2(new_n248_), .ZN(new_n253_));
  NAND2_X1  g180(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND4_X1  g181(.A1(new_n228_), .A2(new_n234_), .A3(new_n242_), .A4(new_n248_), .ZN(new_n255_));
  NAND3_X1  g182(.A1(new_n254_), .A2(new_n219_), .A3(new_n255_), .ZN(new_n256_));
  AND3_X1   g183(.A1(new_n251_), .A2(new_n218_), .A3(new_n256_), .ZN(new_n257_));
  AOI21_X1  g184(.A(new_n218_), .B1(new_n251_), .B2(new_n256_), .ZN(new_n258_));
  NOR2_X1   g185(.A1(new_n257_), .A2(new_n258_), .ZN(RLL_wire_A_27));
  XNOR2_X1 RLL_XNOR_27 (.A(RLL_wire_A_27), .B(KEYINPUT27), .ZN(new_n259_) );
  XNOR2_X1  g186(.A(G22gat), .B(G50gat), .ZN(new_n260_));
  XNOR2_X1  g187(.A(G78gat), .B(G106gat), .ZN(RLL_wire_A_28));
  XOR2_X1 RLL_XOR_28 (.A(RLL_wire_A_28), .B(KEYINPUT28), .Z(new_n261_) );
  XNOR2_X1  g188(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  INV_X1    g189(.A(new_n262_), .ZN(new_n263_));
  NAND2_X1  g190(.A1(G228gat), .A2(G233gat), .ZN(new_n264_));
  NAND2_X1  g191(.A1(new_n252_), .A2(new_n108_), .ZN(new_n265_));
  NAND4_X1  g192(.A1(new_n97_), .A2(new_n228_), .A3(new_n234_), .A4(new_n103_), .ZN(RLL_wire_A_29));
  XOR2_X1 RLL_XOR_29 (.A(RLL_wire_A_29), .B(KEYINPUT29), .Z(new_n266_) );
  AOI21_X1  g193(.A(new_n264_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g194(.A(new_n267_), .ZN(new_n268_));
  NAND3_X1  g195(.A1(new_n265_), .A2(new_n264_), .A3(new_n266_), .ZN(new_n269_));
  NAND3_X1  g196(.A1(new_n268_), .A2(new_n263_), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g197(.A(new_n269_), .ZN(new_n271_));
  OAI21_X1  g198(.A(new_n262_), .B1(new_n271_), .B2(new_n267_), .ZN(new_n272_));
  NAND2_X1  g199(.A1(new_n272_), .A2(new_n270_), .ZN(new_n273_));
  INV_X1    g200(.A(new_n273_), .ZN(new_n274_));
  XOR2_X1   g201(.A(G15gat), .B(G43gat), .Z(new_n275_));
  XNOR2_X1  g202(.A(G71gat), .B(G99gat), .ZN(new_n276_));
  XOR2_X1   g203(.A(new_n275_), .B(new_n276_), .Z(new_n277_));
  INV_X1    g204(.A(new_n277_), .ZN(new_n278_));
  AND2_X1   g205(.A1(G227gat), .A2(G233gat), .ZN(RLL_wire_A_30));
  XOR2_X1 RLL_XOR_30 (.A(RLL_wire_A_30), .B(KEYINPUT30), .Z(new_n279_) );
  XNOR2_X1  g206(.A(new_n107_), .B(new_n253_), .ZN(new_n280_));
  NAND2_X1  g207(.A1(new_n280_), .A2(new_n279_), .ZN(new_n281_));
  NOR2_X1   g208(.A1(new_n280_), .A2(new_n279_), .ZN(new_n282_));
  INV_X1    g209(.A(new_n282_), .ZN(new_n283_));
  NAND3_X1  g210(.A1(new_n283_), .A2(new_n278_), .A3(new_n281_), .ZN(new_n284_));
  INV_X1    g211(.A(new_n281_), .ZN(new_n285_));
  OAI21_X1  g212(.A(new_n277_), .B1(new_n285_), .B2(new_n282_), .ZN(new_n286_));
  NAND2_X1  g213(.A1(new_n286_), .A2(new_n284_), .ZN(RLL_wire_A_31));
  XNOR2_X1 RLL_XNOR_31 (.A(RLL_wire_A_31), .B(KEYINPUT31), .ZN(new_n287_) );
  NAND4_X1  g214(.A1(new_n287_), .A2(new_n114_), .A3(new_n259_), .A4(new_n274_), .ZN(new_n288_));
  INV_X1    g215(.A(new_n287_), .ZN(new_n289_));
  NAND3_X1  g216(.A1(new_n251_), .A2(new_n218_), .A3(new_n256_), .ZN(new_n290_));
  NAND2_X1  g217(.A1(new_n251_), .A2(new_n256_), .ZN(RLL_wire_A_32));
  XNOR2_X1 RLL_XNOR_32 (.A(RLL_wire_A_32), .B(KEYINPUT32), .ZN(new_n291_) );
  NAND2_X1  g218(.A1(new_n291_), .A2(new_n217_), .ZN(new_n292_));
  OAI211_X1 g219(.A(new_n292_), .B(new_n290_), .C1(new_n112_), .C2(new_n113_), .ZN(new_n293_));
  NAND3_X1  g220(.A1(new_n106_), .A2(new_n77_), .A3(new_n111_), .ZN(RLL_wire_A_33));
  XNOR2_X1 RLL_XNOR_33 (.A(RLL_wire_A_33), .B(KEYINPUT33), .ZN(new_n294_) );
  AOI21_X1  g221(.A(new_n78_), .B1(new_n109_), .B2(new_n110_), .ZN(new_n295_));
  NOR3_X1   g222(.A1(new_n105_), .A2(new_n104_), .A3(new_n79_), .ZN(new_n296_));
  OAI21_X1  g223(.A(new_n76_), .B1(new_n296_), .B2(new_n295_), .ZN(new_n297_));
  OAI211_X1 g224(.A(new_n294_), .B(new_n297_), .C1(new_n257_), .C2(new_n258_), .ZN(new_n298_));
  AOI21_X1  g225(.A(new_n273_), .B1(new_n293_), .B2(new_n298_), .ZN(new_n299_));
  AND3_X1   g226(.A1(new_n114_), .A2(new_n259_), .A3(new_n273_), .ZN(new_n300_));
  OAI21_X1  g227(.A(new_n289_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g228(.A(G134gat), .B(G162gat), .ZN(new_n302_));
  XNOR2_X1  g229(.A(G190gat), .B(G218gat), .ZN(new_n303_));
  XNOR2_X1  g230(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  INV_X1    g231(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g232(.A1(G232gat), .A2(G233gat), .ZN(RLL_wire_A_34));
  XNOR2_X1 RLL_XNOR_34 (.A(RLL_wire_A_34), .B(KEYINPUT34), .ZN(new_n306_) );
  NAND2_X1  g233(.A1(new_n191_), .A2(new_n150_), .ZN(new_n307_));
  NAND4_X1  g234(.A1(new_n172_), .A2(new_n127_), .A3(new_n132_), .A4(new_n173_), .ZN(new_n308_));
  AOI21_X1  g235(.A(new_n306_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g236(.A(new_n309_), .ZN(new_n310_));
  NAND3_X1  g237(.A1(new_n307_), .A2(new_n306_), .A3(new_n308_), .ZN(RLL_wire_A_35));
  XNOR2_X1 RLL_XNOR_35 (.A(RLL_wire_A_35), .B(KEYINPUT35), .ZN(new_n311_) );
  NAND3_X1  g238(.A1(new_n310_), .A2(new_n305_), .A3(new_n311_), .ZN(RLL_wire_A_36));
  XOR2_X1 RLL_XOR_36 (.A(RLL_wire_A_36), .B(KEYINPUT36), .Z(new_n312_) );
  INV_X1    g239(.A(new_n311_), .ZN(new_n313_));
  OAI21_X1  g240(.A(new_n304_), .B1(new_n313_), .B2(new_n309_), .ZN(new_n314_));
  NAND2_X1  g241(.A1(new_n314_), .A2(new_n312_), .ZN(new_n315_));
  AOI21_X1  g242(.A(new_n315_), .B1(new_n301_), .B2(new_n288_), .ZN(new_n316_));
  NAND4_X1  g243(.A1(new_n316_), .A2(new_n157_), .A3(new_n199_), .A4(new_n214_), .ZN(new_n317_));
  OAI21_X1  g244(.A(G1gat), .B1(new_n317_), .B2(new_n114_), .ZN(new_n318_));
  INV_X1    g245(.A(new_n114_), .ZN(new_n319_));
  NAND2_X1  g246(.A1(new_n301_), .A2(new_n288_), .ZN(new_n320_));
  AND2_X1   g247(.A1(new_n314_), .A2(new_n312_), .ZN(RLL_wire_A_37));
  XNOR2_X1 RLL_XNOR_37 (.A(RLL_wire_A_37), .B(KEYINPUT37), .ZN(new_n321_) );
  AND4_X1   g248(.A1(new_n199_), .A2(new_n320_), .A3(new_n214_), .A4(new_n321_), .ZN(new_n322_));
  NAND4_X1  g249(.A1(new_n322_), .A2(new_n175_), .A3(new_n319_), .A4(new_n157_), .ZN(RLL_wire_A_38));
  XNOR2_X1 RLL_XNOR_38 (.A(RLL_wire_A_38), .B(KEYINPUT38), .ZN(new_n323_) );
  NAND2_X1  g250(.A1(new_n323_), .A2(new_n318_), .ZN(G1324gat));
  OAI21_X1  g251(.A(G8gat), .B1(new_n317_), .B2(new_n259_), .ZN(RLL_wire_A_39));
  XNOR2_X1 RLL_XNOR_39 (.A(RLL_wire_A_39), .B(KEYINPUT39), .ZN(new_n325_) );
  INV_X1    g252(.A(new_n259_), .ZN(new_n326_));
  NAND4_X1  g253(.A1(new_n322_), .A2(new_n176_), .A3(new_n157_), .A4(new_n326_), .ZN(new_n327_));
  NAND2_X1  g254(.A1(new_n327_), .A2(new_n325_), .ZN(RLL_wire_A_40));
  XOR2_X1 RLL_XOR_40 (.A(RLL_wire_A_40), .B(KEYINPUT40), .Z(G1325gat) );
  OAI21_X1  g255(.A(G15gat), .B1(new_n317_), .B2(new_n289_), .ZN(RLL_wire_A_41));
  XOR2_X1 RLL_XOR_41 (.A(RLL_wire_A_41), .B(KEYINPUT41), .Z(new_n329_) );
  NAND4_X1  g256(.A1(new_n322_), .A2(new_n184_), .A3(new_n157_), .A4(new_n287_), .ZN(new_n330_));
  NAND2_X1  g257(.A1(new_n330_), .A2(new_n329_), .ZN(G1326gat));
  OAI21_X1  g258(.A(G22gat), .B1(new_n317_), .B2(new_n274_), .ZN(RLL_wire_A_42));
  XNOR2_X1 RLL_XNOR_42 (.A(RLL_wire_A_42), .B(KEYINPUT42), .ZN(new_n332_) );
  NAND4_X1  g259(.A1(new_n322_), .A2(new_n185_), .A3(new_n157_), .A4(new_n273_), .ZN(new_n333_));
  NAND2_X1  g260(.A1(new_n333_), .A2(new_n332_), .ZN(G1327gat));
  AOI21_X1  g261(.A(new_n321_), .B1(new_n301_), .B2(new_n288_), .ZN(RLL_wire_A_43));
  XOR2_X1 RLL_XOR_43 (.A(RLL_wire_A_43), .B(KEYINPUT43), .Z(new_n335_) );
  NAND4_X1  g262(.A1(new_n335_), .A2(new_n157_), .A3(new_n199_), .A4(new_n213_), .ZN(RLL_wire_A_44));
  XOR2_X1 RLL_XOR_44 (.A(RLL_wire_A_44), .B(KEYINPUT44), .Z(new_n336_) );
  OAI21_X1  g263(.A(G29gat), .B1(new_n336_), .B2(new_n114_), .ZN(new_n337_));
  INV_X1    g264(.A(G29gat), .ZN(new_n338_));
  AND4_X1   g265(.A1(new_n199_), .A2(new_n320_), .A3(new_n213_), .A4(new_n315_), .ZN(new_n339_));
  NAND4_X1  g266(.A1(new_n339_), .A2(new_n338_), .A3(new_n319_), .A4(new_n157_), .ZN(new_n340_));
  NAND2_X1  g267(.A1(new_n340_), .A2(new_n337_), .ZN(G1328gat));
  OAI21_X1  g268(.A(G36gat), .B1(new_n336_), .B2(new_n259_), .ZN(new_n342_));
  INV_X1    g269(.A(G36gat), .ZN(new_n343_));
  NAND4_X1  g270(.A1(new_n339_), .A2(new_n343_), .A3(new_n157_), .A4(new_n326_), .ZN(RLL_wire_A_45));
  XNOR2_X1 RLL_XNOR_45 (.A(RLL_wire_A_45), .B(KEYINPUT45), .ZN(new_n344_) );
  NAND2_X1  g271(.A1(new_n344_), .A2(new_n342_), .ZN(RLL_wire_A_46));
  XOR2_X1 RLL_XOR_46 (.A(RLL_wire_A_46), .B(KEYINPUT46), .Z(G1329gat) );
  OAI21_X1  g272(.A(G43gat), .B1(new_n336_), .B2(new_n289_), .ZN(new_n346_));
  NAND4_X1  g273(.A1(new_n339_), .A2(new_n168_), .A3(new_n157_), .A4(new_n287_), .ZN(new_n347_));
  NAND2_X1  g274(.A1(new_n347_), .A2(new_n346_), .ZN(RLL_wire_A_47));
  XOR2_X1 RLL_XOR_47 (.A(RLL_wire_A_47), .B(KEYINPUT47), .Z(G1330gat) );
  OAI21_X1  g275(.A(G50gat), .B1(new_n336_), .B2(new_n274_), .ZN(new_n349_));
  NAND4_X1  g276(.A1(new_n339_), .A2(new_n169_), .A3(new_n157_), .A4(new_n273_), .ZN(new_n350_));
  NAND2_X1  g277(.A1(new_n350_), .A2(new_n349_), .ZN(G1331gat));
  INV_X1    g278(.A(new_n157_), .ZN(new_n352_));
  NAND4_X1  g279(.A1(new_n316_), .A2(new_n352_), .A3(new_n198_), .A4(new_n214_), .ZN(new_n353_));
  OAI21_X1  g280(.A(G57gat), .B1(new_n353_), .B2(new_n114_), .ZN(new_n354_));
  AND4_X1   g281(.A1(new_n198_), .A2(new_n320_), .A3(new_n214_), .A4(new_n321_), .ZN(new_n355_));
  NAND4_X1  g282(.A1(new_n355_), .A2(new_n134_), .A3(new_n319_), .A4(new_n352_), .ZN(new_n356_));
  NAND2_X1  g283(.A1(new_n356_), .A2(new_n354_), .ZN(G1332gat));
  OAI21_X1  g284(.A(G64gat), .B1(new_n353_), .B2(new_n259_), .ZN(RLL_wire_A_48));
  XNOR2_X1 RLL_XNOR_48 (.A(RLL_wire_A_48), .B(KEYINPUT48), .ZN(new_n358_) );
  NAND4_X1  g285(.A1(new_n355_), .A2(new_n135_), .A3(new_n352_), .A4(new_n326_), .ZN(new_n359_));
  NAND2_X1  g286(.A1(new_n359_), .A2(new_n358_), .ZN(G1333gat));
  OAI21_X1  g287(.A(G71gat), .B1(new_n353_), .B2(new_n289_), .ZN(RLL_wire_A_49));
  XNOR2_X1 RLL_XNOR_49 (.A(RLL_wire_A_49), .B(KEYINPUT49), .ZN(new_n361_) );
  NAND4_X1  g288(.A1(new_n355_), .A2(new_n143_), .A3(new_n352_), .A4(new_n287_), .ZN(new_n362_));
  NAND2_X1  g289(.A1(new_n362_), .A2(new_n361_), .ZN(G1334gat));
  OAI21_X1  g290(.A(G78gat), .B1(new_n353_), .B2(new_n274_), .ZN(RLL_wire_A_50));
  XNOR2_X1 RLL_XNOR_50 (.A(RLL_wire_A_50), .B(KEYINPUT50), .ZN(new_n364_) );
  NAND4_X1  g291(.A1(new_n355_), .A2(new_n144_), .A3(new_n352_), .A4(new_n273_), .ZN(new_n365_));
  NAND2_X1  g292(.A1(new_n365_), .A2(new_n364_), .ZN(G1335gat));
  NAND4_X1  g293(.A1(new_n335_), .A2(new_n352_), .A3(new_n198_), .A4(new_n213_), .ZN(new_n367_));
  OAI21_X1  g294(.A(G85gat), .B1(new_n367_), .B2(new_n114_), .ZN(new_n368_));
  INV_X1    g295(.A(G85gat), .ZN(new_n369_));
  AND4_X1   g296(.A1(new_n198_), .A2(new_n320_), .A3(new_n213_), .A4(new_n315_), .ZN(new_n370_));
  NAND4_X1  g297(.A1(new_n370_), .A2(new_n369_), .A3(new_n319_), .A4(new_n352_), .ZN(new_n371_));
  NAND2_X1  g298(.A1(new_n371_), .A2(new_n368_), .ZN(G1336gat));
  OAI21_X1  g299(.A(G92gat), .B1(new_n367_), .B2(new_n259_), .ZN(new_n373_));
  INV_X1    g300(.A(G92gat), .ZN(new_n374_));
  NAND4_X1  g301(.A1(new_n370_), .A2(new_n374_), .A3(new_n352_), .A4(new_n326_), .ZN(new_n375_));
  NAND2_X1  g302(.A1(new_n375_), .A2(new_n373_), .ZN(G1337gat));
  OAI21_X1  g303(.A(G99gat), .B1(new_n367_), .B2(new_n289_), .ZN(new_n377_));
  NAND4_X1  g304(.A1(new_n370_), .A2(new_n129_), .A3(new_n352_), .A4(new_n287_), .ZN(new_n378_));
  NAND2_X1  g305(.A1(new_n378_), .A2(new_n377_), .ZN(RLL_wire_A_51));
  XNOR2_X1 RLL_XNOR_51 (.A(RLL_wire_A_51), .B(KEYINPUT51), .ZN(G1338gat) );
  OAI21_X1  g306(.A(G106gat), .B1(new_n367_), .B2(new_n274_), .ZN(RLL_wire_A_52));
  XNOR2_X1 RLL_XNOR_52 (.A(RLL_wire_A_52), .B(KEYINPUT52), .ZN(new_n380_) );
  NAND4_X1  g307(.A1(new_n370_), .A2(new_n130_), .A3(new_n352_), .A4(new_n273_), .ZN(new_n381_));
  NAND2_X1  g308(.A1(new_n381_), .A2(new_n380_), .ZN(RLL_wire_A_53));
  XNOR2_X1 RLL_XNOR_53 (.A(RLL_wire_A_53), .B(KEYINPUT53), .ZN(G1339gat) );
  NAND4_X1  g309(.A1(new_n214_), .A2(new_n157_), .A3(new_n198_), .A4(new_n321_), .ZN(RLL_wire_A_54));
  XNOR2_X1 RLL_XNOR_54 (.A(RLL_wire_A_54), .B(KEYINPUT54), .ZN(new_n383_) );
  NAND3_X1  g310(.A1(new_n149_), .A2(new_n118_), .A3(new_n154_), .ZN(new_n384_));
  AOI21_X1  g311(.A(new_n119_), .B1(new_n152_), .B2(new_n153_), .ZN(new_n385_));
  INV_X1    g312(.A(new_n154_), .ZN(RLL_wire_A_55));
  XNOR2_X1 RLL_XNOR_55 (.A(RLL_wire_A_55), .B(KEYINPUT55), .ZN(new_n386_) );
  OAI21_X1  g313(.A(new_n117_), .B1(new_n386_), .B2(new_n385_), .ZN(RLL_wire_A_56));
  XOR2_X1 RLL_XOR_56 (.A(RLL_wire_A_56), .B(KEYINPUT56), .Z(new_n387_) );
  OAI211_X1 g314(.A(new_n384_), .B(new_n387_), .C1(new_n196_), .C2(new_n197_), .ZN(new_n388_));
  NAND3_X1  g315(.A1(new_n190_), .A2(new_n161_), .A3(new_n195_), .ZN(new_n389_));
  AOI21_X1  g316(.A(new_n162_), .B1(new_n193_), .B2(new_n194_), .ZN(new_n390_));
  NOR3_X1   g317(.A1(new_n189_), .A2(new_n188_), .A3(new_n163_), .ZN(new_n391_));
  OAI21_X1  g318(.A(new_n160_), .B1(new_n391_), .B2(new_n390_), .ZN(new_n392_));
  OAI211_X1 g319(.A(new_n389_), .B(new_n392_), .C1(new_n155_), .C2(new_n156_), .ZN(new_n393_));
  AOI21_X1  g320(.A(new_n315_), .B1(new_n388_), .B2(new_n393_), .ZN(RLL_wire_A_57));
  XNOR2_X1 RLL_XNOR_57 (.A(RLL_wire_A_57), .B(KEYINPUT57), .ZN(new_n394_) );
  NAND4_X1  g321(.A1(new_n387_), .A2(new_n392_), .A3(new_n384_), .A4(new_n389_), .ZN(RLL_wire_A_58));
  XOR2_X1 RLL_XOR_58 (.A(RLL_wire_A_58), .B(KEYINPUT58), .Z(new_n395_) );
  NOR2_X1   g322(.A1(new_n321_), .A2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g323(.A(new_n213_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g324(.A(new_n273_), .B1(new_n397_), .B2(new_n383_), .ZN(new_n398_));
  NAND4_X1  g325(.A1(new_n398_), .A2(new_n319_), .A3(new_n259_), .A4(new_n287_), .ZN(RLL_wire_A_59));
  XNOR2_X1 RLL_XNOR_59 (.A(RLL_wire_A_59), .B(KEYINPUT59), .ZN(new_n399_) );
  OAI21_X1  g326(.A(G113gat), .B1(new_n399_), .B2(new_n198_), .ZN(new_n400_));
  INV_X1    g327(.A(G113gat), .ZN(new_n401_));
  NAND2_X1  g328(.A1(new_n397_), .A2(new_n383_), .ZN(new_n402_));
  AND4_X1   g329(.A1(new_n319_), .A2(new_n402_), .A3(new_n274_), .A4(new_n287_), .ZN(new_n403_));
  NAND4_X1  g330(.A1(new_n403_), .A2(new_n401_), .A3(new_n199_), .A4(new_n259_), .ZN(new_n404_));
  NAND2_X1  g331(.A1(new_n404_), .A2(new_n400_), .ZN(G1340gat));
  OAI21_X1  g332(.A(G120gat), .B1(new_n399_), .B2(new_n157_), .ZN(new_n406_));
  INV_X1    g333(.A(G120gat), .ZN(RLL_wire_A_60));
  XOR2_X1 RLL_XOR_60 (.A(RLL_wire_A_60), .B(KEYINPUT60), .Z(new_n407_) );
  NAND4_X1  g334(.A1(new_n403_), .A2(new_n407_), .A3(new_n352_), .A4(new_n259_), .ZN(new_n408_));
  NAND2_X1  g335(.A1(new_n408_), .A2(new_n406_), .ZN(G1341gat));
  OAI21_X1  g336(.A(G127gat), .B1(new_n399_), .B2(new_n213_), .ZN(new_n410_));
  NAND4_X1  g337(.A1(new_n403_), .A2(new_n84_), .A3(new_n214_), .A4(new_n259_), .ZN(new_n411_));
  NAND2_X1  g338(.A1(new_n411_), .A2(new_n410_), .ZN(G1342gat));
  OAI21_X1  g339(.A(G134gat), .B1(new_n399_), .B2(new_n321_), .ZN(new_n413_));
  NAND4_X1  g340(.A1(new_n403_), .A2(new_n85_), .A3(new_n259_), .A4(new_n315_), .ZN(new_n414_));
  NAND2_X1  g341(.A1(new_n414_), .A2(new_n413_), .ZN(G1343gat));
  AOI21_X1  g342(.A(new_n274_), .B1(new_n397_), .B2(new_n383_), .ZN(new_n416_));
  NAND4_X1  g343(.A1(new_n416_), .A2(new_n319_), .A3(new_n259_), .A4(new_n289_), .ZN(new_n417_));
  OAI21_X1  g344(.A(G141gat), .B1(new_n417_), .B2(new_n198_), .ZN(new_n418_));
  AND4_X1   g345(.A1(new_n319_), .A2(new_n402_), .A3(new_n273_), .A4(new_n289_), .ZN(new_n419_));
  NAND4_X1  g346(.A1(new_n419_), .A2(new_n91_), .A3(new_n199_), .A4(new_n259_), .ZN(new_n420_));
  NAND2_X1  g347(.A1(new_n420_), .A2(new_n418_), .ZN(G1344gat));
  OAI21_X1  g348(.A(G148gat), .B1(new_n417_), .B2(new_n157_), .ZN(new_n422_));
  NAND4_X1  g349(.A1(new_n419_), .A2(new_n92_), .A3(new_n352_), .A4(new_n259_), .ZN(new_n423_));
  NAND2_X1  g350(.A1(new_n423_), .A2(new_n422_), .ZN(G1345gat));
  OAI21_X1  g351(.A(G155gat), .B1(new_n417_), .B2(new_n213_), .ZN(new_n425_));
  NAND4_X1  g352(.A1(new_n419_), .A2(new_n100_), .A3(new_n214_), .A4(new_n259_), .ZN(new_n426_));
  NAND2_X1  g353(.A1(new_n426_), .A2(new_n425_), .ZN(RLL_wire_A_61));
  XNOR2_X1 RLL_XNOR_61 (.A(RLL_wire_A_61), .B(KEYINPUT61), .ZN(G1346gat) );
  OAI21_X1  g354(.A(G162gat), .B1(new_n417_), .B2(new_n321_), .ZN(new_n428_));
  NAND4_X1  g355(.A1(new_n419_), .A2(new_n101_), .A3(new_n259_), .A4(new_n315_), .ZN(new_n429_));
  NAND2_X1  g356(.A1(new_n429_), .A2(new_n428_), .ZN(G1347gat));
  NAND4_X1  g357(.A1(new_n398_), .A2(new_n114_), .A3(new_n326_), .A4(new_n287_), .ZN(new_n431_));
  OAI21_X1  g358(.A(G169gat), .B1(new_n431_), .B2(new_n198_), .ZN(RLL_wire_A_62));
  XNOR2_X1 RLL_XNOR_62 (.A(RLL_wire_A_62), .B(KEYINPUT62), .ZN(new_n432_) );
  AND4_X1   g359(.A1(new_n114_), .A2(new_n402_), .A3(new_n274_), .A4(new_n287_), .ZN(new_n433_));
  NAND4_X1  g360(.A1(new_n433_), .A2(new_n236_), .A3(new_n199_), .A4(new_n326_), .ZN(new_n434_));
  NAND2_X1  g361(.A1(new_n434_), .A2(new_n432_), .ZN(G1348gat));
  OAI21_X1  g362(.A(G176gat), .B1(new_n431_), .B2(new_n157_), .ZN(new_n436_));
  NAND4_X1  g363(.A1(new_n433_), .A2(new_n237_), .A3(new_n352_), .A4(new_n326_), .ZN(new_n437_));
  NAND2_X1  g364(.A1(new_n437_), .A2(new_n436_), .ZN(G1349gat));
  OAI21_X1  g365(.A(G183gat), .B1(new_n431_), .B2(new_n213_), .ZN(new_n439_));
  NAND4_X1  g366(.A1(new_n433_), .A2(new_n245_), .A3(new_n214_), .A4(new_n326_), .ZN(new_n440_));
  NAND2_X1  g367(.A1(new_n440_), .A2(new_n439_), .ZN(G1350gat));
  OAI21_X1  g368(.A(G190gat), .B1(new_n431_), .B2(new_n321_), .ZN(new_n442_));
  NAND4_X1  g369(.A1(new_n433_), .A2(new_n246_), .A3(new_n326_), .A4(new_n315_), .ZN(new_n443_));
  NAND2_X1  g370(.A1(new_n443_), .A2(new_n442_), .ZN(G1351gat));
  NAND4_X1  g371(.A1(new_n416_), .A2(new_n114_), .A3(new_n326_), .A4(new_n289_), .ZN(new_n445_));
  OAI21_X1  g372(.A(G197gat), .B1(new_n445_), .B2(new_n198_), .ZN(new_n446_));
  AND4_X1   g373(.A1(new_n114_), .A2(new_n402_), .A3(new_n273_), .A4(new_n289_), .ZN(new_n447_));
  NAND4_X1  g374(.A1(new_n447_), .A2(new_n222_), .A3(new_n199_), .A4(new_n326_), .ZN(new_n448_));
  NAND2_X1  g375(.A1(new_n448_), .A2(new_n446_), .ZN(G1352gat));
  OAI21_X1  g376(.A(G204gat), .B1(new_n445_), .B2(new_n157_), .ZN(new_n450_));
  NAND4_X1  g377(.A1(new_n447_), .A2(new_n223_), .A3(new_n352_), .A4(new_n326_), .ZN(new_n451_));
  NAND2_X1  g378(.A1(new_n451_), .A2(new_n450_), .ZN(G1353gat));
  OAI21_X1  g379(.A(G211gat), .B1(new_n445_), .B2(new_n213_), .ZN(new_n453_));
  NAND4_X1  g380(.A1(new_n447_), .A2(new_n231_), .A3(new_n214_), .A4(new_n326_), .ZN(RLL_wire_A_63));
  XOR2_X1 RLL_XOR_63 (.A(RLL_wire_A_63), .B(KEYINPUT63), .Z(new_n454_) );
  NAND2_X1  g381(.A1(new_n454_), .A2(new_n453_), .ZN(G1354gat));
  OAI21_X1  g382(.A(G218gat), .B1(new_n445_), .B2(new_n321_), .ZN(new_n456_));
  NAND4_X1  g383(.A1(new_n447_), .A2(new_n232_), .A3(new_n326_), .A4(new_n315_), .ZN(new_n457_));
  NAND2_X1  g384(.A1(new_n457_), .A2(new_n456_), .ZN(G1355gat));

endmodule
