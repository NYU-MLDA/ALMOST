//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 0 1 1 0 0 1 0 1 1 0 0 1 0 1 1 0 1 0 1 0 1 0 1 0 0 1 0 1 0 1 1 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n831_, new_n832_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n841_, new_n842_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n874_, new_n875_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_, new_n904_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(G141gat), .ZN(new_n204_));
  INV_X1    g003(.A(G148gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT90), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n206_), .B1(new_n207_), .B2(KEYINPUT3), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT91), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT2), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n209_), .A2(new_n210_), .A3(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n215_), .A2(new_n204_), .A3(new_n205_), .A4(KEYINPUT90), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n208_), .A2(new_n212_), .A3(new_n214_), .A4(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(KEYINPUT89), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n217_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT89), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n218_), .B(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n220_), .B(KEYINPUT1), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n206_), .B(new_n209_), .C1(new_n223_), .C2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n221_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT4), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G127gat), .B(G134gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G113gat), .B(G120gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n226_), .A2(new_n227_), .A3(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n226_), .A2(new_n231_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n221_), .A2(new_n225_), .A3(new_n230_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n203_), .B(new_n232_), .C1(new_n235_), .C2(new_n227_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n233_), .A2(new_n202_), .A3(new_n234_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G1gat), .B(G29gat), .ZN(new_n238_));
  INV_X1    g037(.A(G85gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT0), .B(G57gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n236_), .A2(new_n237_), .A3(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT33), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT33), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n236_), .A2(new_n237_), .A3(new_n245_), .A4(new_n242_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(G169gat), .ZN(new_n248_));
  INV_X1    g047(.A(G176gat), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G183gat), .A2(G190gat), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT23), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n254_), .B(new_n255_), .C1(G183gat), .C2(G190gat), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n248_), .A2(KEYINPUT85), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT22), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n251_), .B(new_n256_), .C1(new_n259_), .C2(G176gat), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT24), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n262_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT84), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n248_), .A2(new_n249_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n251_), .A2(KEYINPUT24), .A3(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT84), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n262_), .A2(new_n254_), .A3(new_n267_), .A4(new_n255_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n264_), .A2(new_n266_), .A3(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT25), .B(G183gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT26), .B(G190gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT83), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n270_), .A2(new_n271_), .A3(KEYINPUT83), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n260_), .B1(new_n269_), .B2(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(G211gat), .B(G218gat), .Z(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(G197gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(G204gat), .ZN(new_n281_));
  INV_X1    g080(.A(G204gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(G197gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT21), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n282_), .A2(G197gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT92), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT92), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n288_), .B1(G197gat), .B2(new_n282_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n287_), .B1(new_n286_), .B2(new_n289_), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n279_), .B(new_n285_), .C1(new_n290_), .C2(KEYINPUT21), .ZN(new_n291_));
  NOR3_X1   g090(.A1(new_n288_), .A2(new_n282_), .A3(G197gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n283_), .A2(KEYINPUT92), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n292_), .B1(new_n281_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT93), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n278_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT21), .B1(new_n290_), .B2(KEYINPUT93), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n291_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n277_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT99), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT99), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n277_), .A2(new_n298_), .A3(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT20), .ZN(new_n304_));
  INV_X1    g103(.A(new_n263_), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n305_), .A2(new_n266_), .A3(new_n272_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT97), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n258_), .A2(new_n248_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n307_), .B(new_n251_), .C1(new_n310_), .C2(G176gat), .ZN(new_n311_));
  AOI21_X1  g110(.A(G176gat), .B1(new_n308_), .B2(new_n309_), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT97), .B1(new_n312_), .B2(new_n250_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n311_), .A2(new_n313_), .A3(new_n256_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT98), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n311_), .A2(new_n313_), .A3(KEYINPUT98), .A4(new_n256_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n306_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n298_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n304_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G226gat), .A2(G233gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n303_), .A2(new_n320_), .A3(new_n323_), .ZN(new_n324_));
  OR2_X1    g123(.A1(new_n276_), .A2(new_n269_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n279_), .B1(new_n290_), .B2(KEYINPUT93), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n294_), .A2(new_n295_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n326_), .A2(KEYINPUT21), .A3(new_n327_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n325_), .A2(new_n328_), .A3(new_n291_), .A4(new_n260_), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n329_), .B(KEYINPUT20), .C1(new_n318_), .C2(new_n319_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n323_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n324_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G8gat), .B(G36gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(G92gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT18), .B(G64gat), .ZN(new_n336_));
  XOR2_X1   g135(.A(new_n335_), .B(new_n336_), .Z(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n333_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n324_), .A2(new_n332_), .A3(new_n337_), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n235_), .A2(KEYINPUT100), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n235_), .A2(KEYINPUT100), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n341_), .A2(new_n203_), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n242_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n202_), .B(new_n232_), .C1(new_n235_), .C2(new_n227_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n247_), .A2(new_n339_), .A3(new_n340_), .A4(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT101), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G228gat), .A2(G233gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT94), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT95), .B(KEYINPUT28), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n351_), .B(new_n352_), .Z(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n221_), .A2(new_n225_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT29), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n298_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  XOR2_X1   g156(.A(G78gat), .B(G106gat), .Z(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n355_), .A2(new_n356_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G22gat), .B(G50gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n359_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n359_), .A2(new_n362_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n354_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  OR2_X1    g165(.A1(new_n359_), .A2(new_n362_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n367_), .A2(new_n353_), .A3(new_n363_), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n324_), .A2(new_n332_), .A3(new_n337_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n337_), .B1(new_n324_), .B2(new_n332_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n372_), .A2(KEYINPUT101), .A3(new_n346_), .A4(new_n247_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n236_), .A2(new_n237_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(new_n344_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(new_n243_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n337_), .A2(KEYINPUT32), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n377_), .B(KEYINPUT102), .Z(new_n378_));
  INV_X1    g177(.A(new_n314_), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n298_), .A2(new_n379_), .A3(new_n306_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n380_), .B1(new_n300_), .B2(new_n302_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n323_), .B1(new_n381_), .B2(KEYINPUT20), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n330_), .A2(new_n331_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  OAI221_X1 g183(.A(new_n376_), .B1(new_n333_), .B2(new_n378_), .C1(new_n384_), .C2(new_n377_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n349_), .A2(new_n369_), .A3(new_n373_), .A4(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n277_), .B(KEYINPUT30), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT87), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT88), .B(KEYINPUT31), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G71gat), .B(G99gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G15gat), .B(G43gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G227gat), .A2(G233gat), .ZN(new_n395_));
  XOR2_X1   g194(.A(new_n395_), .B(KEYINPUT86), .Z(new_n396_));
  XNOR2_X1  g195(.A(new_n394_), .B(new_n396_), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n389_), .A2(new_n391_), .A3(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n391_), .B1(new_n389_), .B2(new_n397_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n387_), .A2(new_n388_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(new_n231_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n402_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n404_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n366_), .A2(new_n368_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n338_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n408_), .A2(KEYINPUT27), .A3(new_n340_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT27), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n410_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n407_), .B1(new_n412_), .B2(new_n376_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n386_), .A2(new_n406_), .A3(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n407_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n376_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n412_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n414_), .A2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G190gat), .B(G218gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G134gat), .B(G162gat), .ZN(new_n421_));
  XOR2_X1   g220(.A(new_n420_), .B(new_n421_), .Z(new_n422_));
  INV_X1    g221(.A(KEYINPUT36), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  OR2_X1    g223(.A1(new_n422_), .A2(new_n423_), .ZN(new_n425_));
  INV_X1    g224(.A(G92gat), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n239_), .A2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(G85gat), .A2(G92gat), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT9), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT65), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT9), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n431_), .B1(new_n239_), .B2(new_n426_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n429_), .A2(new_n430_), .A3(new_n432_), .ZN(new_n433_));
  AND3_X1   g232(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT66), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G99gat), .A2(G106gat), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT6), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT66), .ZN(new_n440_));
  NAND3_X1  g239(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n439_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n436_), .A2(new_n442_), .ZN(new_n443_));
  XOR2_X1   g242(.A(KEYINPUT10), .B(G99gat), .Z(new_n444_));
  INV_X1    g243(.A(G106gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n427_), .A2(KEYINPUT65), .A3(KEYINPUT9), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n433_), .A2(new_n443_), .A3(new_n446_), .A4(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT69), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NOR3_X1   g250(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT67), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n454_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n439_), .A2(KEYINPUT67), .A3(new_n441_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n453_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n427_), .A2(new_n428_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT8), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n443_), .A2(new_n453_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT8), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(new_n462_), .A3(new_n458_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n449_), .B1(new_n460_), .B2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n462_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n458_), .A2(new_n462_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n466_), .B1(new_n443_), .B2(new_n453_), .ZN(new_n467_));
  NOR3_X1   g266(.A1(new_n465_), .A2(new_n467_), .A3(KEYINPUT69), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n448_), .B1(new_n464_), .B2(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(G43gat), .B(G50gat), .Z(new_n470_));
  INV_X1    g269(.A(G29gat), .ZN(new_n471_));
  INV_X1    g270(.A(G36gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G29gat), .A2(G36gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n470_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G43gat), .B(G50gat), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n477_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n476_), .A2(KEYINPUT15), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(KEYINPUT15), .B1(new_n476_), .B2(new_n478_), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n469_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT76), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n448_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n476_), .A2(new_n478_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G232gat), .A2(G233gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT34), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT75), .B(KEYINPUT35), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n485_), .A2(new_n487_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT76), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n469_), .A2(new_n494_), .A3(new_n481_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n483_), .A2(new_n493_), .A3(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n490_), .A2(new_n492_), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n497_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n482_), .A2(new_n499_), .A3(new_n493_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT77), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n482_), .A2(KEYINPUT77), .A3(new_n499_), .A4(new_n493_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n424_), .B(new_n425_), .C1(new_n498_), .C2(new_n504_), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n502_), .A2(new_n503_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n496_), .A2(new_n497_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n506_), .A2(new_n423_), .A3(new_n422_), .A4(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n505_), .A2(new_n508_), .A3(KEYINPUT78), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT79), .B(KEYINPUT37), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n509_), .B(new_n511_), .ZN(new_n512_));
  AND2_X1   g311(.A1(KEYINPUT80), .A2(G8gat), .ZN(new_n513_));
  NOR2_X1   g312(.A1(KEYINPUT80), .A2(G8gat), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT14), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G15gat), .B(G22gat), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n515_), .A2(G1gat), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(G8gat), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT14), .ZN(new_n519_));
  AND2_X1   g318(.A1(G15gat), .A2(G22gat), .ZN(new_n520_));
  NOR2_X1   g319(.A1(G15gat), .A2(G22gat), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n519_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(G1gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n517_), .A2(new_n518_), .A3(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n518_), .B1(new_n517_), .B2(new_n524_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G231gat), .A2(G233gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G57gat), .B(G64gat), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n530_), .A2(KEYINPUT11), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(KEYINPUT11), .ZN(new_n532_));
  XOR2_X1   g331(.A(G71gat), .B(G78gat), .Z(new_n533_));
  NAND3_X1  g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n532_), .A2(new_n533_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT70), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n529_), .B(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G127gat), .B(G155gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(G211gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT16), .B(G183gat), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n540_), .B(new_n541_), .Z(new_n542_));
  INV_X1    g341(.A(KEYINPUT17), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n538_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n536_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n544_), .B1(new_n529_), .B2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n542_), .A2(new_n543_), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n547_), .B(new_n548_), .C1(new_n546_), .C2(new_n529_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n545_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n419_), .A2(new_n512_), .A3(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G113gat), .B(G141gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G169gat), .B(G197gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT81), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n487_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n557_));
  OR2_X1    g356(.A1(KEYINPUT80), .A2(G8gat), .ZN(new_n558_));
  NAND2_X1  g357(.A1(KEYINPUT80), .A2(G8gat), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n519_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(G1gat), .B1(new_n520_), .B2(new_n521_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(G1gat), .B1(new_n516_), .B2(new_n519_), .ZN(new_n563_));
  OAI21_X1  g362(.A(G8gat), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n517_), .A2(new_n518_), .A3(new_n524_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n564_), .A2(new_n486_), .A3(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n557_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G229gat), .A2(G233gat), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n564_), .B(new_n565_), .C1(new_n479_), .C2(new_n480_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n571_), .A2(new_n557_), .A3(new_n568_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n556_), .B1(new_n570_), .B2(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n568_), .B1(new_n557_), .B2(new_n566_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n574_), .A2(KEYINPUT81), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n555_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT82), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n571_), .A2(new_n557_), .A3(new_n568_), .ZN(new_n578_));
  OAI21_X1  g377(.A(KEYINPUT81), .B1(new_n578_), .B2(new_n574_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n570_), .A2(new_n556_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n555_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n576_), .A2(new_n577_), .A3(new_n582_), .ZN(new_n583_));
  OAI211_X1 g382(.A(KEYINPUT82), .B(new_n555_), .C1(new_n573_), .C2(new_n575_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n552_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT73), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n484_), .A2(new_n546_), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n536_), .B(new_n448_), .C1(new_n465_), .C2(new_n467_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G230gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT64), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n591_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(KEYINPUT68), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n593_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT68), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n469_), .A2(KEYINPUT12), .A3(new_n537_), .ZN(new_n601_));
  OR2_X1    g400(.A1(KEYINPUT71), .A2(KEYINPUT12), .ZN(new_n602_));
  NAND2_X1  g401(.A1(KEYINPUT71), .A2(KEYINPUT12), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n589_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n601_), .A2(new_n593_), .A3(new_n590_), .A4(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G176gat), .B(G204gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G120gat), .B(G148gat), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n608_), .B(new_n609_), .Z(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n600_), .A2(new_n605_), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n611_), .B1(new_n600_), .B2(new_n605_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n588_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  AND4_X1   g414(.A1(new_n593_), .A2(new_n601_), .A3(new_n590_), .A4(new_n604_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n597_), .B(KEYINPUT68), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n610_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n618_), .A2(KEYINPUT73), .A3(new_n612_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n615_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT13), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(KEYINPUT13), .B1(new_n615_), .B2(new_n619_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT74), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n587_), .A2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n627_), .A2(new_n523_), .A3(new_n376_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT38), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n622_), .A2(new_n623_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n630_), .A2(new_n585_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n505_), .A2(new_n508_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n633_), .B1(new_n414_), .B2(new_n418_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n631_), .A2(new_n551_), .A3(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(G1gat), .B1(new_n635_), .B2(new_n416_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n629_), .A2(new_n636_), .ZN(G1324gat));
  NAND2_X1  g436(.A1(new_n558_), .A2(new_n559_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n587_), .A2(new_n638_), .A3(new_n412_), .A4(new_n626_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT103), .Z(new_n640_));
  OAI21_X1  g439(.A(G8gat), .B1(new_n635_), .B2(new_n417_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT104), .ZN(new_n642_));
  OAI21_X1  g441(.A(KEYINPUT39), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n642_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n640_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT40), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n646_), .B(new_n647_), .ZN(G1325gat));
  OAI21_X1  g447(.A(G15gat), .B1(new_n635_), .B2(new_n406_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT41), .Z(new_n650_));
  INV_X1    g449(.A(G15gat), .ZN(new_n651_));
  INV_X1    g450(.A(new_n406_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n627_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n650_), .A2(new_n653_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT105), .Z(G1326gat));
  XNOR2_X1  g454(.A(new_n407_), .B(KEYINPUT106), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G22gat), .B1(new_n635_), .B2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT42), .ZN(new_n659_));
  INV_X1    g458(.A(G22gat), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n627_), .A2(new_n660_), .A3(new_n656_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n661_), .ZN(G1327gat));
  XNOR2_X1  g461(.A(new_n509_), .B(new_n510_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n419_), .A2(new_n663_), .A3(KEYINPUT43), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT43), .B1(new_n419_), .B2(new_n663_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n666_), .A2(KEYINPUT44), .A3(new_n550_), .A4(new_n631_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n419_), .A2(new_n663_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT43), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n419_), .A2(new_n663_), .A3(KEYINPUT43), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n670_), .A2(new_n550_), .A3(new_n631_), .A4(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n667_), .A2(new_n674_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n675_), .A2(new_n471_), .A3(new_n416_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n632_), .B1(new_n414_), .B2(new_n418_), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n631_), .A2(new_n550_), .A3(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(G29gat), .B1(new_n678_), .B2(new_n376_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n676_), .A2(new_n679_), .ZN(G1328gat));
  NOR2_X1   g479(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT109), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT46), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n667_), .A2(new_n674_), .A3(new_n412_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n667_), .A2(new_n674_), .A3(KEYINPUT107), .A4(new_n412_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(G36gat), .A3(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n412_), .B(KEYINPUT108), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n678_), .A2(new_n472_), .A3(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT45), .ZN(new_n692_));
  AOI211_X1 g491(.A(new_n681_), .B(new_n684_), .C1(new_n689_), .C2(new_n692_), .ZN(new_n693_));
  AND4_X1   g492(.A1(new_n682_), .A2(new_n689_), .A3(new_n683_), .A4(new_n692_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1329gat));
  NAND2_X1  g494(.A1(new_n652_), .A2(G43gat), .ZN(new_n696_));
  INV_X1    g495(.A(new_n678_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n697_), .A2(new_n406_), .ZN(new_n698_));
  OAI22_X1  g497(.A1(new_n675_), .A2(new_n696_), .B1(G43gat), .B2(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n699_), .B(new_n700_), .ZN(G1330gat));
  OAI21_X1  g500(.A(G50gat), .B1(new_n675_), .B2(new_n369_), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n657_), .A2(G50gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n697_), .B2(new_n703_), .ZN(G1331gat));
  NOR2_X1   g503(.A1(new_n624_), .A2(new_n586_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n552_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT111), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT111), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n416_), .B1(new_n706_), .B2(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(G57gat), .B1(new_n708_), .B2(new_n710_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n586_), .A2(new_n550_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n625_), .A2(new_n634_), .A3(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT112), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n625_), .A2(KEYINPUT112), .A3(new_n634_), .A4(new_n712_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n376_), .A2(G57gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n711_), .B1(new_n717_), .B2(new_n718_), .ZN(G1332gat));
  INV_X1    g518(.A(G64gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n720_), .B1(new_n717_), .B2(new_n690_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT48), .Z(new_n722_));
  NAND3_X1  g521(.A1(new_n707_), .A2(new_n720_), .A3(new_n690_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1333gat));
  OR3_X1    g523(.A1(new_n706_), .A2(G71gat), .A3(new_n406_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n715_), .A2(new_n652_), .A3(new_n716_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(KEYINPUT113), .B(KEYINPUT49), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n726_), .A2(G71gat), .A3(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n726_), .B2(G71gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT114), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n730_), .B(new_n731_), .ZN(G1334gat));
  INV_X1    g531(.A(G78gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n717_), .B2(new_n656_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT50), .Z(new_n735_));
  NAND3_X1  g534(.A1(new_n707_), .A2(new_n733_), .A3(new_n656_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1335gat));
  AND4_X1   g536(.A1(new_n550_), .A2(new_n625_), .A3(new_n585_), .A4(new_n677_), .ZN(new_n738_));
  AOI21_X1  g537(.A(G85gat), .B1(new_n738_), .B2(new_n376_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n670_), .A2(new_n550_), .A3(new_n671_), .A4(new_n705_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n740_), .A2(new_n239_), .A3(new_n416_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n739_), .A2(new_n741_), .ZN(G1336gat));
  AOI21_X1  g541(.A(G92gat), .B1(new_n738_), .B2(new_n412_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n690_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n740_), .A2(new_n426_), .A3(new_n744_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1337gat));
  NAND3_X1  g545(.A1(new_n738_), .A2(new_n444_), .A3(new_n652_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G99gat), .B1(new_n740_), .B2(new_n406_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g549(.A(G106gat), .B1(new_n740_), .B2(new_n369_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT52), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n738_), .A2(new_n445_), .A3(new_n407_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n754_), .B(new_n755_), .ZN(G1339gat));
  NAND3_X1  g555(.A1(new_n512_), .A2(new_n624_), .A3(new_n712_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT54), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n512_), .A2(new_n624_), .A3(KEYINPUT54), .A4(new_n712_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n612_), .A2(new_n584_), .A3(new_n583_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT116), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n612_), .A2(new_n583_), .A3(KEYINPUT116), .A4(new_n584_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n605_), .A2(KEYINPUT117), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT55), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n601_), .A2(new_n590_), .A3(new_n604_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n594_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT55), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n605_), .A2(KEYINPUT117), .A3(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n768_), .A2(new_n770_), .A3(new_n772_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n773_), .A2(KEYINPUT56), .A3(new_n610_), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT56), .B1(new_n773_), .B2(new_n610_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n766_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT118), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n567_), .A2(new_n568_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n571_), .A2(new_n557_), .A3(new_n569_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(new_n555_), .A3(new_n779_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n582_), .A2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n620_), .A2(new_n777_), .A3(new_n781_), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n613_), .A2(new_n614_), .A3(new_n588_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT73), .B1(new_n618_), .B2(new_n612_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n781_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT118), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n776_), .A2(new_n782_), .A3(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(KEYINPUT57), .A3(new_n632_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT119), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n632_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT57), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n612_), .B(new_n781_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT58), .ZN(new_n794_));
  OR2_X1    g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n794_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n663_), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT119), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n787_), .A2(new_n798_), .A3(KEYINPUT57), .A4(new_n632_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n789_), .A2(new_n792_), .A3(new_n797_), .A4(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n761_), .B1(new_n800_), .B2(new_n550_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n415_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n802_), .A2(new_n412_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n801_), .A2(new_n416_), .A3(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(G113gat), .B1(new_n805_), .B2(new_n586_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n800_), .A2(new_n550_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n761_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n809_), .A2(KEYINPUT120), .A3(new_n376_), .A4(new_n803_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT59), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n805_), .A2(KEYINPUT120), .A3(KEYINPUT59), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n585_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n806_), .B1(new_n814_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g614(.A(KEYINPUT60), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(new_n624_), .B2(G120gat), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n805_), .B(new_n817_), .C1(new_n816_), .C2(G120gat), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n626_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n819_));
  INV_X1    g618(.A(G120gat), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n818_), .B1(new_n819_), .B2(new_n820_), .ZN(G1341gat));
  INV_X1    g620(.A(KEYINPUT121), .ZN(new_n822_));
  NOR4_X1   g621(.A1(new_n801_), .A2(new_n416_), .A3(new_n550_), .A4(new_n804_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n823_), .B2(G127gat), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n809_), .A2(new_n376_), .A3(new_n551_), .A4(new_n803_), .ZN(new_n825_));
  INV_X1    g624(.A(G127gat), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(KEYINPUT121), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n824_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n550_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(G127gat), .B2(new_n829_), .ZN(G1342gat));
  AOI21_X1  g629(.A(G134gat), .B1(new_n805_), .B2(new_n633_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n512_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(G134gat), .ZN(G1343gat));
  NOR3_X1   g632(.A1(new_n801_), .A2(new_n416_), .A3(new_n690_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n652_), .A2(new_n369_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n586_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(G141gat), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n836_), .A2(new_n204_), .A3(new_n586_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(G1344gat));
  NAND3_X1  g639(.A1(new_n834_), .A2(new_n625_), .A3(new_n835_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(KEYINPUT122), .B(G148gat), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n841_), .B(new_n842_), .ZN(G1345gat));
  NAND3_X1  g642(.A1(new_n834_), .A2(new_n551_), .A3(new_n835_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(KEYINPUT61), .B(G155gat), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(G1346gat));
  NAND2_X1  g645(.A1(new_n836_), .A2(new_n633_), .ZN(new_n847_));
  INV_X1    g646(.A(G162gat), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n512_), .A2(new_n848_), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n847_), .A2(new_n848_), .B1(new_n836_), .B2(new_n849_), .ZN(G1347gat));
  NOR2_X1   g649(.A1(new_n744_), .A2(new_n376_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n852_), .A2(new_n406_), .A3(new_n656_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n809_), .A2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n586_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT62), .ZN(new_n857_));
  OR2_X1    g656(.A1(new_n857_), .A2(KEYINPUT123), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(KEYINPUT123), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n856_), .A2(G169gat), .A3(new_n858_), .A4(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n854_), .A2(new_n585_), .ZN(new_n861_));
  OAI211_X1 g660(.A(KEYINPUT123), .B(new_n857_), .C1(new_n861_), .C2(new_n248_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n860_), .B(new_n862_), .C1(new_n310_), .C2(new_n856_), .ZN(G1348gat));
  OAI21_X1  g662(.A(new_n249_), .B1(new_n854_), .B2(new_n624_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT124), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n865_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n801_), .A2(new_n802_), .A3(new_n852_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n626_), .A2(new_n249_), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n866_), .A2(new_n867_), .B1(new_n868_), .B2(new_n869_), .ZN(G1349gat));
  NOR3_X1   g669(.A1(new_n854_), .A2(new_n550_), .A3(new_n270_), .ZN(new_n871_));
  AOI21_X1  g670(.A(G183gat), .B1(new_n868_), .B2(new_n551_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1350gat));
  OAI21_X1  g672(.A(G190gat), .B1(new_n854_), .B2(new_n512_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n633_), .A2(new_n271_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n854_), .B2(new_n875_), .ZN(G1351gat));
  NAND3_X1  g675(.A1(new_n809_), .A2(new_n835_), .A3(new_n851_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT125), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n852_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n880_), .A2(KEYINPUT125), .A3(new_n835_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n882_), .A2(new_n280_), .A3(new_n586_), .ZN(new_n883_));
  AOI21_X1  g682(.A(KEYINPUT125), .B1(new_n880_), .B2(new_n835_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n835_), .ZN(new_n885_));
  NOR4_X1   g684(.A1(new_n801_), .A2(new_n878_), .A3(new_n885_), .A4(new_n852_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n586_), .B1(new_n884_), .B2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(G197gat), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n883_), .A2(new_n888_), .ZN(G1352gat));
  OAI21_X1  g688(.A(new_n625_), .B1(new_n884_), .B2(new_n886_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT126), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n890_), .A2(new_n891_), .A3(G204gat), .ZN(new_n892_));
  OAI221_X1 g691(.A(new_n625_), .B1(KEYINPUT126), .B2(new_n282_), .C1(new_n884_), .C2(new_n886_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(G1353gat));
  OR2_X1    g693(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n895_), .B1(new_n882_), .B2(new_n551_), .ZN(new_n896_));
  XOR2_X1   g695(.A(KEYINPUT63), .B(G211gat), .Z(new_n897_));
  OAI211_X1 g696(.A(new_n551_), .B(new_n897_), .C1(new_n884_), .C2(new_n886_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n896_), .A2(new_n899_), .ZN(G1354gat));
  INV_X1    g699(.A(G218gat), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n633_), .B1(new_n884_), .B2(new_n886_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n663_), .A2(G218gat), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(KEYINPUT127), .ZN(new_n904_));
  AOI22_X1  g703(.A1(new_n901_), .A2(new_n902_), .B1(new_n882_), .B2(new_n904_), .ZN(G1355gat));
endmodule


