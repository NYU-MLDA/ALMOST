//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 0 0 0 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n863_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT64), .Z(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  AND2_X1   g003(.A1(G57gat), .A2(G64gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G57gat), .A2(G64gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT67), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G57gat), .ZN(new_n208_));
  INV_X1    g007(.A(G64gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT67), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G57gat), .A2(G64gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT11), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n207_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G71gat), .A2(G78gat), .ZN(new_n216_));
  INV_X1    g015(.A(G71gat), .ZN(new_n217_));
  INV_X1    g016(.A(G78gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  AND3_X1   g018(.A1(new_n215_), .A2(new_n216_), .A3(new_n219_), .ZN(new_n220_));
  NOR3_X1   g019(.A1(new_n205_), .A2(new_n206_), .A3(KEYINPUT67), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n211_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT11), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT68), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n207_), .A2(new_n213_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT68), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(KEYINPUT11), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n220_), .A2(new_n224_), .A3(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n215_), .A2(new_n216_), .A3(new_n219_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n226_), .B1(new_n225_), .B2(KEYINPUT11), .ZN(new_n230_));
  AOI211_X1 g029(.A(KEYINPUT68), .B(new_n214_), .C1(new_n207_), .C2(new_n213_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n229_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n228_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n234_));
  AND2_X1   g033(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n235_));
  NOR2_X1   g034(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n236_));
  INV_X1    g035(.A(G85gat), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n234_), .B1(new_n238_), .B2(KEYINPUT9), .ZN(new_n239_));
  NOR2_X1   g038(.A1(G85gat), .A2(G92gat), .ZN(new_n240_));
  AND2_X1   g039(.A1(G85gat), .A2(G92gat), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n240_), .B1(new_n241_), .B2(KEYINPUT9), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT9), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT65), .B(G92gat), .ZN(new_n244_));
  OAI211_X1 g043(.A(KEYINPUT66), .B(new_n243_), .C1(new_n244_), .C2(new_n237_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n239_), .A2(new_n242_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G99gat), .A2(G106gat), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT6), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(KEYINPUT10), .B(G99gat), .Z(new_n252_));
  INV_X1    g051(.A(G106gat), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n251_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n246_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT7), .ZN(new_n256_));
  INV_X1    g055(.A(G99gat), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(new_n257_), .A3(new_n253_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n258_), .A2(new_n249_), .A3(new_n250_), .A4(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n241_), .A2(new_n240_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT8), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT8), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n260_), .A2(new_n264_), .A3(new_n261_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n255_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n233_), .A2(new_n267_), .ZN(new_n268_));
  AOI22_X1  g067(.A1(new_n246_), .A2(new_n254_), .B1(new_n263_), .B2(new_n265_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n269_), .A2(new_n228_), .A3(new_n232_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n268_), .A2(KEYINPUT12), .A3(new_n270_), .ZN(new_n271_));
  AOI22_X1  g070(.A1(new_n228_), .A2(new_n232_), .B1(new_n255_), .B2(new_n266_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT12), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n204_), .B1(new_n271_), .B2(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n203_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT69), .B(G204gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT5), .B(G176gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G120gat), .B(G148gat), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n279_), .B(new_n280_), .Z(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  OR3_X1    g081(.A1(new_n275_), .A2(new_n276_), .A3(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n282_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n284_));
  AND3_X1   g083(.A1(new_n283_), .A2(KEYINPUT13), .A3(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(KEYINPUT13), .B1(new_n283_), .B2(new_n284_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G15gat), .B(G22gat), .ZN(new_n288_));
  INV_X1    g087(.A(G1gat), .ZN(new_n289_));
  INV_X1    g088(.A(G8gat), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT14), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n288_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G1gat), .B(G8gat), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n293_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G29gat), .B(G36gat), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G43gat), .B(G50gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(G43gat), .B(G50gat), .Z(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n297_), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n296_), .B(new_n303_), .Z(new_n304_));
  NAND2_X1  g103(.A1(new_n300_), .A2(new_n302_), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n300_), .A2(new_n302_), .A3(KEYINPUT15), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT15), .B1(new_n300_), .B2(new_n302_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  MUX2_X1   g107(.A(new_n305_), .B(new_n308_), .S(new_n296_), .Z(new_n309_));
  NAND2_X1  g108(.A1(G229gat), .A2(G233gat), .ZN(new_n310_));
  MUX2_X1   g109(.A(new_n304_), .B(new_n309_), .S(new_n310_), .Z(new_n311_));
  XNOR2_X1  g110(.A(G113gat), .B(G141gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G169gat), .B(G197gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n311_), .B(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n287_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(G169gat), .ZN(new_n317_));
  INV_X1    g116(.A(G176gat), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NOR3_X1   g120(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT75), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G183gat), .A2(G190gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT23), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT75), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT25), .B(G183gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT74), .ZN(new_n329_));
  INV_X1    g128(.A(G190gat), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n329_), .B1(new_n330_), .B2(KEYINPUT26), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT26), .B(G190gat), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n328_), .B(new_n331_), .C1(new_n332_), .C2(new_n329_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n323_), .A2(new_n325_), .A3(new_n327_), .A4(new_n333_), .ZN(new_n334_));
  OR2_X1    g133(.A1(G183gat), .A2(G190gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n325_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n319_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n317_), .A2(KEYINPUT22), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT76), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n317_), .A2(KEYINPUT22), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n317_), .A2(KEYINPUT76), .A3(KEYINPUT22), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n340_), .A2(new_n341_), .A3(new_n318_), .A4(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n336_), .A2(new_n337_), .A3(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n334_), .A2(new_n344_), .ZN(new_n345_));
  OR2_X1    g144(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n347_));
  AOI21_X1  g146(.A(G197gat), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(G197gat), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT88), .B1(new_n349_), .B2(G204gat), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT88), .ZN(new_n351_));
  INV_X1    g150(.A(G204gat), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(new_n352_), .A3(G197gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n350_), .A2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT21), .B1(new_n348_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT21), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n349_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(G197gat), .A2(G204gat), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n356_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G211gat), .B(G218gat), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n355_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n357_), .A2(new_n358_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n360_), .A2(new_n356_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  AND3_X1   g163(.A1(new_n361_), .A2(KEYINPUT90), .A3(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(KEYINPUT90), .B1(new_n361_), .B2(new_n364_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n345_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G226gat), .A2(G233gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT19), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n361_), .A2(new_n364_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n341_), .A2(new_n318_), .A3(new_n338_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT94), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n325_), .A2(new_n373_), .A3(new_n335_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n373_), .B1(new_n325_), .B2(new_n335_), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n372_), .B(new_n337_), .C1(new_n374_), .C2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n321_), .A2(new_n322_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n332_), .A2(new_n328_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(new_n325_), .A3(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n371_), .A2(new_n376_), .A3(new_n379_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n367_), .A2(KEYINPUT20), .A3(new_n370_), .A4(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT95), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G8gat), .B(G36gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(G92gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT18), .B(G64gat), .ZN(new_n385_));
  XOR2_X1   g184(.A(new_n384_), .B(new_n385_), .Z(new_n386_));
  NAND2_X1  g185(.A1(new_n376_), .A2(new_n379_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n361_), .A2(new_n364_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT90), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n361_), .A2(KEYINPUT90), .A3(new_n364_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  OAI211_X1 g192(.A(KEYINPUT20), .B(new_n389_), .C1(new_n393_), .C2(new_n345_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n369_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n382_), .A2(KEYINPUT100), .A3(new_n386_), .A4(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT20), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n397_), .B1(new_n393_), .B2(new_n345_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n398_), .A2(KEYINPUT95), .A3(new_n370_), .A4(new_n380_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT95), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n381_), .A2(new_n400_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n399_), .A2(new_n401_), .A3(new_n395_), .A4(new_n386_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT100), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n398_), .A2(new_n369_), .A3(new_n380_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n394_), .A2(new_n370_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n386_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n396_), .A2(KEYINPUT27), .A3(new_n404_), .A4(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n399_), .A2(new_n401_), .A3(new_n395_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(new_n408_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n402_), .ZN(new_n413_));
  XOR2_X1   g212(.A(KEYINPUT101), .B(KEYINPUT27), .Z(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n410_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(G228gat), .ZN(new_n417_));
  INV_X1    g216(.A(G233gat), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT29), .ZN(new_n420_));
  AOI21_X1  g219(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT83), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n423_));
  NOR2_X1   g222(.A1(G141gat), .A2(G148gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT82), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT84), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n430_));
  NAND4_X1  g229(.A1(KEYINPUT84), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n429_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT82), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT3), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n434_), .A2(KEYINPUT81), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(KEYINPUT81), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n433_), .B(new_n424_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n422_), .A2(new_n426_), .A3(new_n432_), .A4(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(G155gat), .A2(G162gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT80), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G155gat), .A2(G162gat), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n438_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n424_), .B(KEYINPUT79), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G141gat), .A2(G148gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n442_), .B(KEYINPUT1), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n444_), .B(new_n445_), .C1(new_n440_), .C2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n420_), .B1(new_n443_), .B2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n419_), .B1(new_n448_), .B2(new_n371_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT91), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  OAI211_X1 g250(.A(KEYINPUT91), .B(new_n419_), .C1(new_n448_), .C2(new_n371_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n448_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n419_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n453_), .A2(new_n456_), .ZN(new_n457_));
  XOR2_X1   g256(.A(G78gat), .B(G106gat), .Z(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n457_), .A2(KEYINPUT93), .A3(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n443_), .A2(new_n420_), .A3(new_n447_), .ZN(new_n461_));
  XOR2_X1   g260(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n462_));
  XOR2_X1   g261(.A(new_n461_), .B(new_n462_), .Z(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT87), .B(G50gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT85), .B(G22gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n463_), .B(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT93), .ZN(new_n468_));
  AOI22_X1  g267(.A1(new_n451_), .A2(new_n452_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n469_));
  XOR2_X1   g268(.A(new_n458_), .B(KEYINPUT92), .Z(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n468_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n469_), .A2(new_n458_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n460_), .B(new_n467_), .C1(new_n472_), .C2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT78), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT30), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n334_), .A2(new_n476_), .A3(new_n344_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n476_), .B1(new_n334_), .B2(new_n344_), .ZN(new_n478_));
  OAI21_X1  g277(.A(G43gat), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n345_), .A2(KEYINPUT30), .ZN(new_n480_));
  INV_X1    g279(.A(G43gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n334_), .A2(new_n476_), .A3(new_n344_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n480_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G227gat), .A2(G233gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(G15gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G71gat), .B(G99gat), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n485_), .B(new_n486_), .Z(new_n487_));
  AND3_X1   g286(.A1(new_n479_), .A2(new_n483_), .A3(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n487_), .B1(new_n479_), .B2(new_n483_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n475_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n479_), .A2(new_n483_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n487_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n479_), .A2(new_n483_), .A3(new_n487_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(KEYINPUT78), .A3(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT77), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G127gat), .B(G134gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G113gat), .B(G120gat), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n496_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  XOR2_X1   g298(.A(G127gat), .B(G134gat), .Z(new_n500_));
  XOR2_X1   g299(.A(G113gat), .B(G120gat), .Z(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n499_), .B(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT31), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n490_), .A2(new_n495_), .A3(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n504_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n475_), .B(new_n506_), .C1(new_n488_), .C2(new_n489_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n466_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n463_), .B(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n457_), .A2(new_n470_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n469_), .A2(new_n471_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n510_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n474_), .A2(new_n508_), .A3(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT102), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n500_), .B(new_n498_), .ZN(new_n516_));
  AND3_X1   g315(.A1(new_n443_), .A2(new_n447_), .A3(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n503_), .B1(new_n443_), .B2(new_n447_), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT4), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n443_), .A2(new_n447_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT4), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n521_), .A3(new_n503_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT97), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G225gat), .A2(G233gat), .ZN(new_n524_));
  XOR2_X1   g323(.A(new_n524_), .B(KEYINPUT96), .Z(new_n525_));
  INV_X1    g324(.A(KEYINPUT97), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n520_), .A2(new_n526_), .A3(new_n521_), .A4(new_n503_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n519_), .A2(new_n523_), .A3(new_n525_), .A4(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n524_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT98), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  OAI211_X1 g330(.A(KEYINPUT98), .B(new_n524_), .C1(new_n517_), .C2(new_n518_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n528_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G1gat), .B(G29gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(new_n237_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT0), .B(G57gat), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n535_), .B(new_n536_), .Z(new_n537_));
  NAND2_X1  g336(.A1(new_n533_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n537_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n528_), .A2(new_n531_), .A3(new_n532_), .A4(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n416_), .A2(new_n514_), .A3(new_n515_), .A4(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n410_), .A2(new_n415_), .A3(new_n542_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n474_), .A2(new_n513_), .A3(new_n508_), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT102), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n540_), .B(KEYINPUT33), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n519_), .A2(new_n523_), .A3(new_n524_), .A4(new_n527_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n525_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(new_n537_), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT99), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n548_), .A2(new_n553_), .A3(new_n402_), .A4(new_n412_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n474_), .A2(new_n513_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n386_), .A2(KEYINPUT32), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  AOI22_X1  g356(.A1(new_n538_), .A2(new_n540_), .B1(new_n407_), .B2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n382_), .A2(new_n395_), .A3(new_n556_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n554_), .A2(new_n555_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n474_), .A2(new_n513_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n544_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n508_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n561_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n316_), .B1(new_n547_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G231gat), .A2(G233gat), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n296_), .B(new_n567_), .Z(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(new_n233_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(G127gat), .B(G155gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT73), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G183gat), .B(G211gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n576_), .A2(KEYINPUT17), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(KEYINPUT17), .ZN(new_n578_));
  OR3_X1    g377(.A1(new_n570_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n570_), .A2(new_n577_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n255_), .A2(new_n303_), .A3(new_n266_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT70), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G232gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT34), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n584_), .A2(KEYINPUT35), .A3(new_n586_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n586_), .A2(KEYINPUT35), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n588_), .B1(new_n269_), .B2(new_n308_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n255_), .A2(new_n303_), .A3(new_n266_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n587_), .A2(new_n591_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n583_), .B(new_n588_), .C1(new_n308_), .C2(new_n269_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n593_), .A2(KEYINPUT35), .A3(new_n586_), .A4(new_n584_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n592_), .A2(new_n594_), .A3(KEYINPUT71), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G190gat), .B(G218gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G134gat), .B(G162gat), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n596_), .B(new_n597_), .Z(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n599_), .A2(KEYINPUT36), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n595_), .A2(new_n601_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n592_), .A2(new_n594_), .A3(KEYINPUT71), .A4(new_n600_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n592_), .A2(new_n594_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n605_), .A2(KEYINPUT36), .A3(new_n599_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n582_), .A2(new_n607_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n566_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(G1gat), .B1(new_n610_), .B2(new_n542_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n607_), .A2(KEYINPUT37), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT37), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n604_), .A2(new_n613_), .A3(new_n606_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n615_), .A2(new_n582_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n566_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n617_), .A2(new_n289_), .A3(new_n541_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT103), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n619_), .A2(KEYINPUT38), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(KEYINPUT38), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n611_), .B1(new_n620_), .B2(new_n621_), .ZN(G1324gat));
  INV_X1    g421(.A(KEYINPUT40), .ZN(new_n623_));
  INV_X1    g422(.A(new_n416_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n609_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(G8gat), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n617_), .A2(new_n290_), .A3(new_n624_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT104), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n623_), .B1(new_n628_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n630_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n626_), .B(KEYINPUT39), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n632_), .A2(new_n633_), .A3(KEYINPUT40), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n631_), .A2(new_n634_), .ZN(G1325gat));
  INV_X1    g434(.A(G15gat), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n636_), .B1(new_n609_), .B2(new_n508_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT41), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n617_), .A2(new_n636_), .A3(new_n508_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(G1326gat));
  INV_X1    g439(.A(G22gat), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n617_), .A2(new_n641_), .A3(new_n562_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n641_), .B1(new_n609_), .B2(new_n562_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT105), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT42), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n643_), .A2(new_n644_), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n645_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n646_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n642_), .B1(new_n648_), .B2(new_n649_), .ZN(G1327gat));
  INV_X1    g449(.A(KEYINPUT106), .ZN(new_n651_));
  INV_X1    g450(.A(new_n607_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n581_), .A2(new_n652_), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n566_), .A2(new_n651_), .A3(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n651_), .B1(new_n566_), .B2(new_n653_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(G29gat), .B1(new_n656_), .B2(new_n541_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n316_), .A2(new_n581_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT43), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n547_), .A2(new_n565_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n660_), .B2(new_n615_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n615_), .ZN(new_n662_));
  AOI211_X1 g461(.A(KEYINPUT43), .B(new_n662_), .C1(new_n547_), .C2(new_n565_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n658_), .B1(new_n661_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n666_), .A2(G29gat), .A3(new_n541_), .ZN(new_n667_));
  OAI211_X1 g466(.A(KEYINPUT44), .B(new_n658_), .C1(new_n661_), .C2(new_n663_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n657_), .B1(new_n667_), .B2(new_n668_), .ZN(G1328gat));
  INV_X1    g468(.A(G36gat), .ZN(new_n670_));
  INV_X1    g469(.A(new_n658_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n551_), .B(KEYINPUT99), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n672_), .A2(new_n413_), .ZN(new_n673_));
  AOI22_X1  g472(.A1(new_n673_), .A2(new_n548_), .B1(new_n559_), .B2(new_n558_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n508_), .B1(new_n674_), .B2(new_n555_), .ZN(new_n675_));
  AOI22_X1  g474(.A1(new_n675_), .A2(new_n563_), .B1(new_n546_), .B2(new_n543_), .ZN(new_n676_));
  OAI21_X1  g475(.A(KEYINPUT43), .B1(new_n676_), .B2(new_n662_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n660_), .A2(new_n659_), .A3(new_n615_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n671_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n416_), .B1(new_n679_), .B2(KEYINPUT44), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n670_), .B1(new_n680_), .B2(new_n666_), .ZN(new_n681_));
  XOR2_X1   g480(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n682_));
  NAND4_X1  g481(.A1(new_n656_), .A2(new_n670_), .A3(new_n624_), .A4(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n316_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n660_), .A2(new_n684_), .A3(new_n653_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT106), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n566_), .A2(new_n651_), .A3(new_n653_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n686_), .A2(new_n670_), .A3(new_n624_), .A4(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n682_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n683_), .A2(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n681_), .A2(new_n691_), .A3(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n688_), .B(new_n682_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n668_), .A2(new_n624_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n677_), .A2(new_n678_), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT44), .B1(new_n697_), .B2(new_n658_), .ZN(new_n698_));
  OAI21_X1  g497(.A(G36gat), .B1(new_n696_), .B2(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n692_), .B1(new_n695_), .B2(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n694_), .A2(new_n700_), .ZN(G1329gat));
  NAND4_X1  g500(.A1(new_n666_), .A2(G43gat), .A3(new_n508_), .A4(new_n668_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(KEYINPUT109), .B(G43gat), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n686_), .A2(new_n687_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n704_), .B2(new_n564_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n702_), .A2(new_n705_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g506(.A(G50gat), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n668_), .A2(new_n562_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n708_), .B1(new_n710_), .B2(new_n666_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n562_), .A2(new_n708_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT110), .Z(new_n713_));
  NOR2_X1   g512(.A1(new_n704_), .A2(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(KEYINPUT111), .B1(new_n711_), .B2(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(G50gat), .B1(new_n709_), .B2(new_n698_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT111), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n716_), .B(new_n717_), .C1(new_n704_), .C2(new_n713_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n715_), .A2(new_n718_), .ZN(G1331gat));
  INV_X1    g518(.A(new_n315_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n287_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n616_), .A2(new_n721_), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n660_), .B(new_n720_), .C1(KEYINPUT112), .C2(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n723_), .B1(KEYINPUT112), .B2(new_n722_), .ZN(new_n724_));
  AOI21_X1  g523(.A(G57gat), .B1(new_n724_), .B2(new_n541_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n676_), .A2(new_n315_), .A3(new_n287_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(new_n608_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n542_), .A2(new_n208_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n725_), .B1(new_n727_), .B2(new_n728_), .ZN(G1332gat));
  NAND3_X1  g528(.A1(new_n724_), .A2(new_n209_), .A3(new_n624_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT48), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n727_), .A2(new_n624_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n732_), .B2(G64gat), .ZN(new_n733_));
  AOI211_X1 g532(.A(KEYINPUT48), .B(new_n209_), .C1(new_n727_), .C2(new_n624_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n730_), .B1(new_n733_), .B2(new_n734_), .ZN(G1333gat));
  NAND3_X1  g534(.A1(new_n724_), .A2(new_n217_), .A3(new_n508_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT49), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n727_), .A2(new_n508_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n738_), .B2(G71gat), .ZN(new_n739_));
  AOI211_X1 g538(.A(KEYINPUT49), .B(new_n217_), .C1(new_n727_), .C2(new_n508_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n736_), .B1(new_n739_), .B2(new_n740_), .ZN(G1334gat));
  NAND2_X1  g540(.A1(new_n562_), .A2(new_n218_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT113), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n724_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n727_), .A2(new_n562_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n746_), .B2(G78gat), .ZN(new_n747_));
  AOI211_X1 g546(.A(KEYINPUT50), .B(new_n218_), .C1(new_n727_), .C2(new_n562_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(G1335gat));
  AND2_X1   g548(.A1(new_n726_), .A2(new_n653_), .ZN(new_n750_));
  AOI21_X1  g549(.A(G85gat), .B1(new_n750_), .B2(new_n541_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n287_), .A2(new_n581_), .A3(new_n315_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n697_), .A2(new_n752_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n542_), .A2(new_n237_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n751_), .B1(new_n753_), .B2(new_n754_), .ZN(G1336gat));
  AOI21_X1  g554(.A(G92gat), .B1(new_n750_), .B2(new_n624_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n416_), .A2(new_n244_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n753_), .B2(new_n757_), .ZN(G1337gat));
  AOI21_X1  g557(.A(new_n257_), .B1(new_n753_), .B2(new_n508_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n726_), .A2(new_n252_), .A3(new_n508_), .A4(new_n653_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT114), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  OR3_X1    g563(.A1(new_n759_), .A2(new_n762_), .A3(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n759_), .B2(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(G1338gat));
  NAND3_X1  g566(.A1(new_n750_), .A2(new_n253_), .A3(new_n562_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n562_), .B(new_n752_), .C1(new_n661_), .C2(new_n663_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n769_), .A2(new_n770_), .A3(G106gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n769_), .B2(G106gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g573(.A1(new_n624_), .A2(new_n542_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n269_), .A2(new_n228_), .A3(new_n232_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n777_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n274_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n776_), .B(new_n203_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n271_), .A2(new_n204_), .A3(new_n274_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT55), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n282_), .B(new_n780_), .C1(new_n782_), .C2(new_n275_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT56), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n203_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n785_), .A2(KEYINPUT55), .A3(new_n781_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT56), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n786_), .A2(new_n787_), .A3(new_n282_), .A4(new_n780_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n309_), .A2(G229gat), .A3(G233gat), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n304_), .A2(new_n310_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  MUX2_X1   g590(.A(new_n311_), .B(new_n791_), .S(new_n314_), .Z(new_n792_));
  NAND4_X1  g591(.A1(new_n784_), .A2(new_n283_), .A3(new_n788_), .A4(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT58), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n615_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT117), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n793_), .A2(new_n794_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n795_), .A2(new_n800_), .A3(new_n615_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n797_), .A2(new_n799_), .A3(new_n801_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n784_), .A2(new_n315_), .A3(new_n788_), .A4(new_n283_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n283_), .A2(new_n284_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n792_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT57), .B1(new_n806_), .B2(new_n652_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808_));
  AOI211_X1 g607(.A(new_n808_), .B(new_n607_), .C1(new_n803_), .C2(new_n805_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n581_), .B1(new_n802_), .B2(new_n810_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n612_), .A2(new_n581_), .A3(new_n720_), .A4(new_n614_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(KEYINPUT116), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n812_), .A2(new_n721_), .A3(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(KEYINPUT116), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  OAI211_X1 g616(.A(KEYINPUT116), .B(new_n813_), .C1(new_n812_), .C2(new_n721_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n555_), .B(new_n775_), .C1(new_n811_), .C2(new_n819_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n820_), .A2(new_n564_), .ZN(new_n821_));
  AOI21_X1  g620(.A(G113gat), .B1(new_n821_), .B2(new_n315_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT59), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n820_), .B2(new_n564_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n795_), .A2(new_n800_), .A3(new_n615_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n800_), .B1(new_n795_), .B2(new_n615_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n825_), .A2(new_n826_), .A3(new_n798_), .ZN(new_n827_));
  OR2_X1    g626(.A1(new_n807_), .A2(new_n809_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n582_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n819_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n562_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n831_), .A2(KEYINPUT59), .A3(new_n508_), .A4(new_n775_), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n824_), .A2(new_n832_), .A3(KEYINPUT118), .ZN(new_n833_));
  AOI21_X1  g632(.A(KEYINPUT118), .B1(new_n824_), .B2(new_n832_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n315_), .A2(G113gat), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n822_), .B1(new_n835_), .B2(new_n836_), .ZN(G1340gat));
  NAND2_X1  g636(.A1(new_n824_), .A2(new_n832_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT60), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n839_), .B1(new_n287_), .B2(G120gat), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n821_), .A2(new_n840_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n838_), .A2(new_n721_), .A3(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(G120gat), .ZN(new_n843_));
  OAI22_X1  g642(.A1(new_n842_), .A2(new_n843_), .B1(KEYINPUT60), .B2(new_n841_), .ZN(G1341gat));
  AOI21_X1  g643(.A(G127gat), .B1(new_n821_), .B2(new_n581_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n581_), .A2(new_n846_), .A3(G127gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n846_), .B2(G127gat), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n845_), .B1(new_n835_), .B2(new_n848_), .ZN(G1342gat));
  AOI21_X1  g648(.A(G134gat), .B1(new_n821_), .B2(new_n607_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n615_), .A2(G134gat), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n850_), .B1(new_n835_), .B2(new_n851_), .ZN(G1343gat));
  OAI211_X1 g651(.A(new_n562_), .B(new_n564_), .C1(new_n811_), .C2(new_n819_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n775_), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT120), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n508_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n856_), .A2(new_n857_), .A3(new_n562_), .A4(new_n775_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n720_), .B1(new_n855_), .B2(new_n858_), .ZN(new_n859_));
  XOR2_X1   g658(.A(KEYINPUT121), .B(G141gat), .Z(new_n860_));
  XNOR2_X1  g659(.A(new_n859_), .B(new_n860_), .ZN(G1344gat));
  AOI21_X1  g660(.A(new_n287_), .B1(new_n855_), .B2(new_n858_), .ZN(new_n862_));
  INV_X1    g661(.A(G148gat), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(G1345gat));
  AOI21_X1  g663(.A(new_n582_), .B1(new_n855_), .B2(new_n858_), .ZN(new_n865_));
  XOR2_X1   g664(.A(KEYINPUT61), .B(G155gat), .Z(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1346gat));
  NAND2_X1  g666(.A1(new_n855_), .A2(new_n858_), .ZN(new_n868_));
  AOI21_X1  g667(.A(G162gat), .B1(new_n868_), .B2(new_n607_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n662_), .B1(new_n855_), .B2(new_n858_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(G162gat), .B2(new_n870_), .ZN(G1347gat));
  NOR2_X1   g670(.A1(new_n416_), .A2(new_n541_), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n514_), .B(new_n872_), .C1(new_n811_), .C2(new_n819_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(KEYINPUT123), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n874_), .A2(new_n315_), .A3(new_n338_), .A4(new_n341_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT62), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n876_), .B(G169gat), .C1(new_n873_), .C2(new_n720_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n873_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n315_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n876_), .B1(new_n881_), .B2(G169gat), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n875_), .B1(new_n879_), .B2(new_n882_), .ZN(G1348gat));
  NAND3_X1  g682(.A1(new_n880_), .A2(G176gat), .A3(new_n721_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(KEYINPUT124), .ZN(new_n885_));
  AOI21_X1  g684(.A(G176gat), .B1(new_n874_), .B2(new_n721_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1349gat));
  XOR2_X1   g686(.A(new_n873_), .B(KEYINPUT123), .Z(new_n888_));
  NOR3_X1   g687(.A1(new_n888_), .A2(new_n328_), .A3(new_n582_), .ZN(new_n889_));
  AOI21_X1  g688(.A(G183gat), .B1(new_n880_), .B2(new_n581_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1350gat));
  OAI21_X1  g690(.A(G190gat), .B1(new_n888_), .B2(new_n662_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n607_), .A2(new_n332_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(KEYINPUT125), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n892_), .B1(new_n888_), .B2(new_n894_), .ZN(G1351gat));
  INV_X1    g694(.A(new_n872_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n853_), .A2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n315_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n721_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n900_), .A2(KEYINPUT126), .A3(G204gat), .ZN(new_n901_));
  NAND3_X1  g700(.A1(KEYINPUT89), .A2(KEYINPUT126), .A3(G204gat), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n897_), .A2(new_n721_), .A3(new_n346_), .A4(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n903_), .ZN(G1353gat));
  NAND4_X1  g703(.A1(new_n856_), .A2(new_n562_), .A3(new_n581_), .A4(new_n872_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT63), .ZN(new_n906_));
  INV_X1    g705(.A(G211gat), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(KEYINPUT127), .B1(new_n905_), .B2(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT127), .ZN(new_n911_));
  INV_X1    g710(.A(new_n908_), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n897_), .A2(new_n911_), .A3(new_n581_), .A4(new_n912_), .ZN(new_n913_));
  AND3_X1   g712(.A1(new_n909_), .A2(new_n910_), .A3(new_n913_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n910_), .B1(new_n909_), .B2(new_n913_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1354gat));
  AOI21_X1  g715(.A(G218gat), .B1(new_n897_), .B2(new_n607_), .ZN(new_n917_));
  AND2_X1   g716(.A1(new_n615_), .A2(G218gat), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(new_n897_), .B2(new_n918_), .ZN(G1355gat));
endmodule


