//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n941_;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G78gat), .B(G106gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  XOR2_X1   g006(.A(new_n207_), .B(KEYINPUT3), .Z(new_n208_));
  NAND2_X1  g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  XOR2_X1   g008(.A(new_n209_), .B(KEYINPUT2), .Z(new_n210_));
  OAI211_X1 g009(.A(new_n204_), .B(new_n206_), .C1(new_n208_), .C2(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n205_), .B1(KEYINPUT1), .B2(new_n204_), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n212_), .B1(KEYINPUT1), .B2(new_n204_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n207_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(new_n214_), .A3(new_n209_), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n211_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT29), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G228gat), .ZN(new_n219_));
  INV_X1    g018(.A(G233gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n218_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G197gat), .B(G204gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G211gat), .B(G218gat), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n224_), .A2(new_n226_), .A3(KEYINPUT21), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n225_), .B1(new_n224_), .B2(KEYINPUT21), .ZN(new_n228_));
  INV_X1    g027(.A(G197gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(G204gat), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT21), .B1(new_n230_), .B2(KEYINPUT86), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n231_), .B1(KEYINPUT86), .B2(new_n223_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n227_), .B1(new_n228_), .B2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT87), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n222_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT88), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT88), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n222_), .A2(new_n237_), .A3(new_n234_), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n233_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n221_), .B1(new_n218_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n203_), .B1(new_n239_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n216_), .A2(new_n217_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT28), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G22gat), .B(G50gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n242_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n203_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n243_), .A2(new_n247_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT90), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT90), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n243_), .A2(new_n253_), .A3(new_n247_), .A4(new_n250_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n247_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT89), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n243_), .A2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n257_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(new_n250_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n256_), .B1(new_n258_), .B2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n255_), .A2(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(G127gat), .B(G134gat), .Z(new_n263_));
  XOR2_X1   g062(.A(G113gat), .B(G120gat), .Z(new_n264_));
  XOR2_X1   g063(.A(new_n263_), .B(new_n264_), .Z(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n216_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n211_), .A2(new_n215_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(new_n265_), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n267_), .A2(KEYINPUT4), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT94), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G225gat), .A2(G233gat), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n273_), .B1(new_n269_), .B2(KEYINPUT4), .ZN(new_n274_));
  OR3_X1    g073(.A1(new_n270_), .A2(new_n271_), .A3(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n271_), .B1(new_n270_), .B2(new_n274_), .ZN(new_n276_));
  AND2_X1   g075(.A1(new_n267_), .A2(new_n269_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n272_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n275_), .A2(new_n276_), .A3(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G1gat), .B(G29gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(G85gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT0), .B(G57gat), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n281_), .B(new_n282_), .Z(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n279_), .A2(new_n284_), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n275_), .A2(new_n283_), .A3(new_n276_), .A4(new_n278_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n262_), .A2(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(G8gat), .B(G36gat), .Z(new_n290_));
  XNOR2_X1  g089(.A(G64gat), .B(G92gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n293_));
  XOR2_X1   g092(.A(new_n292_), .B(new_n293_), .Z(new_n294_));
  INV_X1    g093(.A(new_n234_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT83), .ZN(new_n296_));
  INV_X1    g095(.A(G169gat), .ZN(new_n297_));
  INV_X1    g096(.A(G176gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n299_), .A2(KEYINPUT24), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT23), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n301_), .B1(G183gat), .B2(G190gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT79), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  AOI211_X1 g103(.A(KEYINPUT79), .B(new_n301_), .C1(G183gat), .C2(G190gat), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n301_), .A2(G183gat), .A3(G190gat), .ZN(new_n306_));
  NOR3_X1   g105(.A1(new_n304_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT24), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  AOI211_X1 g109(.A(new_n300_), .B(new_n307_), .C1(new_n299_), .C2(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(KEYINPUT77), .B(G183gat), .Z(new_n312_));
  INV_X1    g111(.A(KEYINPUT25), .ZN(new_n313_));
  OR3_X1    g112(.A1(new_n312_), .A2(KEYINPUT78), .A3(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT78), .B1(new_n312_), .B2(new_n313_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(G183gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT26), .B(G190gat), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n314_), .A2(new_n315_), .A3(new_n316_), .A4(new_n317_), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n311_), .A2(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n312_), .A2(G190gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n306_), .B(KEYINPUT82), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n302_), .B(KEYINPUT81), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n320_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  XOR2_X1   g122(.A(KEYINPUT22), .B(G169gat), .Z(new_n324_));
  AND2_X1   g123(.A1(new_n324_), .A2(KEYINPUT80), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n297_), .A2(KEYINPUT22), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n298_), .B1(new_n326_), .B2(KEYINPUT80), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n308_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n323_), .A2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n296_), .B1(new_n319_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n311_), .A2(new_n318_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n329_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n331_), .A2(new_n332_), .A3(KEYINPUT83), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n295_), .B1(new_n330_), .B2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G226gat), .A2(G233gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT19), .ZN(new_n336_));
  NOR2_X1   g135(.A1(G183gat), .A2(G190gat), .ZN(new_n337_));
  OAI221_X1 g136(.A(new_n308_), .B1(G176gat), .B2(new_n324_), .C1(new_n307_), .C2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n321_), .A2(new_n322_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n339_), .B1(KEYINPUT24), .B2(new_n299_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT25), .B(G183gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT91), .ZN(new_n342_));
  INV_X1    g141(.A(new_n317_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n310_), .A2(KEYINPUT92), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n299_), .B1(new_n310_), .B2(KEYINPUT92), .ZN(new_n345_));
  OAI22_X1  g144(.A1(new_n342_), .A2(new_n343_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n338_), .B1(new_n340_), .B2(new_n346_), .ZN(new_n347_));
  OR2_X1    g146(.A1(new_n347_), .A2(new_n233_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT20), .ZN(new_n349_));
  NOR3_X1   g148(.A1(new_n334_), .A2(new_n336_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n336_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n330_), .A2(new_n333_), .A3(new_n295_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT20), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n353_), .B1(new_n347_), .B2(new_n233_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n351_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n294_), .B1(new_n350_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n352_), .A2(new_n354_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(new_n336_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n294_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n333_), .ZN(new_n360_));
  AOI21_X1  g159(.A(KEYINPUT83), .B1(new_n331_), .B2(new_n332_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n234_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n349_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(new_n351_), .A3(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n358_), .A2(new_n359_), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT27), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n356_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT96), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n336_), .B1(new_n334_), .B2(new_n349_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n352_), .A2(new_n351_), .A3(new_n354_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n369_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n369_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n294_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT97), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n365_), .A2(new_n376_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n358_), .A2(KEYINPUT97), .A3(new_n364_), .A4(new_n359_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n375_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n368_), .B1(new_n379_), .B2(KEYINPUT27), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n202_), .B1(new_n289_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n377_), .A2(new_n378_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n352_), .A2(new_n351_), .A3(new_n354_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n351_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT96), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n359_), .B1(new_n385_), .B2(new_n373_), .ZN(new_n386_));
  OAI21_X1  g185(.A(KEYINPUT27), .B1(new_n382_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n367_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n287_), .B1(new_n255_), .B2(new_n261_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(KEYINPUT98), .A3(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT33), .ZN(new_n391_));
  OR2_X1    g190(.A1(new_n286_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n270_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n393_), .B(new_n272_), .C1(KEYINPUT4), .C2(new_n269_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n283_), .B1(new_n277_), .B2(new_n273_), .ZN(new_n395_));
  AOI22_X1  g194(.A1(new_n286_), .A2(new_n391_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n356_), .A2(new_n365_), .A3(new_n392_), .A4(new_n396_), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n397_), .A2(KEYINPUT95), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n359_), .A2(KEYINPUT32), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n399_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n358_), .A2(new_n364_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n400_), .B(new_n287_), .C1(new_n401_), .C2(new_n399_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n397_), .A2(KEYINPUT95), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n398_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n262_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n381_), .A2(new_n390_), .A3(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT84), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT31), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n408_), .B1(new_n266_), .B2(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n410_), .B1(new_n409_), .B2(new_n266_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G71gat), .B(G99gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(G43gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n411_), .B(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G227gat), .A2(G233gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(G15gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT30), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n414_), .B(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n330_), .A2(new_n333_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT85), .ZN(new_n421_));
  OR2_X1    g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n419_), .A2(new_n421_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n407_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n388_), .A2(new_n405_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n424_), .A2(new_n288_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n426_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT9), .ZN(new_n432_));
  INV_X1    g231(.A(G85gat), .ZN(new_n433_));
  INV_X1    g232(.A(G92gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G85gat), .A2(G92gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT65), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n432_), .B(new_n435_), .C1(new_n437_), .C2(new_n438_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n435_), .A2(KEYINPUT65), .A3(KEYINPUT9), .A4(new_n436_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G99gat), .A2(G106gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT6), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT6), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n443_), .A2(G99gat), .A3(G106gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  OR2_X1    g244(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n446_));
  INV_X1    g245(.A(G106gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n446_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n439_), .A2(new_n440_), .A3(new_n445_), .A4(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NOR3_X1   g251(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  AOI211_X1 g253(.A(KEYINPUT8), .B(new_n437_), .C1(new_n454_), .C2(new_n445_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT8), .ZN(new_n456_));
  OR3_X1    g255(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n443_), .B1(G99gat), .B2(G106gat), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n441_), .A2(KEYINPUT6), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n457_), .B(new_n451_), .C1(new_n458_), .C2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n437_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n456_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n450_), .B1(new_n455_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT66), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT66), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n465_), .B(new_n450_), .C1(new_n455_), .C2(new_n462_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(G64gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(G57gat), .ZN(new_n469_));
  INV_X1    g268(.A(G57gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(G64gat), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT67), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n469_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n472_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT11), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n470_), .A2(G64gat), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n468_), .A2(G57gat), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT67), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT11), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n469_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G71gat), .B(G78gat), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n475_), .A2(new_n481_), .A3(new_n483_), .ZN(new_n484_));
  OAI211_X1 g283(.A(KEYINPUT11), .B(new_n482_), .C1(new_n473_), .C2(new_n474_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT68), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT68), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n484_), .A2(new_n488_), .A3(new_n485_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n467_), .A2(new_n490_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n464_), .A2(new_n487_), .A3(new_n489_), .A4(new_n466_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n486_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n494_), .A2(KEYINPUT12), .A3(new_n463_), .ZN(new_n495_));
  AOI22_X1  g294(.A1(new_n464_), .A2(new_n466_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n492_), .B(new_n495_), .C1(new_n496_), .C2(KEYINPUT12), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G230gat), .A2(G233gat), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n498_), .B(KEYINPUT64), .Z(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  MUX2_X1   g299(.A(new_n493_), .B(new_n497_), .S(new_n500_), .Z(new_n501_));
  XNOR2_X1  g300(.A(G120gat), .B(G148gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT5), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G176gat), .B(G204gat), .ZN(new_n504_));
  XOR2_X1   g303(.A(new_n503_), .B(new_n504_), .Z(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(KEYINPUT69), .B1(new_n501_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n501_), .A2(new_n506_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n507_), .B1(new_n501_), .B2(new_n506_), .ZN(new_n511_));
  AND3_X1   g310(.A1(new_n510_), .A2(new_n511_), .A3(KEYINPUT13), .ZN(new_n512_));
  AOI21_X1  g311(.A(KEYINPUT13), .B1(new_n510_), .B2(new_n511_), .ZN(new_n513_));
  OR2_X1    g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT74), .B(G1gat), .ZN(new_n516_));
  INV_X1    g315(.A(G8gat), .ZN(new_n517_));
  OAI21_X1  g316(.A(KEYINPUT14), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G15gat), .B(G22gat), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G1gat), .B(G8gat), .ZN(new_n521_));
  OR2_X1    g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n521_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(G29gat), .B(G36gat), .Z(new_n525_));
  XOR2_X1   g324(.A(G43gat), .B(G50gat), .Z(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n524_), .A2(new_n527_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G229gat), .A2(G233gat), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n524_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n527_), .B(KEYINPUT15), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n536_), .A2(new_n529_), .A3(new_n531_), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n533_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G113gat), .B(G141gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G169gat), .B(G197gat), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n539_), .B(new_n540_), .Z(new_n541_));
  NAND2_X1  g340(.A1(new_n538_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT76), .ZN(new_n543_));
  INV_X1    g342(.A(new_n530_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n537_), .B1(new_n544_), .B2(new_n531_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n541_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n542_), .A2(new_n543_), .A3(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n545_), .A2(KEYINPUT76), .A3(new_n546_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n515_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n431_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G231gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n524_), .B(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n490_), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n556_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G127gat), .B(G155gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT16), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G183gat), .B(G211gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT17), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n557_), .A2(new_n558_), .A3(new_n563_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n555_), .A2(new_n494_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n555_), .A2(new_n494_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT17), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n562_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n565_), .A2(new_n566_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n564_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT75), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT34), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT35), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT70), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  AOI22_X1  g377(.A1(new_n535_), .A2(new_n463_), .B1(new_n575_), .B2(new_n574_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n464_), .A2(new_n527_), .A3(new_n466_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n578_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n576_), .A2(new_n577_), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n582_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(G134gat), .B(G162gat), .Z(new_n586_));
  XNOR2_X1  g385(.A(G190gat), .B(G218gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT36), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n590_), .B(KEYINPUT71), .Z(new_n591_));
  NAND2_X1  g390(.A1(new_n585_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT72), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n588_), .A2(new_n589_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n583_), .A2(new_n584_), .A3(new_n590_), .A4(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n594_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n597_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NOR3_X1   g400(.A1(new_n553_), .A2(new_n571_), .A3(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n602_), .A2(new_n516_), .A3(new_n287_), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n603_), .A2(KEYINPUT99), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(KEYINPUT99), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT38), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n604_), .A2(KEYINPUT38), .A3(new_n605_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n594_), .A2(new_n596_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n611_), .A2(new_n571_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n431_), .A2(new_n552_), .A3(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G1gat), .B1(new_n613_), .B2(new_n288_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n608_), .A2(new_n609_), .A3(new_n614_), .ZN(G1324gat));
  NAND3_X1  g414(.A1(new_n602_), .A2(new_n517_), .A3(new_n380_), .ZN(new_n616_));
  OAI21_X1  g415(.A(G8gat), .B1(new_n613_), .B2(new_n388_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n617_), .A2(KEYINPUT39), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(KEYINPUT39), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n616_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g420(.A(G15gat), .B1(new_n613_), .B2(new_n425_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT41), .Z(new_n623_));
  INV_X1    g422(.A(G15gat), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n602_), .A2(new_n624_), .A3(new_n424_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(G1326gat));
  OAI21_X1  g425(.A(G22gat), .B1(new_n613_), .B2(new_n405_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT42), .ZN(new_n628_));
  INV_X1    g427(.A(G22gat), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n602_), .A2(new_n629_), .A3(new_n262_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(G1327gat));
  NAND2_X1  g430(.A1(new_n611_), .A2(new_n571_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n553_), .A2(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(G29gat), .B1(new_n633_), .B2(new_n287_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n552_), .A2(new_n571_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT43), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n637_), .B1(new_n431_), .B2(new_n601_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n429_), .B1(new_n407_), .B2(new_n425_), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n639_), .A2(KEYINPUT43), .A3(new_n600_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n636_), .B1(new_n638_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT44), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n641_), .A2(KEYINPUT100), .A3(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n388_), .A2(new_n389_), .ZN(new_n645_));
  AOI22_X1  g444(.A1(new_n645_), .A2(new_n202_), .B1(new_n405_), .B2(new_n404_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n424_), .B1(new_n646_), .B2(new_n390_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n637_), .B(new_n601_), .C1(new_n647_), .C2(new_n429_), .ZN(new_n648_));
  OAI21_X1  g447(.A(KEYINPUT43), .B1(new_n639_), .B2(new_n600_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n635_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n644_), .B1(new_n650_), .B2(KEYINPUT44), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n643_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(KEYINPUT44), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n287_), .A2(G29gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n634_), .B1(new_n655_), .B2(new_n656_), .ZN(G1328gat));
  INV_X1    g456(.A(KEYINPUT46), .ZN(new_n658_));
  INV_X1    g457(.A(G36gat), .ZN(new_n659_));
  AOI211_X1 g458(.A(new_n642_), .B(new_n635_), .C1(new_n648_), .C2(new_n649_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n660_), .A2(new_n388_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n659_), .B1(new_n652_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT45), .ZN(new_n663_));
  INV_X1    g462(.A(new_n632_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n388_), .A2(G36gat), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n431_), .A2(new_n552_), .A3(new_n664_), .A4(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT101), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n666_), .A2(KEYINPUT101), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n663_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n669_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n671_), .A2(KEYINPUT45), .A3(new_n667_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n658_), .B1(new_n662_), .B2(new_n673_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n670_), .A2(new_n672_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n653_), .A2(new_n380_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n676_), .B1(new_n651_), .B2(new_n643_), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n675_), .B(KEYINPUT46), .C1(new_n677_), .C2(new_n659_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n674_), .A2(new_n678_), .ZN(G1329gat));
  NAND2_X1  g478(.A1(new_n424_), .A2(G43gat), .ZN(new_n680_));
  AOI211_X1 g479(.A(new_n660_), .B(new_n680_), .C1(new_n643_), .C2(new_n651_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n553_), .A2(new_n425_), .A3(new_n632_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n682_), .A2(G43gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(KEYINPUT47), .B1(new_n681_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT47), .ZN(new_n685_));
  INV_X1    g484(.A(new_n683_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n685_), .B(new_n686_), .C1(new_n654_), .C2(new_n680_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n684_), .A2(new_n687_), .ZN(G1330gat));
  INV_X1    g487(.A(G50gat), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n633_), .A2(new_n689_), .A3(new_n262_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n405_), .B1(new_n650_), .B2(KEYINPUT44), .ZN(new_n691_));
  AOI211_X1 g490(.A(KEYINPUT102), .B(new_n689_), .C1(new_n652_), .C2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT102), .ZN(new_n693_));
  AOI21_X1  g492(.A(KEYINPUT100), .B1(new_n641_), .B2(new_n642_), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n650_), .A2(new_n644_), .A3(KEYINPUT44), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n691_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n693_), .B1(new_n696_), .B2(G50gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n690_), .B1(new_n692_), .B2(new_n697_), .ZN(G1331gat));
  INV_X1    g497(.A(new_n571_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n515_), .A2(new_n600_), .A3(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n551_), .B1(new_n700_), .B2(KEYINPUT103), .ZN(new_n701_));
  AOI211_X1 g500(.A(new_n701_), .B(new_n639_), .C1(KEYINPUT103), .C2(new_n700_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n702_), .A2(new_n470_), .A3(new_n287_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n514_), .A2(new_n550_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n431_), .A2(new_n612_), .A3(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(G57gat), .B1(new_n705_), .B2(new_n288_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n703_), .A2(new_n706_), .ZN(G1332gat));
  OAI21_X1  g506(.A(G64gat), .B1(new_n705_), .B2(new_n388_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT48), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n380_), .A2(new_n468_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT104), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n702_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n709_), .A2(new_n712_), .ZN(G1333gat));
  OAI21_X1  g512(.A(G71gat), .B1(new_n705_), .B2(new_n425_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT49), .ZN(new_n715_));
  INV_X1    g514(.A(G71gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n702_), .A2(new_n716_), .A3(new_n424_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(G1334gat));
  OAI21_X1  g517(.A(G78gat), .B1(new_n705_), .B2(new_n405_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT50), .ZN(new_n720_));
  INV_X1    g519(.A(G78gat), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n702_), .A2(new_n721_), .A3(new_n262_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1335gat));
  NOR4_X1   g522(.A1(new_n639_), .A2(new_n550_), .A3(new_n514_), .A4(new_n632_), .ZN(new_n724_));
  AOI21_X1  g523(.A(G85gat), .B1(new_n724_), .B2(new_n287_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n704_), .A2(new_n571_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n726_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT105), .Z(new_n728_));
  NOR2_X1   g527(.A1(new_n288_), .A2(new_n433_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(G1336gat));
  AOI21_X1  g529(.A(G92gat), .B1(new_n724_), .B2(new_n380_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT106), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n388_), .A2(new_n434_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n728_), .B2(new_n733_), .ZN(G1337gat));
  NAND2_X1  g533(.A1(new_n727_), .A2(new_n424_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(G99gat), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n424_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n738_));
  AOI22_X1  g537(.A1(new_n724_), .A2(new_n737_), .B1(new_n738_), .B2(KEYINPUT51), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n736_), .A2(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n738_), .A2(KEYINPUT51), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n740_), .B(new_n741_), .Z(G1338gat));
  NAND3_X1  g541(.A1(new_n724_), .A2(new_n447_), .A3(new_n262_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT52), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n727_), .A2(new_n262_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n745_), .B2(G106gat), .ZN(new_n746_));
  AOI211_X1 g545(.A(KEYINPUT52), .B(new_n447_), .C1(new_n727_), .C2(new_n262_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n743_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g548(.A1(new_n427_), .A2(new_n288_), .A3(new_n425_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT59), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT54), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n571_), .A2(new_n550_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n514_), .A2(KEYINPUT108), .A3(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n754_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT108), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n755_), .A2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n753_), .B1(new_n759_), .B2(new_n600_), .ZN(new_n760_));
  AOI211_X1 g559(.A(KEYINPUT54), .B(new_n601_), .C1(new_n755_), .C2(new_n758_), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n536_), .A2(new_n529_), .A3(new_n532_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n541_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n764_));
  AOI22_X1  g563(.A1(new_n538_), .A2(new_n541_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n510_), .A2(new_n511_), .A3(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n501_), .A2(new_n506_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n550_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n492_), .A2(new_n495_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT12), .B1(new_n467_), .B2(new_n490_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n499_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n497_), .A2(KEYINPUT109), .A3(new_n499_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(KEYINPUT55), .B1(new_n497_), .B2(new_n499_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n771_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n772_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n779_), .A2(new_n780_), .A3(new_n781_), .A4(new_n500_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n778_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n777_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT110), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT110), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n777_), .A2(new_n783_), .A3(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT56), .B1(new_n788_), .B2(new_n505_), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n777_), .A2(new_n783_), .A3(new_n786_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n786_), .B1(new_n777_), .B2(new_n783_), .ZN(new_n791_));
  OAI211_X1 g590(.A(KEYINPUT56), .B(new_n505_), .C1(new_n790_), .C2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n770_), .B1(new_n789_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n767_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n505_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT56), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n769_), .B1(new_n799_), .B2(new_n792_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT111), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n611_), .B1(new_n796_), .B2(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n802_), .A2(KEYINPUT57), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n766_), .B1(new_n800_), .B2(KEYINPUT111), .ZN(new_n804_));
  AOI211_X1 g603(.A(new_n795_), .B(new_n769_), .C1(new_n799_), .C2(new_n792_), .ZN(new_n805_));
  OAI211_X1 g604(.A(KEYINPUT57), .B(new_n610_), .C1(new_n804_), .C2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n768_), .A2(new_n765_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n799_), .B2(new_n792_), .ZN(new_n808_));
  OR2_X1    g607(.A1(new_n808_), .A2(KEYINPUT58), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(KEYINPUT58), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(new_n601_), .A3(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n806_), .A2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n571_), .B1(new_n803_), .B2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n752_), .B1(new_n762_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n760_), .A2(new_n761_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n806_), .A2(new_n811_), .ZN(new_n817_));
  OAI21_X1  g616(.A(KEYINPUT112), .B1(new_n802_), .B2(KEYINPUT57), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n610_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT112), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n819_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n817_), .A2(new_n818_), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n816_), .B1(new_n823_), .B2(new_n571_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n750_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n815_), .B1(new_n826_), .B2(new_n751_), .ZN(new_n827_));
  OAI21_X1  g626(.A(G113gat), .B1(new_n827_), .B2(new_n551_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n820_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n829_), .A2(new_n812_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n699_), .B1(new_n830_), .B2(new_n822_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n750_), .B1(new_n831_), .B2(new_n816_), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n551_), .A2(G113gat), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n828_), .B1(new_n832_), .B2(new_n833_), .ZN(G1340gat));
  INV_X1    g633(.A(KEYINPUT113), .ZN(new_n835_));
  INV_X1    g634(.A(G120gat), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n814_), .B1(new_n832_), .B2(KEYINPUT59), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(new_n515_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n514_), .A2(KEYINPUT60), .ZN(new_n839_));
  MUX2_X1   g638(.A(KEYINPUT60), .B(new_n839_), .S(new_n836_), .Z(new_n840_));
  NAND2_X1  g639(.A1(new_n826_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n835_), .B1(new_n838_), .B2(new_n842_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n515_), .B(new_n815_), .C1(new_n826_), .C2(new_n751_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(G120gat), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n845_), .A2(KEYINPUT113), .A3(new_n841_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n843_), .A2(new_n846_), .ZN(G1341gat));
  OAI21_X1  g646(.A(G127gat), .B1(new_n827_), .B2(new_n571_), .ZN(new_n848_));
  OR2_X1    g647(.A1(new_n571_), .A2(G127gat), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n832_), .B2(new_n849_), .ZN(G1342gat));
  INV_X1    g649(.A(G134gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n832_), .B2(new_n610_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n600_), .A2(new_n851_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(KEYINPUT114), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n852_), .B1(new_n827_), .B2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(KEYINPUT115), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT115), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n852_), .B(new_n858_), .C1(new_n827_), .C2(new_n855_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(G1343gat));
  NAND4_X1  g659(.A1(new_n388_), .A2(new_n262_), .A3(new_n287_), .A4(new_n425_), .ZN(new_n861_));
  XOR2_X1   g660(.A(new_n861_), .B(KEYINPUT116), .Z(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n824_), .A2(KEYINPUT117), .A3(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT117), .B1(new_n824_), .B2(new_n863_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n551_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT118), .B(G141gat), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(G1344gat));
  INV_X1    g668(.A(new_n866_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n515_), .B1(new_n870_), .B2(new_n864_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G148gat), .ZN(G1345gat));
  AOI21_X1  g671(.A(new_n571_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n873_));
  XOR2_X1   g672(.A(KEYINPUT61), .B(G155gat), .Z(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(KEYINPUT119), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(KEYINPUT120), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n873_), .B(new_n876_), .ZN(G1346gat));
  INV_X1    g676(.A(G162gat), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n878_), .B(new_n611_), .C1(new_n870_), .C2(new_n864_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n600_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(new_n878_), .ZN(G1347gat));
  NAND2_X1  g680(.A1(new_n762_), .A2(new_n813_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n388_), .A2(new_n428_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n262_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n882_), .A2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n550_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n297_), .B1(new_n888_), .B2(KEYINPUT121), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n886_), .A2(new_n551_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n889_), .A2(KEYINPUT62), .A3(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n894_));
  INV_X1    g693(.A(new_n892_), .ZN(new_n895_));
  OAI21_X1  g694(.A(G169gat), .B1(new_n890_), .B2(new_n891_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n894_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n897_));
  OR2_X1    g696(.A1(new_n888_), .A2(new_n324_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n893_), .A2(new_n897_), .A3(new_n898_), .ZN(G1348gat));
  AOI21_X1  g698(.A(G176gat), .B1(new_n887_), .B2(new_n515_), .ZN(new_n900_));
  OR2_X1    g699(.A1(new_n900_), .A2(KEYINPUT122), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(KEYINPUT122), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n903_), .B1(new_n824_), .B2(new_n262_), .ZN(new_n904_));
  OAI211_X1 g703(.A(KEYINPUT123), .B(new_n405_), .C1(new_n831_), .C2(new_n816_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n884_), .A2(new_n298_), .A3(new_n514_), .ZN(new_n907_));
  AOI22_X1  g706(.A1(new_n901_), .A2(new_n902_), .B1(new_n906_), .B2(new_n907_), .ZN(G1349gat));
  NAND3_X1  g707(.A1(new_n887_), .A2(new_n342_), .A3(new_n699_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n883_), .A2(new_n699_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n910_), .B1(new_n904_), .B2(new_n905_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n909_), .B1(new_n911_), .B2(new_n312_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(KEYINPUT124), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n914_));
  OAI211_X1 g713(.A(new_n914_), .B(new_n909_), .C1(new_n911_), .C2(new_n312_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n913_), .A2(new_n915_), .ZN(G1350gat));
  OAI21_X1  g715(.A(G190gat), .B1(new_n886_), .B2(new_n600_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n611_), .A2(new_n317_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n886_), .B2(new_n918_), .ZN(G1351gat));
  INV_X1    g718(.A(new_n824_), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n388_), .A2(new_n289_), .A3(new_n424_), .ZN(new_n921_));
  AND2_X1   g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  NAND4_X1  g721(.A1(new_n922_), .A2(KEYINPUT125), .A3(G197gat), .A4(new_n550_), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT125), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n920_), .A2(new_n550_), .A3(new_n921_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n925_), .B2(new_n229_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n925_), .A2(new_n229_), .ZN(new_n927_));
  AND3_X1   g726(.A1(new_n923_), .A2(new_n926_), .A3(new_n927_), .ZN(G1352gat));
  AND2_X1   g727(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n929_));
  NOR2_X1   g728(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n930_));
  OAI211_X1 g729(.A(new_n922_), .B(new_n515_), .C1(new_n929_), .C2(new_n930_), .ZN(new_n931_));
  AND2_X1   g730(.A1(new_n922_), .A2(new_n515_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n932_), .B2(new_n930_), .ZN(G1353gat));
  AOI21_X1  g732(.A(new_n571_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(KEYINPUT127), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n922_), .A2(new_n935_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  XOR2_X1   g736(.A(new_n936_), .B(new_n937_), .Z(G1354gat));
  INV_X1    g737(.A(G218gat), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n922_), .A2(new_n939_), .A3(new_n611_), .ZN(new_n940_));
  AND2_X1   g739(.A1(new_n922_), .A2(new_n601_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n940_), .B1(new_n941_), .B2(new_n939_), .ZN(G1355gat));
endmodule


