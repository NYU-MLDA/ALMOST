//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 0 0 0 1 0 1 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n899_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT0), .ZN(new_n203_));
  INV_X1    g002(.A(G57gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G85gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT1), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n210_), .B1(G155gat), .B2(G162gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n209_), .A2(KEYINPUT1), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G141gat), .ZN(new_n214_));
  INV_X1    g013(.A(G148gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217_));
  NOR3_X1   g016(.A1(new_n213_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  XOR2_X1   g018(.A(G155gat), .B(G162gat), .Z(new_n220_));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n217_), .A2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n222_), .B(new_n223_), .C1(new_n216_), .C2(KEYINPUT2), .ZN(new_n224_));
  NAND3_X1  g023(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT88), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n220_), .B1(new_n224_), .B2(new_n226_), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n227_), .A2(KEYINPUT89), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(KEYINPUT89), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n219_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT90), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT90), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n232_), .B(new_n219_), .C1(new_n228_), .C2(new_n229_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT4), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G127gat), .B(G134gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G113gat), .B(G120gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n231_), .A2(new_n233_), .A3(new_n234_), .A4(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT98), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G225gat), .A2(G233gat), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n231_), .A2(new_n238_), .A3(new_n233_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n229_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n227_), .A2(KEYINPUT89), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n218_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(new_n237_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n243_), .A2(KEYINPUT4), .A3(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n240_), .A2(new_n242_), .A3(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n243_), .A2(new_n241_), .A3(new_n247_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n208_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT98), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n239_), .B(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n248_), .A2(new_n242_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n250_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n255_), .A2(new_n207_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n251_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT103), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT96), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT21), .ZN(new_n260_));
  INV_X1    g059(.A(G218gat), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n261_), .A2(G211gat), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(G211gat), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n260_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G211gat), .B(G218gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT21), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G197gat), .B(G204gat), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n264_), .A2(new_n266_), .A3(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n265_), .A2(new_n267_), .A3(KEYINPUT21), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(G183gat), .ZN(new_n273_));
  INV_X1    g072(.A(G190gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT23), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT83), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT23), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n277_), .A2(G183gat), .A3(G190gat), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n275_), .A2(new_n276_), .A3(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n273_), .A2(new_n274_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n277_), .A2(KEYINPUT83), .A3(G183gat), .A4(G190gat), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283_));
  INV_X1    g082(.A(G169gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT22), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT22), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(G169gat), .ZN(new_n287_));
  INV_X1    g086(.A(G176gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n285_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n282_), .A2(new_n283_), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT82), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n283_), .A2(KEYINPUT24), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n284_), .A2(new_n288_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT26), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT81), .B1(new_n295_), .B2(G190gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n273_), .A2(KEYINPUT25), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT25), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(G183gat), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n296_), .A2(new_n297_), .A3(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n274_), .A2(KEYINPUT26), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n295_), .A2(G190gat), .ZN(new_n302_));
  AOI21_X1  g101(.A(KEYINPUT81), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n291_), .B(new_n294_), .C1(new_n300_), .C2(new_n303_), .ZN(new_n304_));
  NOR3_X1   g103(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n305_), .B1(new_n275_), .B2(new_n278_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT25), .B(G183gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT26), .B(G190gat), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n296_), .B(new_n308_), .C1(new_n309_), .C2(KEYINPUT81), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n291_), .B1(new_n310_), .B2(new_n294_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n290_), .B1(new_n307_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT84), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT84), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n314_), .B(new_n290_), .C1(new_n307_), .C2(new_n311_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n272_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT95), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n305_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n301_), .A2(new_n302_), .A3(new_n297_), .A4(new_n299_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n318_), .A2(new_n279_), .A3(new_n281_), .A4(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT94), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n289_), .A2(new_n321_), .A3(new_n283_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n278_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n277_), .B1(G183gat), .B2(G190gat), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n280_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n322_), .A2(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n321_), .B1(new_n289_), .B2(new_n283_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n320_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n317_), .B1(new_n328_), .B2(new_n271_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n327_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n330_), .A2(new_n322_), .A3(new_n325_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n272_), .A2(new_n331_), .A3(KEYINPUT95), .A4(new_n320_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G226gat), .A2(G233gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n336_), .A2(KEYINPUT20), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n329_), .A2(new_n332_), .A3(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n259_), .B1(new_n316_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n315_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n294_), .B1(new_n300_), .B2(new_n303_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT82), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(new_n304_), .A3(new_n306_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n314_), .B1(new_n343_), .B2(new_n290_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n271_), .B1(new_n340_), .B2(new_n344_), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n329_), .A2(new_n332_), .A3(new_n337_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(KEYINPUT96), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n339_), .A2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n271_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n328_), .A2(new_n272_), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT20), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(new_n335_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G8gat), .B(G36gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT18), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G64gat), .B(G92gat), .ZN(new_n355_));
  XOR2_X1   g154(.A(new_n354_), .B(new_n355_), .Z(new_n356_));
  AND4_X1   g155(.A1(KEYINPUT97), .A2(new_n348_), .A3(new_n352_), .A4(new_n356_), .ZN(new_n357_));
  AOI22_X1  g156(.A1(new_n339_), .A2(new_n347_), .B1(new_n351_), .B2(new_n335_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT97), .B1(new_n358_), .B2(new_n356_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n356_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n357_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(KEYINPUT102), .B(KEYINPUT27), .Z(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n258_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n358_), .A2(KEYINPUT97), .A3(new_n356_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT97), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n348_), .A2(new_n352_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n356_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n366_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n367_), .A2(new_n368_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n365_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n371_), .A2(KEYINPUT103), .A3(new_n362_), .ZN(new_n372_));
  OAI211_X1 g171(.A(KEYINPUT20), .B(new_n336_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT100), .B(KEYINPUT20), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n271_), .B(KEYINPUT92), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n374_), .B1(new_n375_), .B2(new_n328_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n335_), .B1(new_n316_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n373_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(new_n368_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n360_), .A2(KEYINPUT27), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT101), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT101), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n360_), .A2(new_n382_), .A3(KEYINPUT27), .A4(new_n379_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  AND4_X1   g183(.A1(new_n257_), .A2(new_n364_), .A3(new_n372_), .A4(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G22gat), .B(G50gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT91), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n272_), .B1(G228gat), .B2(G233gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n231_), .A2(new_n233_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT29), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n389_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n375_), .B1(new_n246_), .B2(new_n391_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n393_), .A2(G228gat), .A3(G233gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G78gat), .B(G106gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n396_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n392_), .A2(new_n394_), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n390_), .A2(new_n391_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT28), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT28), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n390_), .A2(new_n402_), .A3(new_n391_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n397_), .A2(new_n399_), .A3(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n404_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n388_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n397_), .A2(new_n399_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n404_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n397_), .A2(new_n404_), .A3(new_n399_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(new_n387_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n407_), .A2(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(KEYINPUT30), .B1(new_n340_), .B2(new_n344_), .ZN(new_n414_));
  XOR2_X1   g213(.A(G71gat), .B(G99gat), .Z(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(G43gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G227gat), .A2(G233gat), .ZN(new_n417_));
  INV_X1    g216(.A(G15gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  XOR2_X1   g218(.A(new_n416_), .B(new_n419_), .Z(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT30), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n313_), .A2(new_n422_), .A3(new_n315_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n414_), .A2(new_n421_), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n414_), .A2(new_n423_), .ZN(new_n425_));
  AOI21_X1  g224(.A(KEYINPUT85), .B1(new_n425_), .B2(new_n420_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT85), .ZN(new_n427_));
  AOI211_X1 g226(.A(new_n427_), .B(new_n421_), .C1(new_n414_), .C2(new_n423_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n424_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT86), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n313_), .A2(new_n422_), .A3(new_n315_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n422_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n420_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n427_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n425_), .A2(KEYINPUT85), .A3(new_n420_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT86), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n437_), .A3(new_n424_), .ZN(new_n438_));
  XOR2_X1   g237(.A(new_n237_), .B(KEYINPUT31), .Z(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n430_), .A2(new_n438_), .A3(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n440_), .B1(new_n430_), .B2(new_n438_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT87), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n437_), .B1(new_n436_), .B2(new_n424_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n424_), .ZN(new_n445_));
  AOI211_X1 g244(.A(KEYINPUT86), .B(new_n445_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n439_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT87), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n430_), .A2(new_n438_), .A3(new_n440_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n413_), .B1(new_n443_), .B2(new_n450_), .ZN(new_n451_));
  AOI22_X1  g250(.A1(new_n407_), .A2(new_n412_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n385_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n443_), .A2(new_n450_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n378_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n356_), .A2(KEYINPUT32), .ZN(new_n456_));
  MUX2_X1   g255(.A(new_n455_), .B(new_n367_), .S(new_n456_), .Z(new_n457_));
  OAI21_X1  g256(.A(new_n457_), .B1(new_n251_), .B2(new_n256_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT33), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n459_), .B1(new_n255_), .B2(new_n207_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n240_), .A2(new_n241_), .A3(new_n248_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n243_), .A2(new_n242_), .A3(new_n247_), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n462_), .A2(KEYINPUT99), .A3(new_n207_), .ZN(new_n463_));
  AOI21_X1  g262(.A(KEYINPUT99), .B1(new_n462_), .B2(new_n207_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n461_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n249_), .A2(KEYINPUT33), .A3(new_n250_), .A4(new_n208_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n460_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n458_), .B1(new_n467_), .B2(new_n371_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n454_), .A2(new_n413_), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n453_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G1gat), .B(G8gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(KEYINPUT76), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G15gat), .B(G22gat), .ZN(new_n474_));
  INV_X1    g273(.A(G1gat), .ZN(new_n475_));
  INV_X1    g274(.A(G8gat), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT14), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n474_), .A2(new_n477_), .ZN(new_n478_));
  OR2_X1    g277(.A1(new_n473_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n473_), .A2(new_n478_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G29gat), .B(G36gat), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G43gat), .B(G50gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n484_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n482_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n481_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT79), .ZN(new_n490_));
  INV_X1    g289(.A(new_n488_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n479_), .A2(new_n491_), .A3(new_n480_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n489_), .A2(new_n490_), .A3(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G229gat), .A2(G233gat), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n481_), .A2(KEYINPUT79), .A3(new_n488_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n493_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT80), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n493_), .A2(KEYINPUT80), .A3(new_n495_), .A4(new_n496_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT15), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n488_), .B(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n481_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n503_), .A2(new_n494_), .A3(new_n492_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n499_), .A2(new_n500_), .A3(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G113gat), .B(G141gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G169gat), .B(G197gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n505_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n508_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n499_), .A2(new_n500_), .A3(new_n504_), .A4(new_n510_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(G127gat), .B(G155gat), .Z(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT16), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G183gat), .B(G211gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT17), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G231gat), .A2(G233gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n481_), .B(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT66), .B(G71gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(G78gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G57gat), .B(G64gat), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n523_), .A2(KEYINPUT11), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(KEYINPUT11), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n522_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(G78gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n521_), .B(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n525_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n520_), .A2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n520_), .A2(new_n532_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n518_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT77), .ZN(new_n536_));
  NOR3_X1   g335(.A1(new_n516_), .A2(new_n536_), .A3(new_n517_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n535_), .B(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G190gat), .B(G218gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G134gat), .B(G162gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n541_), .B(KEYINPUT36), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT75), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT8), .ZN(new_n544_));
  AND2_X1   g343(.A1(G85gat), .A2(G92gat), .ZN(new_n545_));
  NOR2_X1   g344(.A1(G85gat), .A2(G92gat), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT65), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(G92gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n206_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT65), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G85gat), .A2(G92gat), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n549_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n547_), .A2(new_n552_), .A3(KEYINPUT64), .ZN(new_n553_));
  INV_X1    g352(.A(G99gat), .ZN(new_n554_));
  INV_X1    g353(.A(G106gat), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n554_), .A2(new_n555_), .A3(KEYINPUT7), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT7), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n557_), .B1(G99gat), .B2(G106gat), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  AND3_X1   g358(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n560_));
  AOI21_X1  g359(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n559_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n547_), .A2(new_n552_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n544_), .B(new_n553_), .C1(new_n563_), .C2(new_n564_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n547_), .A2(new_n552_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n559_), .A2(new_n562_), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n566_), .B(new_n567_), .C1(KEYINPUT64), .C2(KEYINPUT8), .ZN(new_n568_));
  OR2_X1    g367(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n569_), .A2(new_n555_), .A3(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n549_), .A2(KEYINPUT9), .A3(new_n551_), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n551_), .A2(KEYINPUT9), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n562_), .A2(new_n571_), .A3(new_n572_), .A4(new_n573_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n565_), .A2(new_n568_), .A3(new_n491_), .A4(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT73), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G232gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(KEYINPUT72), .B(KEYINPUT35), .Z(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n574_), .B(KEYINPUT67), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n585_), .A2(new_n568_), .A3(new_n565_), .ZN(new_n586_));
  AOI22_X1  g385(.A1(new_n586_), .A2(new_n502_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n577_), .A2(new_n584_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n584_), .B1(new_n577_), .B2(new_n587_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n543_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n590_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n541_), .A2(KEYINPUT36), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n592_), .A2(new_n593_), .A3(new_n588_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n591_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n591_), .A2(KEYINPUT74), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n595_), .A2(new_n596_), .A3(KEYINPUT37), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT37), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n591_), .B(new_n594_), .C1(KEYINPUT74), .C2(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n538_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT12), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n602_), .B1(new_n527_), .B2(new_n530_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n565_), .A2(new_n568_), .A3(new_n574_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  AOI22_X1  g404(.A1(new_n586_), .A2(new_n603_), .B1(new_n605_), .B2(new_n532_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(G230gat), .A2(G233gat), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n604_), .A2(new_n531_), .ZN(new_n608_));
  AOI21_X1  g407(.A(KEYINPUT68), .B1(new_n608_), .B2(new_n602_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT68), .ZN(new_n610_));
  AOI211_X1 g409(.A(new_n610_), .B(KEYINPUT12), .C1(new_n604_), .C2(new_n531_), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n606_), .B(new_n607_), .C1(new_n609_), .C2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n604_), .B(new_n531_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n613_), .A2(G230gat), .A3(G233gat), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G120gat), .B(G148gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT5), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT69), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G176gat), .B(G204gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n615_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n612_), .A2(new_n614_), .A3(new_n620_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT70), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n625_), .A2(KEYINPUT13), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(KEYINPUT13), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n624_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n622_), .A2(new_n625_), .A3(KEYINPUT13), .A4(new_n623_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n601_), .A2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT78), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n471_), .A2(new_n512_), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n257_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n634_), .A2(new_n475_), .A3(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT38), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n595_), .B(KEYINPUT104), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n631_), .A2(new_n512_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n641_), .A2(new_n538_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n470_), .A2(new_n639_), .A3(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G1gat), .B1(new_n643_), .B2(new_n257_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT105), .Z(new_n645_));
  NAND2_X1  g444(.A1(new_n637_), .A2(new_n645_), .ZN(G1324gat));
  AND2_X1   g445(.A1(new_n372_), .A2(new_n384_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n647_), .A2(new_n364_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n634_), .A2(new_n476_), .A3(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n643_), .A2(new_n648_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n476_), .B1(new_n651_), .B2(KEYINPUT106), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT39), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT106), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n654_), .B1(new_n643_), .B2(new_n648_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n652_), .A2(new_n653_), .A3(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n653_), .B1(new_n652_), .B2(new_n655_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n650_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT40), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  OAI211_X1 g459(.A(KEYINPUT40), .B(new_n650_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1325gat));
  INV_X1    g461(.A(new_n454_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n634_), .A2(new_n418_), .A3(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT107), .ZN(new_n665_));
  INV_X1    g464(.A(new_n643_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n418_), .B1(new_n666_), .B2(new_n663_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n668_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n665_), .A2(new_n669_), .A3(new_n670_), .ZN(G1326gat));
  INV_X1    g470(.A(G22gat), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n407_), .A2(new_n412_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n634_), .A2(new_n672_), .A3(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n666_), .A2(new_n673_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n676_), .B2(G22gat), .ZN(new_n677_));
  AOI211_X1 g476(.A(KEYINPUT42), .B(new_n672_), .C1(new_n666_), .C2(new_n673_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n674_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT108), .ZN(G1327gat));
  INV_X1    g479(.A(new_n538_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n681_), .A2(new_n595_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n471_), .A2(new_n641_), .A3(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(G29gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n684_), .A2(new_n685_), .A3(new_n635_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n597_), .A2(new_n599_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n364_), .A2(new_n372_), .A3(new_n384_), .A4(new_n257_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n441_), .A2(new_n442_), .A3(KEYINPUT87), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n448_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n673_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n452_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n693_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n469_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n692_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT110), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n470_), .A2(KEYINPUT110), .A3(new_n692_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n688_), .B(KEYINPUT109), .Z(new_n704_));
  OAI21_X1  g503(.A(new_n704_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n705_));
  AOI22_X1  g504(.A1(new_n702_), .A2(new_n703_), .B1(KEYINPUT43), .B2(new_n705_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n641_), .A2(new_n681_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n687_), .B1(new_n706_), .B2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n705_), .A2(KEYINPUT43), .ZN(new_n710_));
  AOI21_X1  g509(.A(KEYINPUT110), .B1(new_n470_), .B2(new_n692_), .ZN(new_n711_));
  AOI211_X1 g510(.A(new_n701_), .B(new_n691_), .C1(new_n453_), .C2(new_n469_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n710_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(KEYINPUT44), .A3(new_n707_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n709_), .A2(new_n635_), .A3(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT111), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n715_), .A2(new_n716_), .A3(G29gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n715_), .B2(G29gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n686_), .B1(new_n717_), .B2(new_n718_), .ZN(G1328gat));
  INV_X1    g518(.A(KEYINPUT46), .ZN(new_n720_));
  INV_X1    g519(.A(G36gat), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n713_), .A2(new_n707_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n648_), .B1(new_n722_), .B2(new_n687_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n721_), .B1(new_n723_), .B2(new_n714_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n684_), .A2(new_n721_), .A3(new_n649_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT45), .Z(new_n726_));
  OAI21_X1  g525(.A(new_n720_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n709_), .A2(new_n649_), .A3(new_n714_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(G36gat), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n725_), .B(KEYINPUT45), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n729_), .A2(KEYINPUT46), .A3(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n727_), .A2(new_n731_), .ZN(G1329gat));
  AOI21_X1  g531(.A(G43gat), .B1(new_n684_), .B2(new_n663_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT112), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n441_), .A2(new_n442_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n709_), .A2(new_n714_), .A3(G43gat), .A4(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n734_), .A2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT47), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT47), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n734_), .A2(new_n737_), .A3(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(G1330gat));
  AOI21_X1  g541(.A(G50gat), .B1(new_n684_), .B2(new_n673_), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n709_), .A2(G50gat), .A3(new_n673_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n744_), .B2(new_n714_), .ZN(G1331gat));
  NOR2_X1   g544(.A1(new_n471_), .A2(new_n638_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n631_), .A2(new_n512_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n747_), .A2(new_n538_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n746_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(G57gat), .B1(new_n750_), .B2(new_n257_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n631_), .A2(new_n600_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n512_), .B1(new_n752_), .B2(KEYINPUT113), .ZN(new_n753_));
  AOI211_X1 g552(.A(new_n753_), .B(new_n471_), .C1(KEYINPUT113), .C2(new_n752_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(new_n204_), .A3(new_n635_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n751_), .A2(new_n755_), .ZN(G1332gat));
  INV_X1    g555(.A(G64gat), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n757_), .B1(new_n749_), .B2(new_n649_), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT48), .Z(new_n759_));
  NAND2_X1  g558(.A1(new_n649_), .A2(new_n757_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT114), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n754_), .A2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n759_), .A2(new_n762_), .ZN(G1333gat));
  INV_X1    g562(.A(G71gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n764_), .B1(new_n749_), .B2(new_n663_), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT49), .Z(new_n766_));
  NAND3_X1  g565(.A1(new_n754_), .A2(new_n764_), .A3(new_n663_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(G1334gat));
  AOI21_X1  g567(.A(new_n528_), .B1(new_n749_), .B2(new_n673_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT50), .Z(new_n770_));
  NAND3_X1  g569(.A1(new_n754_), .A2(new_n528_), .A3(new_n673_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(G1335gat));
  NOR2_X1   g571(.A1(new_n747_), .A2(new_n681_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n713_), .A2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(G85gat), .B1(new_n774_), .B2(new_n257_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n471_), .A2(new_n683_), .A3(new_n747_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n776_), .A2(new_n206_), .A3(new_n635_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(G1336gat));
  OAI21_X1  g577(.A(G92gat), .B1(new_n774_), .B2(new_n648_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n776_), .A2(new_n548_), .A3(new_n649_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(G1337gat));
  OAI21_X1  g580(.A(G99gat), .B1(new_n774_), .B2(new_n454_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n776_), .A2(new_n736_), .A3(new_n569_), .A4(new_n570_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT115), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT51), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n782_), .A2(new_n783_), .A3(new_n785_), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n784_), .A2(KEYINPUT51), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n786_), .B(new_n787_), .ZN(G1338gat));
  NAND3_X1  g587(.A1(new_n776_), .A2(new_n555_), .A3(new_n673_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n713_), .A2(new_n673_), .A3(new_n773_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n790_), .A2(new_n791_), .A3(G106gat), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n790_), .B2(G106gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n789_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT53), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n796_), .B(new_n789_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(G1339gat));
  NAND2_X1  g597(.A1(new_n648_), .A2(new_n635_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n799_), .A2(new_n697_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n623_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n512_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n612_), .A2(KEYINPUT117), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT55), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n606_), .B1(new_n609_), .B2(new_n611_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(G230gat), .A3(G233gat), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT118), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n612_), .A2(KEYINPUT117), .A3(new_n810_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n806_), .A2(KEYINPUT118), .A3(G230gat), .A4(G233gat), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n805_), .A2(new_n809_), .A3(new_n811_), .A4(new_n812_), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n813_), .A2(KEYINPUT56), .A3(new_n621_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT56), .B1(new_n813_), .B2(new_n621_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n803_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT119), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n503_), .A2(new_n817_), .A3(new_n492_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n817_), .B1(new_n503_), .B2(new_n492_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n495_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n493_), .A2(new_n494_), .A3(new_n496_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n508_), .A3(new_n821_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n511_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n624_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n816_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n595_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(KEYINPUT120), .A3(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n595_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n829_), .B1(new_n816_), .B2(new_n824_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT120), .ZN(new_n831_));
  OAI21_X1  g630(.A(KEYINPUT57), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n823_), .A2(KEYINPUT121), .A3(new_n623_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT121), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n511_), .A2(new_n822_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(new_n802_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n833_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n815_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n813_), .A2(KEYINPUT56), .A3(new_n621_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n837_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n688_), .B1(new_n840_), .B2(KEYINPUT58), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n814_), .A2(new_n815_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n837_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n841_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n828_), .A2(new_n832_), .A3(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n538_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n600_), .A2(new_n630_), .A3(new_n848_), .A4(new_n512_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT116), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n600_), .A2(new_n630_), .A3(new_n512_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT54), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n849_), .A2(new_n850_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  AOI211_X1 g656(.A(KEYINPUT59), .B(new_n801_), .C1(new_n847_), .C2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n859_), .B1(new_n847_), .B2(new_n857_), .ZN(new_n860_));
  AOI211_X1 g659(.A(KEYINPUT122), .B(new_n856_), .C1(new_n846_), .C2(new_n538_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n800_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n858_), .B1(new_n862_), .B2(KEYINPUT59), .ZN(new_n863_));
  INV_X1    g662(.A(new_n512_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(G113gat), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n866_), .ZN(new_n867_));
  OAI22_X1  g666(.A1(new_n865_), .A2(new_n866_), .B1(new_n862_), .B2(new_n867_), .ZN(G1340gat));
  AOI21_X1  g667(.A(new_n831_), .B1(new_n825_), .B2(new_n595_), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n869_), .A2(new_n827_), .B1(new_n841_), .B2(new_n844_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n681_), .B1(new_n870_), .B2(new_n832_), .ZN(new_n871_));
  OAI21_X1  g670(.A(KEYINPUT122), .B1(new_n871_), .B2(new_n856_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n847_), .A2(new_n859_), .A3(new_n857_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT60), .ZN(new_n875_));
  INV_X1    g674(.A(G120gat), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n631_), .A2(new_n875_), .A3(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n874_), .A2(new_n800_), .A3(new_n878_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n863_), .A2(new_n631_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(new_n876_), .ZN(G1341gat));
  INV_X1    g680(.A(G127gat), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(new_n862_), .B2(new_n538_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(KEYINPUT123), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT123), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n885_), .B(new_n882_), .C1(new_n862_), .C2(new_n538_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n538_), .A2(new_n882_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(KEYINPUT124), .ZN(new_n888_));
  AOI22_X1  g687(.A1(new_n884_), .A2(new_n886_), .B1(new_n863_), .B2(new_n888_), .ZN(G1342gat));
  AND2_X1   g688(.A1(new_n863_), .A2(new_n689_), .ZN(new_n890_));
  INV_X1    g689(.A(G134gat), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n638_), .A2(new_n891_), .ZN(new_n892_));
  OAI22_X1  g691(.A1(new_n890_), .A2(new_n891_), .B1(new_n862_), .B2(new_n892_), .ZN(G1343gat));
  AOI21_X1  g692(.A(new_n696_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n799_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n512_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(new_n214_), .ZN(G1344gat));
  NOR2_X1   g697(.A1(new_n896_), .A2(new_n630_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n215_), .ZN(G1345gat));
  NOR2_X1   g699(.A1(new_n896_), .A2(new_n538_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT61), .B(G155gat), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n901_), .B(new_n903_), .ZN(G1346gat));
  INV_X1    g703(.A(new_n896_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n638_), .ZN(new_n906_));
  INV_X1    g705(.A(G162gat), .ZN(new_n907_));
  AND2_X1   g706(.A1(new_n704_), .A2(G162gat), .ZN(new_n908_));
  AOI22_X1  g707(.A1(new_n906_), .A2(new_n907_), .B1(new_n905_), .B2(new_n908_), .ZN(G1347gat));
  NOR2_X1   g708(.A1(new_n648_), .A2(new_n635_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n663_), .ZN(new_n911_));
  AOI211_X1 g710(.A(new_n673_), .B(new_n911_), .C1(new_n847_), .C2(new_n857_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n284_), .B1(new_n912_), .B2(new_n864_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n913_), .B(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT125), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n912_), .B(new_n916_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n864_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n915_), .B1(new_n917_), .B2(new_n918_), .ZN(G1348gat));
  XNOR2_X1  g718(.A(new_n912_), .B(KEYINPUT125), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n631_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n673_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n911_), .A2(new_n288_), .A3(new_n630_), .ZN(new_n923_));
  AOI22_X1  g722(.A1(new_n921_), .A2(new_n288_), .B1(new_n922_), .B2(new_n923_), .ZN(G1349gat));
  NOR2_X1   g723(.A1(new_n538_), .A2(new_n308_), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n922_), .A2(new_n663_), .A3(new_n681_), .A4(new_n910_), .ZN(new_n926_));
  AOI22_X1  g725(.A1(new_n920_), .A2(new_n925_), .B1(new_n926_), .B2(new_n273_), .ZN(G1350gat));
  OAI21_X1  g726(.A(G190gat), .B1(new_n917_), .B2(new_n688_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n920_), .A2(new_n309_), .A3(new_n638_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(G1351gat));
  OAI211_X1 g729(.A(new_n451_), .B(new_n910_), .C1(new_n860_), .C2(new_n861_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n864_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(G197gat), .ZN(G1352gat));
  AOI21_X1  g733(.A(new_n630_), .B1(KEYINPUT126), .B2(G204gat), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n932_), .A2(new_n935_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT126), .ZN(new_n937_));
  INV_X1    g736(.A(G204gat), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(new_n938_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n936_), .B(new_n939_), .ZN(G1353gat));
  NOR2_X1   g739(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n941_), .B1(new_n931_), .B2(new_n538_), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT127), .ZN(new_n943_));
  XOR2_X1   g742(.A(KEYINPUT63), .B(G211gat), .Z(new_n944_));
  NAND4_X1  g743(.A1(new_n894_), .A2(new_n681_), .A3(new_n910_), .A4(new_n944_), .ZN(new_n945_));
  AND3_X1   g744(.A1(new_n942_), .A2(new_n943_), .A3(new_n945_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n943_), .B1(new_n942_), .B2(new_n945_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n946_), .A2(new_n947_), .ZN(G1354gat));
  OAI21_X1  g747(.A(G218gat), .B1(new_n931_), .B2(new_n688_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n638_), .A2(new_n261_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n949_), .B1(new_n931_), .B2(new_n950_), .ZN(G1355gat));
endmodule


