//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 0 1 0 0 1 1 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 1 1 0 0 0 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n936_, new_n937_, new_n938_, new_n940_, new_n941_, new_n943_,
    new_n944_, new_n946_, new_n947_, new_n948_, new_n949_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n966_, new_n967_, new_n969_, new_n970_, new_n971_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n980_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n988_,
    new_n989_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XOR2_X1   g006(.A(new_n206_), .B(new_n207_), .Z(new_n208_));
  XNOR2_X1  g007(.A(G43gat), .B(G50gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G36gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G29gat), .ZN(new_n212_));
  INV_X1    g011(.A(G29gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(G36gat), .ZN(new_n214_));
  AND3_X1   g013(.A1(new_n212_), .A2(new_n214_), .A3(KEYINPUT71), .ZN(new_n215_));
  AOI21_X1  g014(.A(KEYINPUT71), .B1(new_n212_), .B2(new_n214_), .ZN(new_n216_));
  NOR3_X1   g015(.A1(new_n215_), .A2(new_n216_), .A3(KEYINPUT72), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT72), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT71), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n213_), .A2(G36gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n211_), .A2(G29gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n219_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n212_), .A2(new_n214_), .A3(KEYINPUT71), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n218_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n210_), .B1(new_n217_), .B2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT72), .B1(new_n215_), .B2(new_n216_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n222_), .A2(new_n218_), .A3(new_n223_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(new_n227_), .A3(new_n209_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n225_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT15), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n225_), .A2(KEYINPUT15), .A3(new_n228_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n208_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n228_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n209_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(new_n208_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G229gat), .A2(G233gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n233_), .A2(new_n239_), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n236_), .A2(new_n208_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(new_n237_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n238_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n240_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G113gat), .B(G141gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G169gat), .B(G197gat), .ZN(new_n247_));
  XOR2_X1   g046(.A(new_n246_), .B(new_n247_), .Z(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n245_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n240_), .A2(new_n244_), .A3(new_n248_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n252_), .B(KEYINPUT78), .Z(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT85), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT25), .ZN(new_n256_));
  INV_X1    g055(.A(G190gat), .ZN(new_n257_));
  OAI22_X1  g056(.A1(new_n256_), .A2(G183gat), .B1(new_n257_), .B2(KEYINPUT26), .ZN(new_n258_));
  INV_X1    g057(.A(G183gat), .ZN(new_n259_));
  NOR3_X1   g058(.A1(new_n259_), .A2(KEYINPUT79), .A3(KEYINPUT25), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n256_), .A2(G183gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n257_), .A2(KEYINPUT26), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT80), .ZN(new_n264_));
  AOI22_X1  g063(.A1(KEYINPUT79), .A2(new_n262_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n257_), .A2(KEYINPUT80), .A3(KEYINPUT26), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n261_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT23), .B1(new_n259_), .B2(new_n257_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n259_), .A2(KEYINPUT23), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT82), .B1(new_n269_), .B2(G190gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT23), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n271_), .A2(G183gat), .A3(G190gat), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT82), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n268_), .B1(new_n270_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(G169gat), .ZN(new_n276_));
  INV_X1    g075(.A(G176gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(new_n277_), .A3(KEYINPUT81), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT81), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n279_), .B1(G169gat), .B2(G176gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT24), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT24), .B1(new_n276_), .B2(new_n277_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n285_), .A2(new_n278_), .A3(new_n280_), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n267_), .A2(new_n275_), .A3(new_n283_), .A4(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(G169gat), .ZN(new_n289_));
  AND2_X1   g088(.A1(new_n268_), .A2(new_n272_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n289_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  AND2_X1   g091(.A1(new_n287_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT84), .B(G43gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G227gat), .A2(G233gat), .ZN(new_n296_));
  INV_X1    g095(.A(G15gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(G71gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(G99gat), .ZN(new_n300_));
  INV_X1    g099(.A(G71gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n298_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(G99gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n300_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT83), .B(KEYINPUT30), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n306_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n300_), .A2(new_n304_), .A3(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n295_), .A2(new_n310_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n295_), .A2(new_n310_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G127gat), .B(G134gat), .Z(new_n313_));
  XOR2_X1   g112(.A(G113gat), .B(G120gat), .Z(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT31), .ZN(new_n316_));
  OR4_X1    g115(.A1(new_n255_), .A2(new_n311_), .A3(new_n312_), .A4(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n255_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n295_), .A2(new_n310_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n295_), .A2(new_n310_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(KEYINPUT85), .A3(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n318_), .A2(new_n321_), .A3(new_n316_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n317_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT86), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n317_), .A2(new_n322_), .A3(KEYINPUT86), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G78gat), .B(G106gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G22gat), .B(G50gat), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n328_), .B(new_n329_), .Z(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G197gat), .B(G204gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G211gat), .B(G218gat), .ZN(new_n333_));
  OAI211_X1 g132(.A(KEYINPUT21), .B(new_n332_), .C1(new_n333_), .C2(KEYINPUT90), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT21), .ZN(new_n335_));
  INV_X1    g134(.A(G218gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(G211gat), .ZN(new_n337_));
  INV_X1    g136(.A(G211gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(G218gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT90), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n335_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  AND2_X1   g141(.A1(G197gat), .A2(G204gat), .ZN(new_n343_));
  NOR2_X1   g142(.A1(G197gat), .A2(G204gat), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n345_), .B1(new_n333_), .B2(KEYINPUT21), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n334_), .B1(new_n342_), .B2(new_n346_), .ZN(new_n347_));
  OR2_X1    g146(.A1(new_n347_), .A2(KEYINPUT91), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(KEYINPUT91), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(KEYINPUT87), .A2(G155gat), .A3(G162gat), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT87), .B1(G155gat), .B2(G162gat), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT1), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G155gat), .A2(G162gat), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT87), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT1), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n359_), .A2(new_n360_), .A3(new_n351_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n354_), .A2(new_n356_), .A3(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G141gat), .A2(G148gat), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(G141gat), .A2(G148gat), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT88), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT2), .B1(new_n364_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT2), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n363_), .A2(KEYINPUT88), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT3), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n365_), .A2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n368_), .A2(new_n370_), .A3(new_n372_), .A4(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n355_), .B1(new_n359_), .B2(new_n351_), .ZN(new_n375_));
  AOI22_X1  g174(.A1(new_n362_), .A2(new_n366_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT29), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  OAI211_X1 g177(.A(G228gat), .B(G233gat), .C1(new_n350_), .C2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n376_), .A2(new_n377_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT28), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT89), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n382_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n362_), .A2(new_n366_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n374_), .A2(new_n375_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(KEYINPUT89), .A3(KEYINPUT29), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G228gat), .A2(G233gat), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n383_), .A2(new_n387_), .A3(new_n347_), .A4(new_n388_), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n379_), .A2(new_n381_), .A3(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n381_), .B1(new_n379_), .B2(new_n389_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n331_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n379_), .A2(new_n389_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n381_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n379_), .A2(new_n381_), .A3(new_n389_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n395_), .A2(new_n396_), .A3(new_n330_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n392_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G1gat), .B(G29gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(G85gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT0), .B(G57gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G225gat), .A2(G233gat), .ZN(new_n405_));
  INV_X1    g204(.A(new_n315_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n386_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n376_), .A2(new_n315_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n408_), .A3(KEYINPUT4), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n315_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT4), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n405_), .B1(new_n409_), .B2(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n386_), .A2(new_n406_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n405_), .B1(new_n414_), .B2(new_n410_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n404_), .B1(new_n413_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT33), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT33), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n419_), .B(new_n404_), .C1(new_n413_), .C2(new_n416_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n409_), .A2(new_n405_), .A3(new_n412_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n414_), .A2(new_n410_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n405_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n404_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n418_), .A2(new_n420_), .B1(new_n421_), .B2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G226gat), .A2(G233gat), .ZN(new_n427_));
  XOR2_X1   g226(.A(new_n426_), .B(new_n427_), .Z(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(KEYINPUT93), .ZN(new_n429_));
  INV_X1    g228(.A(new_n347_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(new_n287_), .A3(new_n292_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n431_), .A2(KEYINPUT94), .A3(KEYINPUT20), .ZN(new_n432_));
  INV_X1    g231(.A(new_n268_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n269_), .A2(KEYINPUT82), .A3(G190gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n272_), .A2(new_n273_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n433_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n289_), .B1(new_n436_), .B2(new_n291_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT25), .B(G183gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT26), .B(G190gat), .ZN(new_n439_));
  AOI22_X1  g238(.A1(new_n438_), .A2(new_n439_), .B1(new_n268_), .B2(new_n272_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n284_), .A2(KEYINPUT95), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n441_), .A2(new_n278_), .A3(new_n280_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n284_), .A2(KEYINPUT95), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n283_), .B(new_n440_), .C1(new_n442_), .C2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n437_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(new_n347_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n432_), .A2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT94), .B1(new_n431_), .B2(KEYINPUT20), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n429_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT20), .B1(new_n293_), .B2(new_n430_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n428_), .B1(new_n445_), .B2(new_n347_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(G8gat), .B(G36gat), .Z(new_n454_));
  XNOR2_X1  g253(.A(G64gat), .B(G92gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n449_), .A2(new_n453_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n458_), .B1(new_n449_), .B2(new_n453_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT97), .ZN(new_n462_));
  NOR3_X1   g261(.A1(new_n460_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n449_), .A2(new_n453_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n458_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(KEYINPUT97), .B1(new_n466_), .B2(new_n459_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n425_), .B1(new_n463_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n428_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n445_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n469_), .B1(new_n450_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT98), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n431_), .A2(KEYINPUT20), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT94), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n429_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n476_), .A2(new_n446_), .A3(new_n432_), .A4(new_n477_), .ZN(new_n478_));
  OAI211_X1 g277(.A(KEYINPUT98), .B(new_n469_), .C1(new_n450_), .C2(new_n470_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n473_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n458_), .A2(KEYINPUT32), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT99), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n476_), .A2(new_n446_), .A3(new_n432_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n452_), .B1(new_n486_), .B2(new_n429_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(new_n481_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n413_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n489_), .A2(new_n403_), .A3(new_n415_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(new_n417_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n480_), .A2(KEYINPUT99), .A3(new_n482_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n485_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n399_), .B1(new_n468_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n480_), .A2(new_n465_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT27), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n497_), .B1(new_n487_), .B2(new_n458_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n497_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n491_), .B1(new_n392_), .B2(new_n397_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n327_), .B1(new_n495_), .B2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n398_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT100), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n491_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n323_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n398_), .A2(new_n499_), .A3(new_n500_), .A4(KEYINPUT100), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .A4(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n254_), .B1(new_n505_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT66), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT7), .ZN(new_n516_));
  INV_X1    g315(.A(G106gat), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n516_), .A2(new_n303_), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT6), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n519_), .B1(G99gat), .B2(G106gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G99gat), .A2(G106gat), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n521_), .A2(KEYINPUT6), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n515_), .B(new_n518_), .C1(new_n520_), .C2(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(G85gat), .B(G92gat), .Z(new_n524_));
  AOI21_X1  g323(.A(new_n514_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT8), .ZN(new_n526_));
  NAND3_X1  g325(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT65), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(G85gat), .ZN(new_n530_));
  INV_X1    g329(.A(G92gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  AND2_X1   g331(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n533_));
  NOR2_X1   g332(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n534_));
  OAI22_X1  g333(.A1(new_n533_), .A2(new_n534_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n529_), .A2(new_n532_), .A3(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(KEYINPUT10), .B(G99gat), .Z(new_n537_));
  NAND2_X1  g336(.A1(new_n521_), .A2(KEYINPUT6), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n519_), .A2(G99gat), .A3(G106gat), .ZN(new_n539_));
  AOI22_X1  g338(.A1(new_n537_), .A2(new_n517_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n525_), .A2(new_n526_), .B1(new_n536_), .B2(new_n540_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n538_), .A2(new_n539_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n518_), .A2(new_n515_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n524_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT66), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n523_), .A2(new_n514_), .A3(new_n524_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n545_), .A2(KEYINPUT8), .A3(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G57gat), .B(G64gat), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n548_), .A2(KEYINPUT11), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(KEYINPUT11), .ZN(new_n550_));
  XOR2_X1   g349(.A(G71gat), .B(G78gat), .Z(new_n551_));
  NAND3_X1  g350(.A1(new_n549_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n550_), .A2(new_n551_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n541_), .A2(new_n547_), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n554_), .B1(new_n541_), .B2(new_n547_), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT12), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G230gat), .A2(G233gat), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT12), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n523_), .A2(new_n514_), .A3(new_n524_), .ZN(new_n560_));
  NOR3_X1   g359(.A1(new_n560_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n544_), .A2(KEYINPUT66), .A3(new_n526_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n536_), .A2(new_n540_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n559_), .B1(new_n565_), .B2(new_n554_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n557_), .A2(new_n558_), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT67), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n554_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n570_), .B1(new_n561_), .B2(new_n564_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n541_), .A2(new_n547_), .A3(new_n554_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n558_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n557_), .A2(new_n566_), .A3(KEYINPUT67), .A4(new_n558_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n569_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(G176gat), .B(G204gat), .Z(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT69), .ZN(new_n579_));
  XOR2_X1   g378(.A(G120gat), .B(G148gat), .Z(new_n580_));
  XOR2_X1   g379(.A(new_n579_), .B(new_n580_), .Z(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n577_), .A2(new_n584_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n569_), .A2(new_n575_), .A3(new_n576_), .A4(new_n583_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(KEYINPUT70), .A3(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT70), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n577_), .A2(new_n588_), .A3(new_n584_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n587_), .A2(KEYINPUT13), .A3(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(KEYINPUT13), .B1(new_n587_), .B2(new_n589_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(G190gat), .B(G218gat), .Z(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT73), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G134gat), .B(G162gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT36), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G232gat), .A2(G233gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT34), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT35), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  AOI22_X1  g401(.A1(new_n231_), .A2(new_n232_), .B1(new_n547_), .B2(new_n541_), .ZN(new_n603_));
  OAI21_X1  g402(.A(KEYINPUT74), .B1(new_n599_), .B2(KEYINPUT35), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n541_), .A2(new_n547_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n605_), .B1(new_n606_), .B2(new_n229_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n602_), .B1(new_n603_), .B2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n596_), .A2(KEYINPUT36), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n604_), .B1(new_n565_), .B2(new_n236_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n602_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n234_), .A2(new_n235_), .A3(new_n230_), .ZN(new_n612_));
  AOI21_X1  g411(.A(KEYINPUT15), .B1(new_n225_), .B2(new_n228_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n606_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n610_), .A2(new_n611_), .A3(new_n614_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n608_), .A2(new_n609_), .A3(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n609_), .B1(new_n608_), .B2(new_n615_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n597_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT76), .ZN(new_n619_));
  OAI21_X1  g418(.A(KEYINPUT37), .B1(new_n616_), .B2(KEYINPUT75), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT76), .ZN(new_n622_));
  OAI211_X1 g421(.A(new_n622_), .B(new_n597_), .C1(new_n616_), .C2(new_n617_), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n619_), .A2(new_n621_), .A3(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n621_), .B1(new_n619_), .B2(new_n623_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n208_), .B(new_n554_), .Z(new_n627_));
  NAND2_X1  g426(.A1(G231gat), .A2(G233gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT17), .ZN(new_n630_));
  XOR2_X1   g429(.A(G127gat), .B(G155gat), .Z(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT16), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G183gat), .B(G211gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  OR3_X1    g433(.A1(new_n629_), .A2(new_n630_), .A3(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(KEYINPUT17), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n629_), .A2(new_n636_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT77), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n592_), .A2(new_n626_), .A3(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n513_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n642_), .A2(new_n203_), .A3(new_n491_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n644_), .A2(KEYINPUT38), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT101), .Z(new_n646_));
  AOI21_X1  g445(.A(new_n618_), .B1(new_n505_), .B2(new_n512_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n592_), .ZN(new_n648_));
  AND4_X1   g447(.A1(new_n252_), .A2(new_n647_), .A3(new_n638_), .A4(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n203_), .B1(new_n649_), .B2(new_n491_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n650_), .B1(new_n644_), .B2(KEYINPUT38), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n646_), .A2(new_n651_), .ZN(G1324gat));
  AOI21_X1  g451(.A(new_n204_), .B1(new_n649_), .B2(new_n501_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT39), .Z(new_n654_));
  NAND3_X1  g453(.A1(new_n642_), .A2(new_n204_), .A3(new_n501_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n654_), .A2(new_n655_), .A3(new_n657_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1325gat));
  AND3_X1   g460(.A1(new_n317_), .A2(new_n322_), .A3(KEYINPUT86), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT86), .B1(new_n317_), .B2(new_n322_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n297_), .B1(new_n649_), .B2(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT41), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n642_), .A2(new_n297_), .A3(new_n664_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1326gat));
  INV_X1    g467(.A(G22gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n669_), .B1(new_n649_), .B2(new_n399_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT42), .Z(new_n671_));
  NAND3_X1  g470(.A1(new_n642_), .A2(new_n669_), .A3(new_n399_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1327gat));
  INV_X1    g472(.A(new_n639_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n618_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n513_), .A2(new_n648_), .A3(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n513_), .A2(KEYINPUT106), .A3(new_n648_), .A4(new_n676_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(G29gat), .B1(new_n681_), .B2(new_n491_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n480_), .A2(KEYINPUT99), .A3(new_n482_), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT99), .B1(new_n480_), .B2(new_n482_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n488_), .A2(new_n491_), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n683_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n418_), .A2(new_n420_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n424_), .A2(new_n421_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n462_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n466_), .A2(KEYINPUT97), .A3(new_n459_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n689_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n398_), .B1(new_n686_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n504_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n664_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n512_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT103), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n624_), .A2(new_n625_), .A3(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n619_), .A2(new_n623_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(new_n620_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n619_), .A2(new_n623_), .A3(new_n621_), .ZN(new_n701_));
  AOI21_X1  g500(.A(KEYINPUT103), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  OAI22_X1  g501(.A1(new_n695_), .A2(new_n696_), .B1(new_n698_), .B2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT43), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n505_), .A2(new_n512_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n705_), .A2(new_n706_), .A3(new_n626_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n704_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT105), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n648_), .A2(new_n252_), .A3(new_n639_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n708_), .A2(new_n709_), .A3(KEYINPUT44), .A4(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n697_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n700_), .A2(new_n701_), .A3(KEYINPUT103), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n706_), .B1(new_n705_), .B2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n626_), .A2(new_n706_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n717_), .B1(new_n505_), .B2(new_n512_), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n711_), .B(KEYINPUT44), .C1(new_n716_), .C2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT105), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n711_), .B1(new_n716_), .B2(new_n718_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n722_));
  AOI22_X1  g521(.A1(new_n712_), .A2(new_n720_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n509_), .A2(new_n213_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n682_), .B1(new_n723_), .B2(new_n724_), .ZN(G1328gat));
  NAND2_X1  g524(.A1(new_n712_), .A2(new_n720_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n501_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n727_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(G36gat), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT107), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT46), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n679_), .A2(new_n211_), .A3(new_n501_), .A4(new_n680_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT45), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n730_), .A2(new_n731_), .A3(new_n732_), .A4(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n731_), .A2(new_n732_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n211_), .B1(new_n726_), .B2(new_n728_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n733_), .B(new_n739_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n736_), .B(new_n737_), .C1(new_n738_), .C2(new_n740_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n735_), .A2(new_n741_), .ZN(G1329gat));
  AND3_X1   g541(.A1(new_n723_), .A2(G43gat), .A3(new_n510_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n679_), .A2(new_n664_), .A3(new_n680_), .ZN(new_n744_));
  INV_X1    g543(.A(G43gat), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT108), .ZN(new_n747_));
  OAI21_X1  g546(.A(KEYINPUT47), .B1(new_n743_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n746_), .B(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT47), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n723_), .A2(G43gat), .A3(new_n510_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n750_), .A2(new_n751_), .A3(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n748_), .A2(new_n753_), .ZN(G1330gat));
  INV_X1    g553(.A(G50gat), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n681_), .A2(new_n755_), .A3(new_n399_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n723_), .A2(new_n399_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n757_), .A2(KEYINPUT109), .A3(G50gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT109), .B1(new_n757_), .B2(G50gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n756_), .B1(new_n758_), .B2(new_n759_), .ZN(G1331gat));
  INV_X1    g559(.A(new_n252_), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n705_), .A2(new_n761_), .A3(new_n592_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n626_), .A2(new_n639_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(G57gat), .B1(new_n765_), .B2(new_n491_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT110), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n647_), .A2(new_n254_), .A3(new_n674_), .A4(new_n592_), .ZN(new_n768_));
  XOR2_X1   g567(.A(KEYINPUT111), .B(G57gat), .Z(new_n769_));
  NOR3_X1   g568(.A1(new_n768_), .A2(new_n509_), .A3(new_n769_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n767_), .A2(new_n770_), .ZN(G1332gat));
  OAI21_X1  g570(.A(G64gat), .B1(new_n768_), .B2(new_n727_), .ZN(new_n772_));
  XOR2_X1   g571(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n773_));
  XNOR2_X1  g572(.A(new_n772_), .B(new_n773_), .ZN(new_n774_));
  OR2_X1    g573(.A1(new_n727_), .A2(G64gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n764_), .B2(new_n775_), .ZN(G1333gat));
  OAI21_X1  g575(.A(G71gat), .B1(new_n768_), .B2(new_n327_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT49), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n765_), .A2(new_n301_), .A3(new_n664_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(G1334gat));
  OAI21_X1  g579(.A(G78gat), .B1(new_n768_), .B2(new_n398_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT50), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n398_), .A2(G78gat), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT113), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n782_), .B1(new_n764_), .B2(new_n784_), .ZN(G1335gat));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n716_), .A2(new_n718_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n648_), .A2(new_n252_), .A3(new_n674_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n786_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n708_), .A2(KEYINPUT114), .A3(new_n788_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(G85gat), .B1(new_n792_), .B2(new_n509_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n762_), .A2(new_n676_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n795_), .A2(new_n530_), .A3(new_n491_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n793_), .A2(new_n796_), .ZN(G1336gat));
  OAI21_X1  g596(.A(G92gat), .B1(new_n792_), .B2(new_n727_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n795_), .A2(new_n531_), .A3(new_n501_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(G1337gat));
  NAND3_X1  g599(.A1(new_n795_), .A2(new_n510_), .A3(new_n537_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n327_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(new_n303_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g603(.A1(new_n795_), .A2(new_n517_), .A3(new_n399_), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n399_), .B(new_n788_), .C1(new_n716_), .C2(new_n718_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT115), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n806_), .A2(new_n807_), .A3(G106gat), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n807_), .B1(new_n806_), .B2(G106gat), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n809_), .A2(new_n810_), .A3(KEYINPUT52), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n806_), .A2(G106gat), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT115), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n812_), .B1(new_n814_), .B2(new_n808_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n805_), .B1(new_n811_), .B2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT53), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n818_), .B(new_n805_), .C1(new_n811_), .C2(new_n815_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(G1339gat));
  INV_X1    g619(.A(KEYINPUT122), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n640_), .A2(new_n254_), .ZN(new_n822_));
  XOR2_X1   g621(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n640_), .B(new_n254_), .C1(KEYINPUT116), .C2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n252_), .A2(new_n586_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  XOR2_X1   g629(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n831_));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n569_), .A2(new_n832_), .A3(new_n576_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n559_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT12), .B1(new_n606_), .B2(new_n570_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n574_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  OAI211_X1 g637(.A(KEYINPUT117), .B(new_n574_), .C1(new_n834_), .C2(new_n835_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NOR4_X1   g639(.A1(new_n834_), .A2(new_n835_), .A3(new_n832_), .A4(new_n574_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n833_), .A2(new_n840_), .A3(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n831_), .B1(new_n843_), .B2(new_n584_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT56), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n841_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n846_));
  AOI211_X1 g645(.A(new_n845_), .B(new_n583_), .C1(new_n846_), .C2(new_n833_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n830_), .B1(new_n844_), .B2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n248_), .B1(new_n242_), .B2(new_n238_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n237_), .A2(new_n243_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n233_), .B2(new_n850_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n851_), .A2(new_n251_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n587_), .A2(new_n589_), .A3(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n618_), .B1(new_n848_), .B2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(KEYINPUT57), .B1(new_n854_), .B2(KEYINPUT119), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n843_), .A2(new_n584_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n831_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n843_), .A2(KEYINPUT56), .A3(new_n584_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n829_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n853_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n675_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n855_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n618_), .A2(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n867_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n848_), .A2(new_n853_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n871_), .A2(KEYINPUT120), .A3(new_n867_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n872_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n852_), .A2(new_n586_), .ZN(new_n874_));
  AOI21_X1  g673(.A(KEYINPUT56), .B1(new_n843_), .B2(new_n584_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(new_n847_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT58), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  OAI211_X1 g677(.A(KEYINPUT58), .B(new_n874_), .C1(new_n875_), .C2(new_n847_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n878_), .A2(new_n626_), .A3(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n865_), .A2(new_n873_), .A3(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n638_), .B1(new_n881_), .B2(KEYINPUT121), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT121), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n865_), .A2(new_n873_), .A3(new_n883_), .A4(new_n880_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n828_), .B1(new_n882_), .B2(new_n884_), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n508_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n491_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n821_), .B1(new_n885_), .B2(new_n887_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n675_), .B(KEYINPUT119), .C1(new_n860_), .C2(new_n861_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n866_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n854_), .A2(KEYINPUT119), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(KEYINPUT120), .B1(new_n871_), .B2(new_n867_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n867_), .ZN(new_n894_));
  AOI211_X1 g693(.A(new_n869_), .B(new_n894_), .C1(new_n848_), .C2(new_n853_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n880_), .B1(new_n893_), .B2(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(KEYINPUT121), .B1(new_n892_), .B2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n638_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n897_), .A2(new_n898_), .A3(new_n884_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n827_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n887_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n900_), .A2(KEYINPUT122), .A3(new_n901_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n888_), .A2(new_n252_), .A3(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(G113gat), .ZN(new_n904_));
  OR2_X1    g703(.A1(new_n887_), .A2(KEYINPUT123), .ZN(new_n905_));
  AOI21_X1  g704(.A(KEYINPUT59), .B1(new_n887_), .B2(KEYINPUT123), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n881_), .A2(new_n639_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(new_n827_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n900_), .A2(new_n901_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(new_n910_), .B2(KEYINPUT59), .ZN(new_n911_));
  XNOR2_X1  g710(.A(KEYINPUT124), .B(G113gat), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n253_), .A2(new_n912_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(KEYINPUT125), .ZN(new_n914_));
  AOI22_X1  g713(.A1(new_n903_), .A2(new_n904_), .B1(new_n911_), .B2(new_n914_), .ZN(G1340gat));
  INV_X1    g714(.A(new_n909_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n887_), .B1(new_n899_), .B2(new_n827_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT59), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n916_), .B1(new_n917_), .B2(new_n918_), .ZN(new_n919_));
  OAI21_X1  g718(.A(G120gat), .B1(new_n919_), .B2(new_n648_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT60), .ZN(new_n921_));
  AOI21_X1  g720(.A(G120gat), .B1(new_n592_), .B2(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n922_), .B1(new_n921_), .B2(G120gat), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n888_), .A2(new_n902_), .A3(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n920_), .A2(new_n924_), .ZN(G1341gat));
  INV_X1    g724(.A(G127gat), .ZN(new_n926_));
  NAND4_X1  g725(.A1(new_n888_), .A2(new_n926_), .A3(new_n674_), .A4(new_n902_), .ZN(new_n927_));
  OAI211_X1 g726(.A(new_n638_), .B(new_n916_), .C1(new_n917_), .C2(new_n918_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n927_), .B1(new_n929_), .B2(new_n926_), .ZN(G1342gat));
  INV_X1    g729(.A(G134gat), .ZN(new_n931_));
  NAND4_X1  g730(.A1(new_n888_), .A2(new_n931_), .A3(new_n618_), .A4(new_n902_), .ZN(new_n932_));
  OAI211_X1 g731(.A(new_n626_), .B(new_n916_), .C1(new_n917_), .C2(new_n918_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n933_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n932_), .B1(new_n934_), .B2(new_n931_), .ZN(G1343gat));
  NOR4_X1   g734(.A1(new_n664_), .A2(new_n509_), .A3(new_n398_), .A4(new_n501_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n900_), .A2(new_n252_), .A3(new_n936_), .ZN(new_n937_));
  XOR2_X1   g736(.A(KEYINPUT126), .B(G141gat), .Z(new_n938_));
  XNOR2_X1  g737(.A(new_n937_), .B(new_n938_), .ZN(G1344gat));
  NAND3_X1  g738(.A1(new_n900_), .A2(new_n592_), .A3(new_n936_), .ZN(new_n940_));
  XOR2_X1   g739(.A(KEYINPUT127), .B(G148gat), .Z(new_n941_));
  XNOR2_X1  g740(.A(new_n940_), .B(new_n941_), .ZN(G1345gat));
  NAND3_X1  g741(.A1(new_n900_), .A2(new_n674_), .A3(new_n936_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(KEYINPUT61), .B(G155gat), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n943_), .B(new_n944_), .ZN(G1346gat));
  AND2_X1   g744(.A1(new_n900_), .A2(new_n936_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(new_n618_), .ZN(new_n947_));
  INV_X1    g746(.A(G162gat), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n948_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n949_));
  AOI22_X1  g748(.A1(new_n947_), .A2(new_n948_), .B1(new_n946_), .B2(new_n949_), .ZN(G1347gat));
  NAND2_X1  g749(.A1(new_n908_), .A2(new_n827_), .ZN(new_n951_));
  NOR3_X1   g750(.A1(new_n327_), .A2(new_n491_), .A3(new_n727_), .ZN(new_n952_));
  INV_X1    g751(.A(new_n952_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n953_), .A2(new_n399_), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n951_), .A2(new_n252_), .A3(new_n954_), .ZN(new_n955_));
  OAI21_X1  g754(.A(KEYINPUT62), .B1(new_n955_), .B2(KEYINPUT22), .ZN(new_n956_));
  OAI21_X1  g755(.A(G169gat), .B1(new_n955_), .B2(KEYINPUT62), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n956_), .A2(new_n957_), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n958_), .B1(new_n276_), .B2(new_n956_), .ZN(G1348gat));
  NAND2_X1  g758(.A1(new_n951_), .A2(new_n954_), .ZN(new_n960_));
  INV_X1    g759(.A(new_n960_), .ZN(new_n961_));
  AOI21_X1  g760(.A(G176gat), .B1(new_n961_), .B2(new_n592_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n885_), .A2(new_n399_), .ZN(new_n963_));
  NOR3_X1   g762(.A1(new_n953_), .A2(new_n648_), .A3(new_n277_), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n962_), .B1(new_n963_), .B2(new_n964_), .ZN(G1349gat));
  NOR3_X1   g764(.A1(new_n960_), .A2(new_n438_), .A3(new_n898_), .ZN(new_n966_));
  NAND3_X1  g765(.A1(new_n963_), .A2(new_n674_), .A3(new_n952_), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n966_), .B1(new_n967_), .B2(new_n259_), .ZN(G1350gat));
  INV_X1    g767(.A(new_n626_), .ZN(new_n969_));
  OAI21_X1  g768(.A(G190gat), .B1(new_n960_), .B2(new_n969_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n618_), .A2(new_n439_), .ZN(new_n971_));
  OAI21_X1  g770(.A(new_n970_), .B1(new_n960_), .B2(new_n971_), .ZN(G1351gat));
  NOR3_X1   g771(.A1(new_n664_), .A2(new_n503_), .A3(new_n727_), .ZN(new_n973_));
  AND2_X1   g772(.A1(new_n900_), .A2(new_n973_), .ZN(new_n974_));
  AOI21_X1  g773(.A(G197gat), .B1(new_n974_), .B2(new_n252_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n900_), .A2(new_n973_), .ZN(new_n976_));
  INV_X1    g775(.A(G197gat), .ZN(new_n977_));
  NOR3_X1   g776(.A1(new_n976_), .A2(new_n977_), .A3(new_n761_), .ZN(new_n978_));
  NOR2_X1   g777(.A1(new_n975_), .A2(new_n978_), .ZN(G1352gat));
  NAND3_X1  g778(.A1(new_n900_), .A2(new_n592_), .A3(new_n973_), .ZN(new_n980_));
  XNOR2_X1  g779(.A(new_n980_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g780(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n982_));
  AND2_X1   g781(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n983_));
  NOR4_X1   g782(.A1(new_n976_), .A2(new_n898_), .A3(new_n982_), .A4(new_n983_), .ZN(new_n984_));
  INV_X1    g783(.A(new_n982_), .ZN(new_n985_));
  AOI21_X1  g784(.A(new_n985_), .B1(new_n974_), .B2(new_n638_), .ZN(new_n986_));
  NOR2_X1   g785(.A1(new_n984_), .A2(new_n986_), .ZN(G1354gat));
  NAND3_X1  g786(.A1(new_n974_), .A2(new_n336_), .A3(new_n618_), .ZN(new_n988_));
  OAI21_X1  g787(.A(G218gat), .B1(new_n976_), .B2(new_n969_), .ZN(new_n989_));
  NAND2_X1  g788(.A1(new_n988_), .A2(new_n989_), .ZN(G1355gat));
endmodule


