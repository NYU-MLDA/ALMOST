//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 0 1 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 1 0 1 1 1 0 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 1 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n631_, new_n632_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n658_, new_n659_, new_n660_, new_n661_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n770_, new_n771_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n807_, new_n808_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n827_, new_n828_, new_n829_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G8gat), .B(G36gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n206_));
  XOR2_X1   g005(.A(new_n205_), .B(new_n206_), .Z(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT26), .B(G190gat), .ZN(new_n208_));
  INV_X1    g007(.A(G183gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT76), .B1(new_n209_), .B2(KEYINPUT25), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT25), .B(G183gat), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n208_), .B(new_n210_), .C1(new_n211_), .C2(KEYINPUT76), .ZN(new_n212_));
  XOR2_X1   g011(.A(G169gat), .B(G176gat), .Z(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT24), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n215_), .A2(KEYINPUT77), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT23), .ZN(new_n218_));
  OR3_X1    g017(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n215_), .A2(KEYINPUT77), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n216_), .A2(new_n218_), .A3(new_n219_), .A4(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n218_), .B1(G183gat), .B2(G190gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n223_));
  INV_X1    g022(.A(G169gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n223_), .B(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n222_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n221_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G211gat), .B(G218gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT87), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G197gat), .B(G204gat), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT21), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n230_), .A2(new_n233_), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n231_), .A2(new_n232_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n230_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n228_), .A2(new_n238_), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n225_), .B(KEYINPUT90), .Z(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(new_n222_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n242_));
  OR3_X1    g041(.A1(new_n242_), .A2(G169gat), .A3(G176gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n213_), .A2(new_n242_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n211_), .A2(new_n208_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n218_), .A4(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n241_), .A2(new_n237_), .A3(new_n246_), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n239_), .A2(KEYINPUT20), .A3(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G226gat), .A2(G233gat), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n249_), .B(KEYINPUT88), .Z(new_n250_));
  XOR2_X1   g049(.A(new_n250_), .B(KEYINPUT19), .Z(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n248_), .A2(new_n252_), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n221_), .A2(new_n227_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(new_n237_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n241_), .A2(new_n246_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(new_n238_), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n255_), .A2(KEYINPUT20), .A3(new_n252_), .A4(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n207_), .B1(new_n253_), .B2(new_n259_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n255_), .A2(KEYINPUT20), .A3(new_n251_), .A4(new_n257_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n261_), .B1(new_n248_), .B2(new_n251_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n207_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n260_), .A2(new_n264_), .A3(KEYINPUT27), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT95), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n258_), .B(new_n263_), .C1(new_n248_), .C2(new_n252_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n260_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT27), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G22gat), .B(G50gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT84), .ZN(new_n272_));
  INV_X1    g071(.A(G233gat), .ZN(new_n273_));
  OR2_X1    g072(.A1(KEYINPUT85), .A2(G228gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(KEYINPUT85), .A2(G228gat), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n273_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(new_n272_), .B(new_n276_), .Z(new_n277_));
  NAND2_X1  g076(.A1(G141gat), .A2(G148gat), .ZN(new_n278_));
  INV_X1    g077(.A(G141gat), .ZN(new_n279_));
  INV_X1    g078(.A(G148gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(G155gat), .A2(G162gat), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT82), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n284_), .B1(KEYINPUT1), .B2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(KEYINPUT1), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT83), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n278_), .B(new_n281_), .C1(new_n286_), .C2(new_n289_), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n281_), .A2(KEYINPUT3), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT2), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n278_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n281_), .A2(KEYINPUT3), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n291_), .A2(new_n293_), .A3(new_n294_), .A4(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n296_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n290_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT29), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n238_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n298_), .A2(KEYINPUT29), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NOR3_X1   g101(.A1(new_n238_), .A2(KEYINPUT29), .A3(new_n298_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n277_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n303_), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n298_), .A2(KEYINPUT29), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(new_n299_), .A3(new_n238_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n277_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n305_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n304_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G78gat), .B(G106gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n310_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n304_), .A2(new_n313_), .A3(new_n309_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT95), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n260_), .A2(new_n264_), .A3(new_n318_), .A4(KEYINPUT27), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n266_), .A2(new_n270_), .A3(new_n317_), .A4(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT96), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G127gat), .B(G134gat), .ZN(new_n323_));
  INV_X1    g122(.A(G113gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(G120gat), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(new_n298_), .B2(KEYINPUT92), .ZN(new_n327_));
  INV_X1    g126(.A(G120gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n325_), .B(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT92), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n329_), .A2(new_n330_), .A3(new_n290_), .A4(new_n297_), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n327_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G225gat), .A2(G233gat), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n327_), .A2(new_n331_), .A3(KEYINPUT4), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT4), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n298_), .A2(new_n326_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(new_n334_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G1gat), .B(G29gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(G85gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT0), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n344_), .B(G57gat), .Z(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n336_), .A2(new_n341_), .A3(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n333_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n345_), .B1(new_n335_), .B2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n347_), .A2(new_n349_), .A3(KEYINPUT94), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT94), .B1(new_n347_), .B2(new_n349_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(G71gat), .B(G99gat), .Z(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT30), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n228_), .B(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT78), .B(G43gat), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT79), .B(G15gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G227gat), .A2(G233gat), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n360_), .B(new_n361_), .Z(new_n362_));
  NOR2_X1   g161(.A1(new_n254_), .A2(new_n355_), .ZN(new_n363_));
  AND3_X1   g162(.A1(new_n221_), .A2(new_n227_), .A3(new_n355_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n357_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n359_), .A2(new_n362_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n362_), .B1(new_n359_), .B2(new_n365_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n326_), .B(KEYINPUT31), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT81), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  OAI22_X1  g170(.A1(new_n367_), .A2(new_n368_), .B1(KEYINPUT80), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n368_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n369_), .B1(KEYINPUT80), .B2(new_n370_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(new_n366_), .A3(new_n374_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n353_), .A2(new_n372_), .A3(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n321_), .A2(new_n322_), .A3(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n353_), .A2(new_n372_), .A3(new_n375_), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT96), .B1(new_n320_), .B2(new_n378_), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n351_), .A2(new_n352_), .A3(new_n317_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n380_), .A2(new_n270_), .A3(new_n266_), .A4(new_n319_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n347_), .A2(new_n349_), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n207_), .A2(KEYINPUT32), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n262_), .A2(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n253_), .A2(new_n259_), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n382_), .B(new_n384_), .C1(new_n385_), .C2(new_n383_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT33), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n349_), .A2(new_n387_), .ZN(new_n388_));
  OAI211_X1 g187(.A(KEYINPUT33), .B(new_n345_), .C1(new_n335_), .C2(new_n348_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n260_), .A2(new_n388_), .A3(new_n267_), .A4(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n332_), .A2(new_n334_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n337_), .A2(new_n333_), .A3(new_n339_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n392_), .A3(new_n346_), .ZN(new_n393_));
  XOR2_X1   g192(.A(new_n393_), .B(KEYINPUT93), .Z(new_n394_));
  OAI21_X1  g193(.A(new_n386_), .B1(new_n390_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n317_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n381_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n372_), .A2(new_n375_), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n377_), .A2(new_n379_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  XOR2_X1   g198(.A(G85gat), .B(G92gat), .Z(new_n400_));
  XOR2_X1   g199(.A(KEYINPUT10), .B(G99gat), .Z(new_n401_));
  INV_X1    g200(.A(G106gat), .ZN(new_n402_));
  AOI22_X1  g201(.A1(KEYINPUT9), .A2(new_n400_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT9), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n404_), .A2(G85gat), .A3(G92gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G99gat), .A2(G106gat), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT6), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT64), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT64), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT6), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n406_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n408_), .A2(new_n410_), .A3(new_n406_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n403_), .B(new_n405_), .C1(new_n411_), .C2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT65), .ZN(new_n414_));
  OAI22_X1  g213(.A1(new_n414_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n414_), .B1(KEYINPUT66), .B2(KEYINPUT7), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  OAI221_X1 g216(.A(new_n414_), .B1(KEYINPUT66), .B2(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n417_), .B(new_n418_), .C1(new_n412_), .C2(new_n411_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT8), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n419_), .A2(new_n420_), .A3(new_n400_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n420_), .B1(new_n419_), .B2(new_n400_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n413_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G57gat), .B(G64gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT11), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G71gat), .B(G78gat), .ZN(new_n426_));
  OR2_X1    g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n424_), .A2(KEYINPUT11), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n425_), .A2(new_n426_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n423_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n430_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n432_), .B(new_n413_), .C1(new_n421_), .C2(new_n422_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(KEYINPUT12), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT12), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n423_), .A2(new_n435_), .A3(new_n430_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(G230gat), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n438_), .A2(new_n273_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  AOI211_X1 g239(.A(new_n438_), .B(new_n273_), .C1(new_n431_), .C2(new_n433_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(G148gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G176gat), .B(G204gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT68), .B(G120gat), .ZN(new_n447_));
  XOR2_X1   g246(.A(new_n446_), .B(new_n447_), .Z(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n442_), .A2(new_n449_), .ZN(new_n450_));
  NOR3_X1   g249(.A1(new_n440_), .A2(new_n441_), .A3(new_n448_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  OR2_X1    g251(.A1(new_n452_), .A2(KEYINPUT13), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(KEYINPUT13), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G29gat), .B(G36gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(G43gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(G50gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G1gat), .B(G8gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT73), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G15gat), .B(G22gat), .ZN(new_n461_));
  INV_X1    g260(.A(G8gat), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n460_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n460_), .A2(new_n464_), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n458_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n458_), .B(KEYINPUT15), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n465_), .A2(new_n466_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n467_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G229gat), .A2(G233gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(new_n469_), .B(new_n458_), .Z(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(G229gat), .A3(G233gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G113gat), .B(G141gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(new_n224_), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n477_), .B(G197gat), .Z(new_n478_));
  NAND2_X1  g277(.A1(new_n475_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n478_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n472_), .A2(new_n474_), .A3(new_n480_), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n455_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n399_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n423_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n458_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n468_), .A2(new_n423_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G232gat), .A2(G233gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT34), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n490_), .A2(KEYINPUT35), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT70), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n487_), .A2(new_n488_), .A3(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n490_), .A2(KEYINPUT35), .ZN(new_n494_));
  XOR2_X1   g293(.A(new_n494_), .B(KEYINPUT69), .Z(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n493_), .B(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT72), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G190gat), .B(G218gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT71), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(G134gat), .ZN(new_n501_));
  INV_X1    g300(.A(G162gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT36), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n503_), .A2(new_n504_), .ZN(new_n506_));
  NOR4_X1   g305(.A1(new_n497_), .A2(new_n498_), .A3(new_n505_), .A4(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT72), .B1(new_n497_), .B2(new_n505_), .ZN(new_n508_));
  OR3_X1    g307(.A1(new_n497_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n507_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G127gat), .B(G155gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT16), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(new_n209_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(G211gat), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT75), .B1(new_n516_), .B2(KEYINPUT17), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G231gat), .A2(G233gat), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n518_), .B(KEYINPUT74), .Z(new_n519_));
  XNOR2_X1  g318(.A(new_n430_), .B(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n520_), .B(new_n469_), .Z(new_n521_));
  XNOR2_X1  g320(.A(new_n517_), .B(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n522_), .B1(KEYINPUT17), .B2(new_n516_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n511_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n485_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT98), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT98), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n485_), .A2(new_n528_), .A3(new_n525_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n353_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n202_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT99), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n497_), .A2(new_n505_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n509_), .A2(KEYINPUT37), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT37), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n536_), .B1(new_n510_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NOR4_X1   g338(.A1(new_n399_), .A2(new_n539_), .A3(new_n484_), .A4(new_n524_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n540_), .A2(new_n202_), .A3(new_n531_), .ZN(new_n541_));
  XOR2_X1   g340(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n533_), .A2(new_n543_), .ZN(G1324gat));
  AND3_X1   g343(.A1(new_n266_), .A2(new_n270_), .A3(new_n319_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n540_), .A2(new_n462_), .A3(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n485_), .A2(new_n546_), .A3(new_n525_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT100), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n548_), .A2(new_n549_), .A3(G8gat), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n549_), .B1(new_n548_), .B2(G8gat), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT39), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NOR3_X1   g353(.A1(new_n550_), .A2(new_n551_), .A3(KEYINPUT39), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n547_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n556_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g356(.A(G15gat), .ZN(new_n558_));
  INV_X1    g357(.A(new_n398_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n540_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n527_), .A2(new_n559_), .A3(new_n529_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT102), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n561_), .A2(new_n562_), .A3(G15gat), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n562_), .B1(new_n561_), .B2(G15gat), .ZN(new_n565_));
  OAI21_X1  g364(.A(KEYINPUT101), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n565_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT101), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(new_n568_), .A3(new_n563_), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n566_), .A2(new_n569_), .A3(KEYINPUT41), .ZN(new_n570_));
  AOI21_X1  g369(.A(KEYINPUT41), .B1(new_n566_), .B2(new_n569_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n560_), .B1(new_n570_), .B2(new_n571_), .ZN(G1326gat));
  INV_X1    g371(.A(G22gat), .ZN(new_n573_));
  INV_X1    g372(.A(new_n317_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n573_), .B1(new_n530_), .B2(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n575_), .B(KEYINPUT42), .Z(new_n576_));
  NAND3_X1  g375(.A1(new_n540_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(G1327gat));
  NOR2_X1   g377(.A1(new_n510_), .A2(new_n523_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n485_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT104), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n485_), .A2(KEYINPUT104), .A3(new_n579_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(G29gat), .B1(new_n584_), .B2(new_n531_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT44), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT43), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n377_), .A2(new_n379_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n397_), .A2(new_n398_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n538_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT103), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n587_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  OAI211_X1 g391(.A(KEYINPUT103), .B(KEYINPUT43), .C1(new_n399_), .C2(new_n538_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n483_), .A2(new_n524_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n586_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n596_), .A2(G29gat), .A3(new_n531_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n595_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT44), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n585_), .B1(new_n598_), .B2(new_n600_), .ZN(G1328gat));
  INV_X1    g400(.A(G36gat), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n582_), .A2(new_n602_), .A3(new_n546_), .A4(new_n583_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(KEYINPUT106), .B(KEYINPUT107), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT45), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n603_), .B(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT105), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n545_), .B1(new_n599_), .B2(KEYINPUT44), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n596_), .A2(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n607_), .B1(new_n609_), .B2(G36gat), .ZN(new_n610_));
  AOI211_X1 g409(.A(KEYINPUT105), .B(new_n602_), .C1(new_n596_), .C2(new_n608_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n606_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT46), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  OAI211_X1 g413(.A(KEYINPUT46), .B(new_n606_), .C1(new_n610_), .C2(new_n611_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(G1329gat));
  OAI21_X1  g415(.A(G43gat), .B1(new_n599_), .B2(KEYINPUT44), .ZN(new_n617_));
  AOI211_X1 g416(.A(new_n586_), .B(new_n595_), .C1(new_n592_), .C2(new_n593_), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n617_), .A2(new_n398_), .A3(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n582_), .A2(new_n559_), .A3(new_n583_), .ZN(new_n620_));
  INV_X1    g419(.A(G43gat), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(KEYINPUT108), .B1(new_n619_), .B2(new_n623_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n596_), .A2(G43gat), .A3(new_n600_), .A4(new_n559_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT108), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n625_), .A2(new_n626_), .A3(new_n622_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n624_), .A2(KEYINPUT47), .A3(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT47), .B1(new_n624_), .B2(new_n627_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1330gat));
  AOI21_X1  g429(.A(G50gat), .B1(new_n584_), .B2(new_n574_), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n596_), .A2(G50gat), .A3(new_n600_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n631_), .B1(new_n632_), .B2(new_n574_), .ZN(G1331gat));
  INV_X1    g432(.A(new_n399_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n455_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n482_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n634_), .A2(new_n637_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n638_), .A2(new_n511_), .A3(new_n524_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n639_), .A2(G57gat), .A3(new_n531_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT109), .Z(new_n641_));
  NOR3_X1   g440(.A1(new_n638_), .A2(new_n524_), .A3(new_n539_), .ZN(new_n642_));
  AOI21_X1  g441(.A(G57gat), .B1(new_n642_), .B2(new_n531_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n641_), .A2(new_n643_), .ZN(G1332gat));
  INV_X1    g443(.A(G64gat), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n642_), .A2(new_n645_), .A3(new_n546_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n639_), .B2(new_n546_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT111), .Z(new_n648_));
  XNOR2_X1  g447(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n648_), .A2(new_n649_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n646_), .B1(new_n650_), .B2(new_n651_), .ZN(G1333gat));
  INV_X1    g451(.A(G71gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(new_n639_), .B2(new_n559_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT49), .Z(new_n655_));
  NAND3_X1  g454(.A1(new_n642_), .A2(new_n653_), .A3(new_n559_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1334gat));
  INV_X1    g456(.A(G78gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n658_), .B1(new_n639_), .B2(new_n574_), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n659_), .B(KEYINPUT50), .Z(new_n660_));
  NAND3_X1  g459(.A1(new_n642_), .A2(new_n658_), .A3(new_n574_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1335gat));
  NAND2_X1  g461(.A1(new_n455_), .A2(new_n482_), .ZN(new_n663_));
  AOI211_X1 g462(.A(new_n523_), .B(new_n663_), .C1(new_n592_), .C2(new_n593_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(new_n531_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n638_), .A2(new_n510_), .A3(new_n523_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n353_), .A2(G85gat), .ZN(new_n667_));
  AOI22_X1  g466(.A1(new_n665_), .A2(G85gat), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT112), .ZN(G1336gat));
  AOI21_X1  g468(.A(G92gat), .B1(new_n666_), .B2(new_n546_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT113), .Z(new_n671_));
  AND2_X1   g470(.A1(new_n546_), .A2(G92gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n664_), .B2(new_n672_), .ZN(G1337gat));
  NAND3_X1  g472(.A1(new_n666_), .A2(new_n401_), .A3(new_n559_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT114), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n664_), .A2(new_n559_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n676_), .B2(G99gat), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT51), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n677_), .B(new_n678_), .ZN(G1338gat));
  NAND3_X1  g478(.A1(new_n666_), .A2(new_n402_), .A3(new_n574_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT52), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n664_), .A2(new_n574_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n682_), .B2(G106gat), .ZN(new_n683_));
  AOI211_X1 g482(.A(KEYINPUT52), .B(new_n402_), .C1(new_n664_), .C2(new_n574_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n680_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g485(.A1(new_n320_), .A2(new_n398_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT57), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n482_), .A2(new_n451_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n434_), .A2(new_n439_), .A3(new_n436_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT115), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n690_), .A2(new_n691_), .A3(KEYINPUT55), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n691_), .B1(new_n690_), .B2(KEYINPUT55), .ZN(new_n693_));
  OAI22_X1  g492(.A1(new_n692_), .A2(new_n693_), .B1(new_n439_), .B2(new_n437_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n690_), .A2(KEYINPUT55), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT115), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n690_), .A2(new_n691_), .A3(KEYINPUT55), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n696_), .A2(new_n440_), .A3(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n694_), .A2(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(KEYINPUT56), .B1(new_n699_), .B2(new_n448_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT56), .ZN(new_n701_));
  AOI211_X1 g500(.A(new_n701_), .B(new_n449_), .C1(new_n694_), .C2(new_n698_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n689_), .B1(new_n700_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT116), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n473_), .A2(new_n471_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n470_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n478_), .B(new_n706_), .C1(new_n707_), .C2(new_n471_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n708_), .A2(new_n481_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n709_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n710_));
  OAI211_X1 g509(.A(KEYINPUT116), .B(new_n689_), .C1(new_n700_), .C2(new_n702_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n705_), .A2(new_n710_), .A3(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n510_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n688_), .B1(new_n713_), .B2(KEYINPUT117), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT117), .ZN(new_n715_));
  AOI211_X1 g514(.A(new_n715_), .B(KEYINPUT57), .C1(new_n712_), .C2(new_n510_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n714_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT118), .ZN(new_n718_));
  OR3_X1    g517(.A1(new_n700_), .A2(new_n702_), .A3(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n451_), .B1(new_n702_), .B2(new_n718_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n719_), .A2(new_n720_), .A3(new_n709_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT58), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n719_), .A2(new_n720_), .A3(KEYINPUT58), .A4(new_n709_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n723_), .A2(new_n539_), .A3(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n523_), .B1(new_n717_), .B2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n538_), .A2(new_n482_), .A3(new_n523_), .ZN(new_n727_));
  OR3_X1    g526(.A1(new_n727_), .A2(KEYINPUT54), .A3(new_n455_), .ZN(new_n728_));
  OAI21_X1  g527(.A(KEYINPUT54), .B1(new_n727_), .B2(new_n455_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n531_), .B(new_n687_), .C1(new_n726_), .C2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT59), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n713_), .A2(KEYINPUT117), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT57), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n713_), .A2(KEYINPUT117), .A3(new_n688_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(new_n725_), .A3(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n524_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(new_n730_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT59), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n739_), .A2(new_n740_), .A3(new_n531_), .A4(new_n687_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n482_), .A2(new_n324_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT119), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n733_), .A2(new_n741_), .A3(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n324_), .B1(new_n732_), .B2(new_n482_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT120), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT120), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n744_), .A2(new_n748_), .A3(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1340gat));
  INV_X1    g549(.A(KEYINPUT60), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n751_), .B1(new_n635_), .B2(G120gat), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n739_), .A2(new_n531_), .A3(new_n687_), .A4(new_n752_), .ZN(new_n753_));
  AND4_X1   g552(.A1(new_n455_), .A2(new_n733_), .A3(new_n741_), .A4(new_n753_), .ZN(new_n754_));
  OAI22_X1  g553(.A1(new_n754_), .A2(new_n328_), .B1(KEYINPUT60), .B2(new_n753_), .ZN(G1341gat));
  NAND4_X1  g554(.A1(new_n733_), .A2(new_n741_), .A3(G127gat), .A4(new_n523_), .ZN(new_n756_));
  INV_X1    g555(.A(G127gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n757_), .B1(new_n732_), .B2(new_n524_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1342gat));
  NAND4_X1  g558(.A1(new_n733_), .A2(new_n741_), .A3(G134gat), .A4(new_n539_), .ZN(new_n760_));
  INV_X1    g559(.A(G134gat), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n761_), .B1(new_n732_), .B2(new_n510_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1343gat));
  NOR2_X1   g562(.A1(new_n546_), .A2(new_n317_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n739_), .A2(new_n531_), .A3(new_n398_), .A4(new_n764_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n765_), .A2(new_n482_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(new_n279_), .ZN(G1344gat));
  NOR2_X1   g566(.A1(new_n765_), .A2(new_n635_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(new_n280_), .ZN(G1345gat));
  NOR2_X1   g568(.A1(new_n765_), .A2(new_n524_), .ZN(new_n770_));
  XOR2_X1   g569(.A(KEYINPUT61), .B(G155gat), .Z(new_n771_));
  XNOR2_X1  g570(.A(new_n770_), .B(new_n771_), .ZN(G1346gat));
  NOR3_X1   g571(.A1(new_n765_), .A2(new_n502_), .A3(new_n538_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n502_), .B1(new_n765_), .B2(new_n510_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT121), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  OAI211_X1 g575(.A(KEYINPUT121), .B(new_n502_), .C1(new_n765_), .C2(new_n510_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(G1347gat));
  NOR2_X1   g577(.A1(new_n545_), .A2(new_n378_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n739_), .A2(new_n636_), .A3(new_n317_), .A4(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(G169gat), .ZN(new_n781_));
  XOR2_X1   g580(.A(KEYINPUT122), .B(KEYINPUT62), .Z(new_n782_));
  NOR2_X1   g581(.A1(new_n782_), .A2(KEYINPUT123), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  XOR2_X1   g583(.A(KEYINPUT22), .B(G169gat), .Z(new_n785_));
  NAND2_X1  g584(.A1(new_n782_), .A2(KEYINPUT123), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n780_), .A2(G169gat), .A3(new_n786_), .ZN(new_n787_));
  OAI221_X1 g586(.A(new_n784_), .B1(new_n780_), .B2(new_n785_), .C1(new_n783_), .C2(new_n787_), .ZN(G1348gat));
  AOI21_X1  g587(.A(new_n731_), .B1(new_n524_), .B2(new_n737_), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT124), .B1(new_n789_), .B2(new_n574_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT124), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n739_), .A2(new_n791_), .A3(new_n317_), .ZN(new_n792_));
  INV_X1    g591(.A(G176gat), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n635_), .A2(new_n793_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n790_), .A2(new_n792_), .A3(new_n779_), .A4(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n739_), .A2(new_n317_), .A3(new_n779_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n793_), .B1(new_n796_), .B2(new_n635_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n795_), .A2(new_n797_), .ZN(G1349gat));
  NAND4_X1  g597(.A1(new_n790_), .A2(new_n792_), .A3(new_n523_), .A4(new_n779_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n209_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT125), .ZN(new_n801_));
  INV_X1    g600(.A(new_n211_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n739_), .A2(new_n317_), .A3(new_n802_), .A4(new_n779_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n801_), .B1(new_n803_), .B2(new_n524_), .ZN(new_n804_));
  OR3_X1    g603(.A1(new_n803_), .A2(new_n801_), .A3(new_n524_), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n800_), .A2(new_n804_), .A3(new_n805_), .ZN(G1350gat));
  OAI21_X1  g605(.A(G190gat), .B1(new_n796_), .B2(new_n538_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n511_), .A2(new_n208_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n807_), .B1(new_n796_), .B2(new_n808_), .ZN(G1351gat));
  NOR2_X1   g608(.A1(new_n545_), .A2(new_n559_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n380_), .B(new_n810_), .C1(new_n726_), .C2(new_n731_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT126), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n739_), .A2(KEYINPUT126), .A3(new_n380_), .A4(new_n810_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  AND3_X1   g614(.A1(new_n815_), .A2(G197gat), .A3(new_n636_), .ZN(new_n816_));
  AOI21_X1  g615(.A(G197gat), .B1(new_n815_), .B2(new_n636_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(G1352gat));
  AOI21_X1  g617(.A(new_n635_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n819_));
  INV_X1    g618(.A(G204gat), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n819_), .B(new_n820_), .ZN(G1353gat));
  XNOR2_X1  g620(.A(KEYINPUT63), .B(G211gat), .ZN(new_n822_));
  AOI211_X1 g621(.A(new_n524_), .B(new_n822_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n815_), .A2(new_n523_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n823_), .B1(new_n824_), .B2(new_n825_), .ZN(G1354gat));
  AOI21_X1  g625(.A(G218gat), .B1(new_n815_), .B2(new_n511_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n539_), .A2(G218gat), .ZN(new_n828_));
  XOR2_X1   g627(.A(new_n828_), .B(KEYINPUT127), .Z(new_n829_));
  AOI21_X1  g628(.A(new_n827_), .B1(new_n815_), .B2(new_n829_), .ZN(G1355gat));
endmodule


