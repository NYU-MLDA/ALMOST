//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 0 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n857_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT68), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G71gat), .B(G78gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n205_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n203_), .B(KEYINPUT68), .ZN(new_n210_));
  INV_X1    g009(.A(new_n208_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(G15gat), .B(G22gat), .Z(new_n214_));
  NAND2_X1  g013(.A1(G1gat), .A2(G8gat), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n214_), .B1(KEYINPUT14), .B2(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(new_n216_), .B(KEYINPUT72), .Z(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT73), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n216_), .B(KEYINPUT72), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT73), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n218_), .A2(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(G1gat), .B(G8gat), .Z(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n218_), .A2(new_n223_), .A3(new_n221_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(G231gat), .ZN(new_n228_));
  INV_X1    g027(.A(G233gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n227_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n230_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n232_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n213_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n226_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n223_), .B1(new_n218_), .B2(new_n221_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(new_n232_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n233_), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n209_), .A2(new_n212_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G127gat), .B(G155gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT16), .ZN(new_n243_));
  XOR2_X1   g042(.A(G183gat), .B(G211gat), .Z(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT17), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n234_), .A2(new_n241_), .A3(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT74), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n234_), .A2(new_n241_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n245_), .B(KEYINPUT17), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT75), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT75), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n251_), .A2(new_n255_), .A3(new_n252_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n250_), .A2(new_n254_), .A3(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n255_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n252_), .ZN(new_n259_));
  AOI211_X1 g058(.A(KEYINPUT75), .B(new_n259_), .C1(new_n234_), .C2(new_n241_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n249_), .B1(new_n258_), .B2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n257_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT37), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G190gat), .B(G218gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G134gat), .B(G162gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n266_), .B(KEYINPUT36), .Z(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT71), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT8), .ZN(new_n269_));
  NOR2_X1   g068(.A1(G99gat), .A2(G106gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT7), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G99gat), .A2(G106gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT6), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT6), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n274_), .A2(G99gat), .A3(G106gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n271_), .A2(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(G85gat), .B(G92gat), .Z(new_n278_));
  AOI21_X1  g077(.A(new_n269_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n276_), .B(KEYINPUT67), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n271_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n278_), .A2(new_n269_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n279_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(KEYINPUT10), .B(G99gat), .Z(new_n285_));
  INV_X1    g084(.A(G106gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT65), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT66), .B(G85gat), .ZN(new_n290_));
  INV_X1    g089(.A(G92gat), .ZN(new_n291_));
  NOR3_X1   g090(.A1(new_n290_), .A2(KEYINPUT9), .A3(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n292_), .B1(KEYINPUT9), .B2(new_n278_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n289_), .A2(new_n280_), .A3(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G29gat), .B(G36gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G43gat), .B(G50gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n284_), .A2(new_n294_), .A3(new_n297_), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n298_), .B(KEYINPUT70), .Z(new_n299_));
  NAND2_X1  g098(.A1(G232gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT34), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT35), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n284_), .A2(new_n294_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n297_), .B(KEYINPUT15), .ZN(new_n307_));
  AOI22_X1  g106(.A1(new_n306_), .A2(new_n307_), .B1(new_n303_), .B2(new_n302_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n299_), .A2(new_n305_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n305_), .B1(new_n299_), .B2(new_n308_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n268_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n311_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n266_), .A2(KEYINPUT36), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n313_), .A2(new_n314_), .A3(new_n309_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n263_), .B1(new_n312_), .B2(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n267_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n315_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n316_), .B1(new_n319_), .B2(new_n263_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n262_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n294_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n240_), .B1(new_n322_), .B2(new_n283_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n284_), .A2(new_n294_), .A3(new_n213_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G230gat), .A2(G233gat), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n326_), .B(KEYINPUT64), .Z(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT69), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT69), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n325_), .A2(new_n330_), .A3(new_n327_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n323_), .A2(new_n324_), .A3(KEYINPUT12), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT12), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n306_), .A2(new_n334_), .A3(new_n240_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n327_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G120gat), .B(G148gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT5), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G176gat), .B(G204gat), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n338_), .B(new_n339_), .Z(new_n340_));
  OR3_X1    g139(.A1(new_n332_), .A2(new_n336_), .A3(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n340_), .B1(new_n332_), .B2(new_n336_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT13), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(KEYINPUT13), .B1(new_n341_), .B2(new_n342_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n321_), .A2(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT76), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n297_), .B(KEYINPUT77), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n350_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n350_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n225_), .A2(new_n226_), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n351_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G229gat), .A2(G233gat), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n237_), .A2(KEYINPUT78), .A3(new_n352_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n355_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n237_), .A2(new_n307_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n360_), .A2(new_n356_), .A3(new_n351_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G113gat), .B(G141gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G169gat), .B(G197gat), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n362_), .B(new_n363_), .Z(new_n364_));
  NAND3_X1  g163(.A1(new_n359_), .A2(new_n361_), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n364_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  XOR2_X1   g167(.A(KEYINPUT99), .B(KEYINPUT18), .Z(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT100), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G8gat), .B(G36gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G64gat), .B(G92gat), .ZN(new_n373_));
  XOR2_X1   g172(.A(new_n372_), .B(new_n373_), .Z(new_n374_));
  INV_X1    g173(.A(KEYINPUT20), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT79), .B(G190gat), .ZN(new_n376_));
  INV_X1    g175(.A(G183gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G183gat), .A2(G190gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT23), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT23), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(G183gat), .A3(G190gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  AOI22_X1  g182(.A1(new_n378_), .A2(new_n383_), .B1(G169gat), .B2(G176gat), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT22), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n385_), .A2(G169gat), .ZN(new_n386_));
  INV_X1    g185(.A(G169gat), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n387_), .A2(KEYINPUT22), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT83), .B1(new_n386_), .B2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT84), .B(G176gat), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n389_), .B(new_n390_), .C1(KEYINPUT83), .C2(new_n386_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n384_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(G176gat), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n387_), .A2(new_n393_), .A3(KEYINPUT81), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT81), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n395_), .B1(G169gat), .B2(G176gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G169gat), .A2(G176gat), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n394_), .A2(new_n396_), .A3(KEYINPUT24), .A4(new_n397_), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n394_), .A2(new_n396_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n398_), .B1(new_n399_), .B2(KEYINPUT24), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n382_), .A2(KEYINPUT82), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT82), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n402_), .A2(new_n381_), .A3(G183gat), .A4(G190gat), .ZN(new_n403_));
  AOI22_X1  g202(.A1(new_n401_), .A2(new_n403_), .B1(KEYINPUT23), .B2(new_n379_), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n400_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT25), .B(G183gat), .ZN(new_n406_));
  INV_X1    g205(.A(G190gat), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n406_), .B1(KEYINPUT26), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n376_), .A2(KEYINPUT26), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT80), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT80), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n376_), .A2(new_n411_), .A3(KEYINPUT26), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n408_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n392_), .B1(new_n405_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT21), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G197gat), .B(G204gat), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT92), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G211gat), .B(G218gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n419_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n416_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n415_), .B1(new_n420_), .B2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT21), .B1(new_n418_), .B2(new_n419_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n375_), .B1(new_n414_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G226gat), .A2(G233gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT19), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT97), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n430_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n387_), .A2(KEYINPUT22), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n385_), .A2(G169gat), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(new_n433_), .A3(KEYINPUT97), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n431_), .A2(new_n390_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n397_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(G183gat), .A2(G190gat), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n404_), .A2(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT95), .ZN(new_n441_));
  NOR2_X1   g240(.A1(G169gat), .A2(G176gat), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT24), .ZN(new_n443_));
  AOI221_X4 g242(.A(new_n441_), .B1(new_n442_), .B2(new_n443_), .C1(new_n380_), .C2(new_n382_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n443_), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT95), .B1(new_n383_), .B2(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(KEYINPUT26), .B(G190gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n406_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(new_n398_), .ZN(new_n450_));
  NOR3_X1   g249(.A1(new_n447_), .A2(KEYINPUT96), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT96), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n383_), .A2(new_n445_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n441_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n383_), .A2(KEYINPUT95), .A3(new_n445_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n450_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n452_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n440_), .B1(new_n451_), .B2(new_n458_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n426_), .B(new_n429_), .C1(new_n425_), .C2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT20), .B1(new_n414_), .B2(new_n425_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT98), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n459_), .A2(new_n462_), .A3(new_n425_), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT96), .B1(new_n447_), .B2(new_n450_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n456_), .A2(new_n452_), .A3(new_n457_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n439_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n425_), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT98), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n461_), .B1(new_n463_), .B2(new_n468_), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n374_), .B(new_n460_), .C1(new_n469_), .C2(new_n429_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT107), .ZN(new_n471_));
  INV_X1    g270(.A(new_n461_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n462_), .B1(new_n459_), .B2(new_n425_), .ZN(new_n473_));
  NOR3_X1   g272(.A1(new_n466_), .A2(KEYINPUT98), .A3(new_n467_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n472_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(new_n428_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT107), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n476_), .A2(new_n477_), .A3(new_n374_), .A4(new_n460_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n374_), .ZN(new_n479_));
  AOI211_X1 g278(.A(new_n428_), .B(new_n461_), .C1(new_n463_), .C2(new_n468_), .ZN(new_n480_));
  OAI211_X1 g279(.A(new_n467_), .B(new_n440_), .C1(new_n447_), .C2(new_n450_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n429_), .B1(new_n426_), .B2(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n479_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n471_), .A2(new_n478_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT27), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n460_), .B1(new_n469_), .B2(new_n429_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n479_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT27), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(new_n488_), .A3(new_n470_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n485_), .A2(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G71gat), .B(G99gat), .Z(new_n491_));
  XNOR2_X1  g290(.A(G15gat), .B(G43gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n414_), .B(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(G127gat), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n495_), .A2(G134gat), .ZN(new_n496_));
  INV_X1    g295(.A(G134gat), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n497_), .A2(G127gat), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT86), .B1(new_n496_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(G127gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n495_), .A2(G134gat), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT86), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G113gat), .B(G120gat), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n499_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n504_), .B1(new_n499_), .B2(new_n503_), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n494_), .B(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G227gat), .A2(G233gat), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n509_), .B(KEYINPUT85), .Z(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT30), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT31), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n508_), .B(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(KEYINPUT90), .A2(G228gat), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(KEYINPUT90), .A2(G228gat), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n229_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT91), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT91), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n423_), .A2(new_n424_), .A3(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(G141gat), .A2(G148gat), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G141gat), .A2(G148gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G155gat), .A2(G162gat), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n526_), .A2(KEYINPUT1), .ZN(new_n527_));
  NOR2_X1   g326(.A1(G155gat), .A2(G162gat), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n526_), .B1(new_n528_), .B2(KEYINPUT1), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n527_), .B1(new_n529_), .B2(KEYINPUT87), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT1), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n531_), .B1(G155gat), .B2(G162gat), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT87), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(new_n533_), .A3(new_n526_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n525_), .B1(new_n530_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT3), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n522_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT2), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n524_), .A2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n537_), .A2(new_n539_), .A3(new_n540_), .A4(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n528_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n543_), .A2(new_n526_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT88), .B1(new_n535_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT88), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n532_), .A2(new_n533_), .A3(new_n526_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n533_), .B1(new_n532_), .B2(new_n526_), .ZN(new_n550_));
  NOR3_X1   g349(.A1(new_n549_), .A2(new_n550_), .A3(new_n527_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n548_), .B(new_n545_), .C1(new_n551_), .C2(new_n525_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n547_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT29), .ZN(new_n554_));
  OAI221_X1 g353(.A(new_n519_), .B1(new_n521_), .B2(new_n518_), .C1(new_n553_), .C2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(G78gat), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n535_), .A2(new_n546_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT93), .B(KEYINPUT29), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n425_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(new_n518_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n555_), .A2(new_n556_), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n556_), .B1(new_n555_), .B2(new_n560_), .ZN(new_n563_));
  OAI21_X1  g362(.A(G106gat), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n563_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n565_), .A2(new_n286_), .A3(new_n561_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n553_), .A2(new_n554_), .ZN(new_n568_));
  XOR2_X1   g367(.A(G22gat), .B(G50gat), .Z(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n568_), .A2(new_n569_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n571_), .A2(new_n572_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n574_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n576_), .A2(new_n577_), .A3(KEYINPUT94), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT94), .ZN(new_n579_));
  INV_X1    g378(.A(new_n577_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n579_), .B1(new_n580_), .B2(new_n575_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n567_), .A2(new_n578_), .A3(new_n581_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n580_), .A2(new_n575_), .A3(new_n579_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n583_), .A2(new_n564_), .A3(new_n566_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n514_), .B1(new_n582_), .B2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G1gat), .B(G29gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(G85gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT0), .B(G57gat), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n587_), .B(new_n588_), .Z(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n547_), .A2(new_n552_), .A3(new_n507_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT103), .B(KEYINPUT4), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G225gat), .A2(G233gat), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n505_), .A2(new_n506_), .ZN(new_n597_));
  AOI21_X1  g396(.A(KEYINPUT101), .B1(new_n557_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n591_), .A2(new_n598_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n547_), .A2(new_n552_), .A3(new_n507_), .A4(KEYINPUT101), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT4), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT102), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n601_), .A2(KEYINPUT102), .A3(KEYINPUT4), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n596_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n601_), .A2(new_n594_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n590_), .B1(new_n606_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT106), .ZN(new_n610_));
  INV_X1    g409(.A(new_n596_), .ZN(new_n611_));
  AOI21_X1  g410(.A(KEYINPUT102), .B1(new_n601_), .B2(KEYINPUT4), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT4), .ZN(new_n613_));
  AOI211_X1 g412(.A(new_n603_), .B(new_n613_), .C1(new_n599_), .C2(new_n600_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n611_), .B1(new_n612_), .B2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n615_), .A2(new_n607_), .A3(new_n589_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n609_), .A2(new_n610_), .A3(new_n616_), .ZN(new_n617_));
  OAI211_X1 g416(.A(KEYINPUT106), .B(new_n590_), .C1(new_n606_), .C2(new_n608_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n490_), .A2(new_n585_), .A3(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(KEYINPUT108), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n485_), .A2(new_n489_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT108), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(new_n623_), .A3(new_n585_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n621_), .A2(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n480_), .A2(new_n482_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n374_), .A2(KEYINPUT32), .ZN(new_n627_));
  MUX2_X1   g426(.A(new_n626_), .B(new_n486_), .S(new_n627_), .Z(new_n628_));
  NAND3_X1  g427(.A1(new_n617_), .A2(new_n618_), .A3(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n582_), .A2(new_n584_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n487_), .A2(new_n470_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n593_), .A2(new_n594_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n632_), .B1(new_n612_), .B2(new_n614_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(KEYINPUT105), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT105), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n635_), .B(new_n632_), .C1(new_n612_), .C2(new_n614_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n589_), .B1(new_n601_), .B2(new_n595_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n634_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT104), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n639_), .A2(KEYINPUT33), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n616_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n640_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n615_), .A2(new_n607_), .A3(new_n589_), .A4(new_n642_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n631_), .A2(new_n638_), .A3(new_n641_), .A4(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n629_), .A2(new_n630_), .A3(new_n644_), .ZN(new_n645_));
  OAI211_X1 g444(.A(new_n645_), .B(new_n514_), .C1(new_n630_), .C2(new_n622_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n368_), .B1(new_n625_), .B2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n349_), .A2(new_n647_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n648_), .A2(G1gat), .A3(new_n619_), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n649_), .A2(KEYINPUT109), .A3(KEYINPUT38), .ZN(new_n650_));
  AOI21_X1  g449(.A(KEYINPUT109), .B1(new_n649_), .B2(KEYINPUT38), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT38), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n319_), .B1(new_n625_), .B2(new_n646_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n257_), .A2(new_n261_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n368_), .ZN(new_n655_));
  AND4_X1   g454(.A1(new_n653_), .A2(new_n654_), .A3(new_n655_), .A4(new_n347_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n619_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n652_), .B1(new_n658_), .B2(G1gat), .ZN(new_n659_));
  OAI22_X1  g458(.A1(new_n650_), .A2(new_n651_), .B1(new_n659_), .B2(new_n649_), .ZN(G1324gat));
  OR3_X1    g459(.A1(new_n648_), .A2(G8gat), .A3(new_n490_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n490_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n656_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(G8gat), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n664_), .A2(KEYINPUT39), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(KEYINPUT39), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n661_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT40), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(G1325gat));
  INV_X1    g468(.A(G15gat), .ZN(new_n670_));
  INV_X1    g469(.A(new_n514_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n656_), .B2(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT41), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n670_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n673_), .B1(new_n648_), .B2(new_n674_), .ZN(G1326gat));
  INV_X1    g474(.A(G22gat), .ZN(new_n676_));
  INV_X1    g475(.A(new_n630_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n656_), .B2(new_n677_), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT42), .Z(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n676_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT110), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n679_), .B1(new_n648_), .B2(new_n681_), .ZN(G1327gat));
  NOR2_X1   g481(.A1(new_n654_), .A2(new_n318_), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n647_), .A2(new_n347_), .A3(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G29gat), .B1(new_n684_), .B2(new_n657_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n316_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n686_), .B1(KEYINPUT37), .B2(new_n318_), .ZN(new_n687_));
  AOI211_X1 g486(.A(KEYINPUT43), .B(new_n687_), .C1(new_n625_), .C2(new_n646_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n623_), .B1(new_n622_), .B2(new_n585_), .ZN(new_n690_));
  AND4_X1   g489(.A1(new_n623_), .A2(new_n490_), .A3(new_n585_), .A4(new_n619_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n645_), .A2(new_n514_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n622_), .A2(new_n630_), .ZN(new_n693_));
  OAI22_X1  g492(.A1(new_n690_), .A2(new_n691_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n689_), .B1(new_n694_), .B2(new_n320_), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n688_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n347_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n654_), .A2(new_n697_), .A3(new_n368_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n696_), .A2(KEYINPUT44), .A3(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(KEYINPUT44), .B1(new_n696_), .B2(new_n698_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n657_), .A2(G29gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n685_), .B1(new_n702_), .B2(new_n703_), .ZN(G1328gat));
  INV_X1    g503(.A(KEYINPUT46), .ZN(new_n705_));
  INV_X1    g504(.A(G36gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n702_), .B2(new_n662_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n684_), .A2(new_n706_), .A3(new_n662_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT45), .Z(new_n709_));
  OAI21_X1  g508(.A(new_n705_), .B1(new_n707_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n701_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n699_), .ZN(new_n712_));
  OAI21_X1  g511(.A(G36gat), .B1(new_n712_), .B2(new_n490_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n709_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n713_), .A2(KEYINPUT46), .A3(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n710_), .A2(new_n715_), .ZN(G1329gat));
  AOI21_X1  g515(.A(G43gat), .B1(new_n684_), .B2(new_n671_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT111), .Z(new_n718_));
  NAND2_X1  g517(.A1(new_n671_), .A2(G43gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n712_), .B2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT47), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT47), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n718_), .B(new_n722_), .C1(new_n712_), .C2(new_n719_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(G1330gat));
  AOI21_X1  g523(.A(G50gat), .B1(new_n684_), .B2(new_n677_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n677_), .A2(G50gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n702_), .B2(new_n726_), .ZN(G1331gat));
  NOR3_X1   g526(.A1(new_n262_), .A2(new_n347_), .A3(new_n655_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n653_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(G57gat), .B1(new_n730_), .B2(new_n619_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n655_), .B1(new_n625_), .B2(new_n646_), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n732_), .A2(new_n697_), .A3(new_n321_), .ZN(new_n733_));
  INV_X1    g532(.A(G57gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(new_n734_), .A3(new_n657_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n731_), .A2(new_n735_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT112), .Z(G1332gat));
  OAI21_X1  g536(.A(G64gat), .B1(new_n730_), .B2(new_n490_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n738_), .B(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n490_), .A2(G64gat), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT114), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n733_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n740_), .A2(new_n743_), .ZN(G1333gat));
  INV_X1    g543(.A(G71gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n729_), .B2(new_n671_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT49), .Z(new_n747_));
  NAND3_X1  g546(.A1(new_n733_), .A2(new_n745_), .A3(new_n671_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1334gat));
  AOI21_X1  g548(.A(new_n556_), .B1(new_n729_), .B2(new_n677_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT50), .Z(new_n751_));
  NAND3_X1  g550(.A1(new_n733_), .A2(new_n556_), .A3(new_n677_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1335gat));
  AND3_X1   g552(.A1(new_n732_), .A2(new_n697_), .A3(new_n683_), .ZN(new_n754_));
  AOI21_X1  g553(.A(G85gat), .B1(new_n754_), .B2(new_n657_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n654_), .A2(new_n655_), .A3(new_n347_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n696_), .A2(new_n756_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n619_), .A2(new_n290_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n755_), .B1(new_n757_), .B2(new_n758_), .ZN(G1336gat));
  NAND3_X1  g558(.A1(new_n754_), .A2(new_n291_), .A3(new_n662_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n757_), .A2(new_n662_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(new_n291_), .ZN(G1337gat));
  INV_X1    g561(.A(G99gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n763_), .B1(new_n757_), .B2(new_n671_), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n754_), .A2(new_n285_), .A3(new_n671_), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g566(.A1(new_n754_), .A2(new_n286_), .A3(new_n677_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n677_), .B(new_n756_), .C1(new_n688_), .C2(new_n695_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n769_), .A2(new_n770_), .A3(G106gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n769_), .B2(G106gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT116), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT116), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n775_), .B(new_n768_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n774_), .A2(new_n776_), .A3(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n778_), .A2(new_n779_), .ZN(G1339gat));
  INV_X1    g579(.A(new_n585_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n355_), .A2(new_n356_), .A3(new_n358_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n356_), .B1(new_n227_), .B2(new_n350_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n364_), .B1(new_n783_), .B2(new_n360_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n343_), .A2(new_n365_), .A3(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n333_), .A2(new_n335_), .ZN(new_n788_));
  OAI211_X1 g587(.A(KEYINPUT117), .B(new_n787_), .C1(new_n788_), .C2(new_n327_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT117), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n790_), .B1(new_n336_), .B2(KEYINPUT55), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n788_), .A2(new_n327_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n336_), .A2(KEYINPUT55), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n789_), .A2(new_n791_), .A3(new_n792_), .A4(new_n793_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n794_), .A2(KEYINPUT56), .A3(new_n340_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT56), .B1(new_n794_), .B2(new_n340_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n341_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n786_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT118), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n799_), .A2(new_n318_), .A3(new_n801_), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n341_), .A2(new_n365_), .A3(new_n785_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n803_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT58), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n803_), .B(KEYINPUT58), .C1(new_n795_), .C2(new_n796_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n806_), .A2(new_n320_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n802_), .A2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n801_), .B1(new_n799_), .B2(new_n318_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n262_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n654_), .A2(new_n687_), .A3(new_n368_), .A4(new_n347_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT54), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n321_), .A2(new_n814_), .A3(new_n368_), .A4(new_n347_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n781_), .B1(new_n811_), .B2(new_n816_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n662_), .A2(new_n619_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT59), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n817_), .B(new_n818_), .C1(KEYINPUT119), .C2(new_n819_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n817_), .A2(new_n818_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n820_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(G113gat), .B1(new_n823_), .B2(new_n368_), .ZN(new_n824_));
  INV_X1    g623(.A(G113gat), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n821_), .A2(new_n825_), .A3(new_n655_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(G1340gat));
  XNOR2_X1  g626(.A(KEYINPUT120), .B(G120gat), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(new_n823_), .B2(new_n347_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT60), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n828_), .B1(new_n697_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT121), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT121), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n833_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n821_), .B(new_n832_), .C1(new_n831_), .C2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n829_), .A2(new_n835_), .ZN(G1341gat));
  NOR2_X1   g635(.A1(new_n262_), .A2(KEYINPUT122), .ZN(new_n837_));
  MUX2_X1   g636(.A(KEYINPUT122), .B(new_n837_), .S(G127gat), .Z(new_n838_));
  OAI211_X1 g637(.A(new_n820_), .B(new_n838_), .C1(new_n821_), .C2(new_n822_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n821_), .A2(new_n654_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(G127gat), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT123), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT123), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n839_), .B(new_n843_), .C1(new_n840_), .C2(G127gat), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n844_), .ZN(G1342gat));
  OAI21_X1  g644(.A(G134gat), .B1(new_n823_), .B2(new_n687_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n821_), .A2(new_n497_), .A3(new_n319_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(G1343gat));
  AOI211_X1 g647(.A(new_n630_), .B(new_n671_), .C1(new_n811_), .C2(new_n816_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n818_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT124), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n849_), .A2(KEYINPUT124), .A3(new_n818_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n368_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(G141gat), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n854_), .B(new_n855_), .ZN(G1344gat));
  AOI21_X1  g655(.A(new_n347_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n857_));
  INV_X1    g656(.A(G148gat), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(G1345gat));
  AOI21_X1  g658(.A(new_n262_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT61), .B(G155gat), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n860_), .B(new_n862_), .ZN(G1346gat));
  NAND2_X1  g662(.A1(new_n852_), .A2(new_n853_), .ZN(new_n864_));
  INV_X1    g663(.A(G162gat), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n864_), .A2(new_n865_), .A3(new_n319_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n687_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(new_n865_), .ZN(G1347gat));
  INV_X1    g667(.A(KEYINPUT126), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n811_), .A2(new_n816_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n657_), .A2(new_n490_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n870_), .A2(new_n585_), .A3(new_n655_), .A4(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT125), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n817_), .A2(KEYINPUT125), .A3(new_n655_), .A4(new_n871_), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n874_), .A2(KEYINPUT62), .A3(G169gat), .A4(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n817_), .A2(new_n871_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n878_), .A2(new_n431_), .A3(new_n434_), .A4(new_n655_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n876_), .A2(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n387_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n881_));
  AOI21_X1  g680(.A(KEYINPUT62), .B1(new_n881_), .B2(new_n875_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n869_), .B1(new_n880_), .B2(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n874_), .A2(G169gat), .A3(new_n875_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT62), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n886_), .A2(KEYINPUT126), .A3(new_n879_), .A4(new_n876_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n883_), .A2(new_n887_), .ZN(G1348gat));
  NAND2_X1  g687(.A1(new_n870_), .A2(new_n630_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(KEYINPUT127), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n657_), .A2(new_n490_), .A3(new_n514_), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n697_), .A2(new_n891_), .A3(G176gat), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n878_), .A2(new_n697_), .ZN(new_n893_));
  AOI22_X1  g692(.A1(new_n890_), .A2(new_n892_), .B1(new_n893_), .B2(new_n390_), .ZN(G1349gat));
  NOR3_X1   g693(.A1(new_n877_), .A2(new_n406_), .A3(new_n262_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n890_), .A2(new_n654_), .A3(new_n891_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n895_), .B1(new_n896_), .B2(new_n377_), .ZN(G1350gat));
  OAI21_X1  g696(.A(G190gat), .B1(new_n877_), .B2(new_n687_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n319_), .A2(new_n448_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n877_), .B2(new_n899_), .ZN(G1351gat));
  AND2_X1   g699(.A1(new_n849_), .A2(new_n871_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n655_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n697_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g704(.A1(new_n901_), .A2(new_n654_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n907_));
  AND2_X1   g706(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n906_), .A2(new_n907_), .A3(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n909_), .B1(new_n906_), .B2(new_n907_), .ZN(G1354gat));
  INV_X1    g709(.A(G218gat), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n901_), .A2(new_n911_), .A3(new_n319_), .ZN(new_n912_));
  AND2_X1   g711(.A1(new_n901_), .A2(new_n320_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n911_), .ZN(G1355gat));
endmodule


