//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 0 0 0 0 1 1 1 0 1 1 0 1 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 1 0 1 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n773_, new_n774_, new_n775_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n897_, new_n898_, new_n900_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G29gat), .B(G36gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G43gat), .B(G50gat), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n204_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT15), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G15gat), .B(G22gat), .ZN(new_n209_));
  INV_X1    g008(.A(G1gat), .ZN(new_n210_));
  INV_X1    g009(.A(G8gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT14), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G1gat), .B(G8gat), .ZN(new_n214_));
  XOR2_X1   g013(.A(new_n213_), .B(new_n214_), .Z(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n208_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT80), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n207_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n205_), .A2(KEYINPUT80), .A3(new_n206_), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(KEYINPUT81), .B1(new_n221_), .B2(new_n215_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n215_), .A2(new_n220_), .A3(new_n219_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT81), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n202_), .B(new_n217_), .C1(new_n222_), .C2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G113gat), .B(G141gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G169gat), .B(G197gat), .ZN(new_n228_));
  XOR2_X1   g027(.A(new_n227_), .B(new_n228_), .Z(new_n229_));
  NOR2_X1   g028(.A1(new_n221_), .A2(new_n215_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n223_), .A2(new_n224_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n221_), .A2(KEYINPUT81), .A3(new_n215_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n230_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n226_), .B(new_n229_), .C1(new_n233_), .C2(new_n202_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT82), .ZN(new_n235_));
  OAI22_X1  g034(.A1(new_n222_), .A2(new_n225_), .B1(new_n215_), .B2(new_n221_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n202_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT82), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n238_), .A2(new_n239_), .A3(new_n226_), .A4(new_n229_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n235_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n238_), .A2(new_n226_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n229_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(G211gat), .B(G218gat), .Z(new_n247_));
  INV_X1    g046(.A(KEYINPUT21), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G197gat), .B(G204gat), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n249_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT21), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n251_), .A2(new_n247_), .A3(KEYINPUT21), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  AND2_X1   g054(.A1(KEYINPUT94), .A2(G233gat), .ZN(new_n256_));
  NOR2_X1   g055(.A1(KEYINPUT94), .A2(G233gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(G228gat), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT91), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT91), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n261_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G141gat), .A2(G148gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT2), .ZN(new_n265_));
  NOR3_X1   g064(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT90), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NOR4_X1   g067(.A1(KEYINPUT90), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n263_), .B(new_n265_), .C1(new_n268_), .C2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT92), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G155gat), .A2(G162gat), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT88), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(KEYINPUT88), .A2(G155gat), .A3(G162gat), .ZN(new_n275_));
  INV_X1    g074(.A(G155gat), .ZN(new_n276_));
  INV_X1    g075(.A(G162gat), .ZN(new_n277_));
  AOI22_X1  g076(.A1(new_n274_), .A2(new_n275_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n270_), .A2(new_n271_), .A3(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n271_), .B1(new_n270_), .B2(new_n278_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n275_), .ZN(new_n281_));
  AOI21_X1  g080(.A(KEYINPUT88), .B1(G155gat), .B2(G162gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT1), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT1), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n274_), .A2(new_n284_), .A3(new_n275_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n276_), .A2(new_n277_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n283_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  XOR2_X1   g086(.A(G141gat), .B(G148gat), .Z(new_n288_));
  AND3_X1   g087(.A1(new_n287_), .A2(KEYINPUT89), .A3(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(KEYINPUT89), .B1(new_n287_), .B2(new_n288_), .ZN(new_n290_));
  OAI22_X1  g089(.A1(new_n279_), .A2(new_n280_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT29), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n255_), .B(new_n258_), .C1(new_n292_), .C2(new_n293_), .ZN(new_n294_));
  XOR2_X1   g093(.A(new_n255_), .B(KEYINPUT95), .Z(new_n295_));
  AOI21_X1  g094(.A(new_n295_), .B1(KEYINPUT29), .B2(new_n291_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n294_), .B1(new_n296_), .B2(new_n258_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G78gat), .B(G106gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT96), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n291_), .A2(KEYINPUT29), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT93), .B(KEYINPUT28), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G22gat), .B(G50gat), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n302_), .B(new_n303_), .Z(new_n304_));
  XNOR2_X1  g103(.A(new_n301_), .B(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n300_), .A2(new_n305_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n297_), .A2(new_n298_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n299_), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n306_), .A2(new_n308_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G1gat), .B(G29gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(G85gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT0), .B(G57gat), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n313_), .B(new_n314_), .Z(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(G127gat), .B(G134gat), .Z(new_n317_));
  XOR2_X1   g116(.A(G113gat), .B(G120gat), .Z(new_n318_));
  XOR2_X1   g117(.A(new_n317_), .B(new_n318_), .Z(new_n319_));
  NAND2_X1  g118(.A1(new_n291_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n319_), .ZN(new_n321_));
  OAI221_X1 g120(.A(new_n321_), .B1(new_n289_), .B2(new_n290_), .C1(new_n279_), .C2(new_n280_), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G225gat), .A2(G233gat), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT4), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n291_), .A2(new_n328_), .A3(new_n319_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT103), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n320_), .A2(new_n322_), .A3(KEYINPUT4), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT102), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT102), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n320_), .A2(new_n322_), .A3(new_n333_), .A4(KEYINPUT4), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n330_), .B1(new_n332_), .B2(new_n334_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n316_), .B(new_n327_), .C1(new_n335_), .C2(new_n324_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n332_), .A2(new_n334_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT103), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n329_), .B(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n324_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n315_), .B1(new_n340_), .B2(new_n326_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n336_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G226gat), .A2(G233gat), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n343_), .B(new_n344_), .Z(new_n345_));
  INV_X1    g144(.A(G169gat), .ZN(new_n346_));
  INV_X1    g145(.A(G176gat), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT24), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT84), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n349_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT84), .B1(G169gat), .B2(G176gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  MUX2_X1   g151(.A(KEYINPUT24), .B(new_n348_), .S(new_n352_), .Z(new_n353_));
  NAND2_X1  g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT23), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT23), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n356_), .A2(G183gat), .A3(G190gat), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT25), .B(G183gat), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT26), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(G190gat), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(G190gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT26), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT83), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n358_), .B1(new_n362_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT85), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n358_), .A2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(G183gat), .A2(G190gat), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  OR2_X1    g169(.A1(new_n357_), .A2(new_n367_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n368_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(G169gat), .ZN(new_n374_));
  AOI22_X1  g173(.A1(new_n353_), .A2(new_n366_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n255_), .ZN(new_n376_));
  OAI211_X1 g175(.A(KEYINPUT20), .B(new_n345_), .C1(new_n375_), .C2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n361_), .A2(new_n364_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(new_n359_), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n368_), .A2(new_n371_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n353_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n355_), .A2(new_n357_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(new_n370_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n384_), .A2(KEYINPUT98), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(KEYINPUT98), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n374_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n376_), .A2(new_n382_), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT99), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n388_), .A2(new_n389_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n378_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT20), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n382_), .A2(new_n387_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n394_), .B1(new_n395_), .B2(new_n255_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n375_), .A2(new_n376_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n345_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  XOR2_X1   g199(.A(G8gat), .B(G36gat), .Z(new_n401_));
  XNOR2_X1  g200(.A(G64gat), .B(G92gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT32), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n393_), .A2(new_n400_), .A3(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n398_), .A2(new_n399_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n395_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n394_), .B1(new_n295_), .B2(new_n409_), .ZN(new_n410_));
  OR2_X1    g209(.A1(new_n410_), .A2(KEYINPUT105), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n295_), .A2(new_n409_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n412_), .A2(KEYINPUT105), .A3(KEYINPUT20), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n411_), .B(new_n413_), .C1(new_n376_), .C2(new_n375_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n408_), .B1(new_n414_), .B2(new_n399_), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n342_), .B(new_n407_), .C1(new_n415_), .C2(new_n406_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n405_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n409_), .A2(KEYINPUT99), .A3(new_n376_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n377_), .B1(new_n418_), .B2(new_n390_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n345_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n417_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n393_), .A2(new_n400_), .A3(new_n405_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT101), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  OAI211_X1 g223(.A(KEYINPUT101), .B(new_n417_), .C1(new_n419_), .C2(new_n420_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n337_), .A2(new_n324_), .A3(new_n339_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n315_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n426_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n341_), .A2(KEYINPUT33), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT33), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n432_), .B(new_n315_), .C1(new_n340_), .C2(new_n326_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n430_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT104), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n416_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  AOI211_X1 g235(.A(KEYINPUT104), .B(new_n430_), .C1(new_n431_), .C2(new_n433_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n311_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n311_), .A2(new_n342_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n422_), .A2(KEYINPUT27), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n414_), .A2(new_n399_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n408_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  XOR2_X1   g242(.A(new_n405_), .B(KEYINPUT106), .Z(new_n444_));
  AOI21_X1  g243(.A(new_n440_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT27), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n424_), .A2(new_n446_), .A3(new_n425_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT107), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  OR2_X1    g248(.A1(new_n447_), .A2(new_n448_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n445_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n439_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n438_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G227gat), .A2(G233gat), .ZN(new_n454_));
  INV_X1    g253(.A(G15gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n375_), .B(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT86), .B(KEYINPUT30), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(KEYINPUT87), .B1(new_n319_), .B2(KEYINPUT31), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n460_), .B1(KEYINPUT31), .B2(new_n319_), .ZN(new_n461_));
  XOR2_X1   g260(.A(new_n459_), .B(new_n461_), .Z(new_n462_));
  XNOR2_X1  g261(.A(G71gat), .B(G99gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(G43gat), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  OR2_X1    g264(.A1(new_n462_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n462_), .A2(new_n465_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n453_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n445_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n450_), .A2(new_n449_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n311_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n468_), .A2(new_n342_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n246_), .B1(new_n469_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(G99gat), .ZN(new_n478_));
  INV_X1    g277(.A(G106gat), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n478_), .A2(new_n479_), .A3(KEYINPUT67), .A4(KEYINPUT7), .ZN(new_n480_));
  NAND2_X1  g279(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n481_), .B1(G99gat), .B2(G106gat), .ZN(new_n482_));
  NOR2_X1   g281(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n480_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G99gat), .A2(G106gat), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT6), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT66), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT66), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT6), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n486_), .A2(new_n488_), .A3(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n489_), .A2(KEYINPUT6), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n487_), .A2(KEYINPUT66), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n485_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n484_), .A2(new_n491_), .A3(new_n494_), .ZN(new_n495_));
  AND2_X1   g294(.A1(G85gat), .A2(G92gat), .ZN(new_n496_));
  NOR2_X1   g295(.A1(G85gat), .A2(G92gat), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n495_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT8), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n495_), .A2(KEYINPUT8), .A3(new_n498_), .ZN(new_n502_));
  INV_X1    g301(.A(G92gat), .ZN(new_n503_));
  OAI22_X1  g302(.A1(new_n496_), .A2(new_n497_), .B1(KEYINPUT9), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(G85gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n503_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT9), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G85gat), .A2(G92gat), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n506_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n504_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT65), .ZN(new_n511_));
  INV_X1    g310(.A(new_n491_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n486_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT65), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n504_), .A2(new_n509_), .A3(new_n515_), .ZN(new_n516_));
  OR2_X1    g315(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n479_), .A2(KEYINPUT64), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT64), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(G106gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n517_), .A2(new_n518_), .A3(new_n520_), .A4(new_n521_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n511_), .A2(new_n514_), .A3(new_n516_), .A4(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G57gat), .B(G64gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G71gat), .B(G78gat), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n524_), .A2(new_n525_), .A3(KEYINPUT11), .ZN(new_n526_));
  INV_X1    g325(.A(new_n525_), .ZN(new_n527_));
  INV_X1    g326(.A(G64gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(G57gat), .ZN(new_n529_));
  INV_X1    g328(.A(G57gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(G64gat), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n529_), .A2(new_n531_), .A3(KEYINPUT11), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n527_), .A2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n524_), .A2(KEYINPUT11), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n526_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n501_), .A2(new_n502_), .A3(new_n523_), .A4(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT70), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G230gat), .A2(G233gat), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n537_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n501_), .A2(new_n502_), .A3(new_n523_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n535_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT12), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n535_), .A2(KEYINPUT69), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT69), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n548_), .B(new_n526_), .C1(new_n533_), .C2(new_n534_), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n547_), .A2(KEYINPUT12), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n542_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n546_), .A2(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(KEYINPUT71), .B1(new_n541_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n538_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n504_), .A2(new_n509_), .A3(new_n515_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n494_), .A2(new_n522_), .A3(new_n491_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  AOI22_X1  g356(.A1(new_n511_), .A2(new_n557_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n535_), .B1(new_n558_), .B2(new_n502_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n536_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n554_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT68), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  OAI211_X1 g362(.A(KEYINPUT68), .B(new_n554_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  AOI22_X1  g364(.A1(new_n544_), .A2(new_n545_), .B1(new_n542_), .B2(new_n550_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT71), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n566_), .B(new_n567_), .C1(new_n540_), .C2(new_n539_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n553_), .A2(new_n565_), .A3(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(G120gat), .B(G148gat), .Z(new_n570_));
  XNOR2_X1  g369(.A(G176gat), .B(G204gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n572_), .B(new_n573_), .Z(new_n574_));
  NAND2_X1  g373(.A1(new_n569_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n574_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n553_), .A2(new_n565_), .A3(new_n568_), .A4(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n575_), .A2(KEYINPUT73), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT73), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n569_), .A2(new_n579_), .A3(new_n574_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT13), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT74), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n583_), .A2(new_n584_), .ZN(new_n587_));
  NOR3_X1   g386(.A1(new_n586_), .A2(KEYINPUT75), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT75), .ZN(new_n589_));
  INV_X1    g388(.A(new_n583_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(KEYINPUT74), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n589_), .B1(new_n591_), .B2(new_n585_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n588_), .A2(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(G127gat), .B(G155gat), .Z(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT16), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G183gat), .B(G211gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT17), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n600_), .B(KEYINPUT79), .Z(new_n601_));
  XOR2_X1   g400(.A(new_n215_), .B(new_n601_), .Z(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n599_), .B1(new_n535_), .B2(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n604_), .B1(new_n535_), .B2(new_n603_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n547_), .A2(new_n549_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  AOI211_X1 g406(.A(new_n598_), .B(new_n597_), .C1(new_n602_), .C2(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n608_), .B1(new_n607_), .B2(new_n602_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n605_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n558_), .A2(new_n207_), .A3(new_n502_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n542_), .A2(new_n208_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(G232gat), .A2(G233gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT34), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n615_), .A2(KEYINPUT35), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n616_), .A2(KEYINPUT77), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n612_), .A2(new_n613_), .A3(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n615_), .A2(KEYINPUT35), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(G190gat), .B(G218gat), .Z(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT76), .ZN(new_n622_));
  XOR2_X1   g421(.A(G134gat), .B(G162gat), .Z(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT36), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n620_), .A2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n620_), .A2(new_n625_), .A3(new_n624_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT78), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n630_), .A2(KEYINPUT37), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(KEYINPUT37), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n629_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n627_), .A2(new_n630_), .A3(KEYINPUT37), .A4(new_n628_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  AND4_X1   g435(.A1(new_n477_), .A2(new_n593_), .A3(new_n611_), .A4(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n637_), .A2(new_n210_), .A3(new_n342_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(KEYINPUT108), .B(KEYINPUT38), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n639_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n629_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n642_), .B1(new_n469_), .B2(new_n476_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n586_), .A2(new_n587_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n644_), .A2(new_n246_), .A3(new_n610_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n643_), .A2(new_n645_), .A3(new_n342_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(G1gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n640_), .A2(new_n641_), .A3(new_n647_), .ZN(G1324gat));
  XNOR2_X1  g447(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n643_), .A2(new_n645_), .A3(new_n472_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(G8gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT39), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n637_), .A2(new_n211_), .A3(new_n472_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n649_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n651_), .A2(KEYINPUT39), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT39), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n656_), .B1(new_n650_), .B2(G8gat), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n653_), .B(new_n649_), .C1(new_n655_), .C2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n654_), .A2(new_n659_), .ZN(G1325gat));
  INV_X1    g459(.A(new_n468_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n637_), .A2(new_n455_), .A3(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n643_), .A2(new_n645_), .A3(new_n661_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n663_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT41), .B1(new_n663_), .B2(G15gat), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n662_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT110), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n666_), .B(new_n667_), .ZN(G1326gat));
  INV_X1    g467(.A(G22gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n637_), .A2(new_n669_), .A3(new_n473_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n643_), .A2(new_n645_), .A3(new_n473_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(G22gat), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n672_), .A2(KEYINPUT42), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n672_), .A2(KEYINPUT42), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n670_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT111), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n675_), .B(new_n676_), .ZN(G1327gat));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n635_), .B(KEYINPUT112), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n661_), .B1(new_n438_), .B2(new_n452_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n475_), .A2(new_n311_), .A3(new_n451_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n679_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n426_), .A2(new_n429_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n327_), .B1(new_n335_), .B2(new_n324_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n432_), .B1(new_n684_), .B2(new_n315_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n433_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n683_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT104), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n434_), .A2(new_n435_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n688_), .A2(new_n689_), .A3(new_n416_), .ZN(new_n690_));
  AOI22_X1  g489(.A1(new_n690_), .A2(new_n311_), .B1(new_n439_), .B2(new_n451_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n476_), .B1(new_n691_), .B2(new_n661_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n636_), .A2(KEYINPUT43), .ZN(new_n693_));
  AOI22_X1  g492(.A1(new_n682_), .A2(KEYINPUT43), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n644_), .A2(new_n246_), .A3(new_n611_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n678_), .B1(new_n694_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n692_), .B2(new_n679_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n693_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n700_), .B1(new_n469_), .B2(new_n476_), .ZN(new_n701_));
  OAI211_X1 g500(.A(KEYINPUT44), .B(new_n695_), .C1(new_n699_), .C2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n697_), .A2(new_n342_), .A3(new_n702_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n703_), .A2(KEYINPUT113), .ZN(new_n704_));
  OAI21_X1  g503(.A(G29gat), .B1(new_n703_), .B2(KEYINPUT113), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n629_), .A2(new_n611_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n644_), .A2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n477_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n342_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n710_), .A2(G29gat), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT114), .Z(new_n712_));
  OAI22_X1  g511(.A1(new_n704_), .A2(new_n705_), .B1(new_n709_), .B2(new_n712_), .ZN(G1328gat));
  NAND3_X1  g512(.A1(new_n697_), .A2(new_n472_), .A3(new_n702_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(G36gat), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n451_), .A2(G36gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n477_), .A2(new_n708_), .A3(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT45), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n715_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT46), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n715_), .A2(KEYINPUT46), .A3(new_n718_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1329gat));
  NOR3_X1   g522(.A1(new_n709_), .A2(G43gat), .A3(new_n468_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n697_), .A2(new_n661_), .A3(new_n702_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n725_), .B2(G43gat), .ZN(new_n726_));
  XNOR2_X1  g525(.A(KEYINPUT115), .B(KEYINPUT47), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n726_), .B(new_n728_), .ZN(G1330gat));
  NAND4_X1  g528(.A1(new_n697_), .A2(G50gat), .A3(new_n702_), .A4(new_n473_), .ZN(new_n730_));
  INV_X1    g529(.A(G50gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n731_), .B1(new_n709_), .B2(new_n311_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n730_), .A2(new_n732_), .ZN(G1331gat));
  AOI21_X1  g532(.A(new_n245_), .B1(new_n469_), .B2(new_n476_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n734_), .A2(KEYINPUT116), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n734_), .A2(KEYINPUT116), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n644_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n738_), .A2(new_n610_), .A3(new_n635_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n740_), .A2(G57gat), .A3(new_n710_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n593_), .ZN(new_n742_));
  AND4_X1   g541(.A1(new_n246_), .A2(new_n643_), .A3(new_n742_), .A4(new_n611_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n530_), .B1(new_n743_), .B2(new_n342_), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n741_), .A2(new_n744_), .ZN(G1332gat));
  INV_X1    g544(.A(KEYINPUT48), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n743_), .A2(new_n472_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n747_), .B2(G64gat), .ZN(new_n748_));
  AOI211_X1 g547(.A(KEYINPUT48), .B(new_n528_), .C1(new_n743_), .C2(new_n472_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n472_), .A2(new_n528_), .ZN(new_n750_));
  OAI22_X1  g549(.A1(new_n748_), .A2(new_n749_), .B1(new_n740_), .B2(new_n750_), .ZN(G1333gat));
  INV_X1    g550(.A(KEYINPUT49), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n743_), .A2(new_n661_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n753_), .B2(G71gat), .ZN(new_n754_));
  INV_X1    g553(.A(G71gat), .ZN(new_n755_));
  AOI211_X1 g554(.A(KEYINPUT49), .B(new_n755_), .C1(new_n743_), .C2(new_n661_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n661_), .A2(new_n755_), .ZN(new_n757_));
  OAI22_X1  g556(.A1(new_n754_), .A2(new_n756_), .B1(new_n740_), .B2(new_n757_), .ZN(G1334gat));
  INV_X1    g557(.A(KEYINPUT50), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n743_), .A2(new_n473_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n760_), .B2(G78gat), .ZN(new_n761_));
  INV_X1    g560(.A(G78gat), .ZN(new_n762_));
  AOI211_X1 g561(.A(KEYINPUT50), .B(new_n762_), .C1(new_n743_), .C2(new_n473_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n473_), .A2(new_n762_), .ZN(new_n764_));
  OAI22_X1  g563(.A1(new_n761_), .A2(new_n763_), .B1(new_n740_), .B2(new_n764_), .ZN(G1335gat));
  NOR2_X1   g564(.A1(new_n593_), .A2(new_n707_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n737_), .A2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n767_), .A2(new_n505_), .A3(new_n342_), .ZN(new_n768_));
  NOR4_X1   g567(.A1(new_n694_), .A2(new_n245_), .A3(new_n738_), .A4(new_n611_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n342_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n768_), .B1(new_n505_), .B2(new_n771_), .ZN(G1336gat));
  NAND3_X1  g571(.A1(new_n767_), .A2(new_n503_), .A3(new_n472_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n769_), .A2(new_n472_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n773_), .B1(new_n503_), .B2(new_n775_), .ZN(G1337gat));
  INV_X1    g575(.A(KEYINPUT117), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n777_), .A2(KEYINPUT51), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n738_), .A2(new_n245_), .A3(new_n611_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n779_), .B(new_n661_), .C1(new_n699_), .C2(new_n701_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(G99gat), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n661_), .A2(new_n517_), .A3(new_n521_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n766_), .B(new_n782_), .C1(new_n735_), .C2(new_n736_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n778_), .B1(new_n781_), .B2(new_n783_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n777_), .A2(KEYINPUT51), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n784_), .B(new_n785_), .ZN(G1338gat));
  AND3_X1   g585(.A1(new_n473_), .A2(new_n518_), .A3(new_n520_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n737_), .A2(new_n766_), .A3(new_n787_), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n779_), .B(new_n473_), .C1(new_n699_), .C2(new_n701_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n789_), .A2(new_n790_), .A3(G106gat), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n789_), .B2(G106gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n788_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT53), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n788_), .B(new_n795_), .C1(new_n792_), .C2(new_n791_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(G1339gat));
  INV_X1    g596(.A(KEYINPUT122), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n474_), .A2(new_n342_), .A3(new_n661_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n217_), .B1(new_n222_), .B2(new_n225_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n202_), .B1(new_n800_), .B2(KEYINPUT119), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n801_), .B1(KEYINPUT119), .B2(new_n800_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n229_), .B1(new_n236_), .B2(new_n202_), .ZN(new_n803_));
  AOI22_X1  g602(.A1(new_n235_), .A2(new_n240_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n578_), .A2(new_n580_), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT120), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT120), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n578_), .A2(new_n807_), .A3(new_n580_), .A4(new_n804_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n245_), .A2(new_n577_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n553_), .A2(new_n811_), .A3(new_n568_), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n566_), .B(KEYINPUT55), .C1(new_n540_), .C2(new_n539_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n546_), .A2(new_n551_), .A3(new_n536_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n554_), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n813_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n812_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n574_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT56), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n817_), .A2(KEYINPUT56), .A3(new_n574_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n810_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n809_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n629_), .A2(KEYINPUT57), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n824_), .A2(KEYINPUT121), .A3(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT121), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n822_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(new_n825_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n827_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n820_), .A2(new_n821_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n804_), .A2(new_n577_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT58), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n832_), .A2(KEYINPUT58), .A3(new_n833_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(new_n635_), .A3(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n642_), .B1(new_n809_), .B2(new_n823_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n839_), .B2(KEYINPUT57), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n610_), .B1(new_n831_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n246_), .B2(new_n611_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n245_), .A2(KEYINPUT118), .A3(new_n610_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n635_), .A2(new_n843_), .A3(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n583_), .A2(new_n845_), .A3(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n846_), .B1(new_n583_), .B2(new_n845_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n799_), .B1(new_n841_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n798_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n829_), .B2(new_n642_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n827_), .A2(new_n856_), .A3(new_n830_), .A4(new_n838_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n850_), .B1(new_n857_), .B2(new_n610_), .ZN(new_n858_));
  OAI211_X1 g657(.A(KEYINPUT122), .B(KEYINPUT59), .C1(new_n858_), .C2(new_n799_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n854_), .A2(new_n859_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n857_), .A2(KEYINPUT123), .A3(new_n610_), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT123), .B1(new_n857_), .B2(new_n610_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n851_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n799_), .A2(KEYINPUT59), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n860_), .A2(new_n245_), .A3(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(G113gat), .ZN(new_n867_));
  INV_X1    g666(.A(new_n852_), .ZN(new_n868_));
  OR2_X1    g667(.A1(new_n246_), .A2(G113gat), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n867_), .B1(new_n868_), .B2(new_n869_), .ZN(G1340gat));
  AOI21_X1  g669(.A(new_n593_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n860_), .A2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT124), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n860_), .A2(new_n871_), .A3(KEYINPUT124), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n874_), .A2(G120gat), .A3(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(G120gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(new_n738_), .B2(KEYINPUT60), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n852_), .B(new_n878_), .C1(KEYINPUT60), .C2(new_n877_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n876_), .A2(new_n879_), .ZN(G1341gat));
  NAND3_X1  g679(.A1(new_n860_), .A2(new_n611_), .A3(new_n865_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(G127gat), .ZN(new_n882_));
  OR2_X1    g681(.A1(new_n610_), .A2(G127gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n868_), .B2(new_n883_), .ZN(G1342gat));
  NAND3_X1  g683(.A1(new_n860_), .A2(new_n635_), .A3(new_n865_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(G134gat), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n629_), .A2(G134gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n868_), .B2(new_n887_), .ZN(G1343gat));
  NOR2_X1   g687(.A1(new_n858_), .A2(new_n661_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n472_), .A2(new_n311_), .A3(new_n710_), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n889_), .A2(KEYINPUT125), .A3(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(KEYINPUT125), .B1(new_n889_), .B2(new_n890_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n245_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G141gat), .ZN(G1344gat));
  OAI21_X1  g693(.A(new_n742_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G148gat), .ZN(G1345gat));
  OAI21_X1  g695(.A(new_n611_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT61), .B(G155gat), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n897_), .B(new_n898_), .ZN(G1346gat));
  OR2_X1    g698(.A1(new_n891_), .A2(new_n892_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n642_), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n679_), .A2(G162gat), .ZN(new_n902_));
  AOI22_X1  g701(.A1(new_n901_), .A2(new_n277_), .B1(new_n900_), .B2(new_n902_), .ZN(G1347gat));
  NAND2_X1  g702(.A1(new_n475_), .A2(new_n472_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n863_), .A2(new_n245_), .A3(new_n311_), .A4(new_n905_), .ZN(new_n906_));
  OAI211_X1 g705(.A(KEYINPUT62), .B(new_n346_), .C1(new_n906_), .C2(KEYINPUT22), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(KEYINPUT62), .B1(new_n906_), .B2(KEYINPUT22), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n906_), .A2(KEYINPUT62), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n910_), .A2(new_n346_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n908_), .B1(new_n909_), .B2(new_n911_), .ZN(G1348gat));
  AND2_X1   g711(.A1(new_n863_), .A2(new_n311_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n913_), .A2(new_n644_), .A3(new_n905_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n858_), .A2(new_n473_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n593_), .A2(new_n347_), .A3(new_n904_), .ZN(new_n916_));
  AOI22_X1  g715(.A1(new_n914_), .A2(new_n347_), .B1(new_n915_), .B2(new_n916_), .ZN(G1349gat));
  NOR2_X1   g716(.A1(new_n904_), .A2(new_n610_), .ZN(new_n918_));
  AOI21_X1  g717(.A(G183gat), .B1(new_n915_), .B2(new_n918_), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n904_), .A2(new_n359_), .A3(new_n610_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n919_), .B1(new_n913_), .B2(new_n920_), .ZN(G1350gat));
  NAND2_X1  g720(.A1(new_n913_), .A2(new_n905_), .ZN(new_n922_));
  OAI21_X1  g721(.A(G190gat), .B1(new_n922_), .B2(new_n636_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n642_), .A2(new_n379_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n922_), .B2(new_n924_), .ZN(G1351gat));
  AND3_X1   g724(.A1(new_n889_), .A2(new_n439_), .A3(new_n472_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n245_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(G197gat), .ZN(G1352gat));
  AND2_X1   g727(.A1(new_n926_), .A2(new_n742_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT126), .ZN(new_n930_));
  AND2_X1   g729(.A1(new_n930_), .A2(G204gat), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n930_), .A2(G204gat), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n929_), .B1(new_n931_), .B2(new_n932_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n933_), .B1(new_n929_), .B2(new_n932_), .ZN(G1353gat));
  NAND2_X1  g733(.A1(new_n926_), .A2(new_n611_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(KEYINPUT63), .B(G211gat), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n937_), .B1(new_n935_), .B2(new_n938_), .ZN(G1354gat));
  NAND2_X1  g738(.A1(new_n926_), .A2(new_n642_), .ZN(new_n940_));
  XOR2_X1   g739(.A(KEYINPUT127), .B(G218gat), .Z(new_n941_));
  NOR2_X1   g740(.A1(new_n636_), .A2(new_n941_), .ZN(new_n942_));
  AOI22_X1  g741(.A1(new_n940_), .A2(new_n941_), .B1(new_n926_), .B2(new_n942_), .ZN(G1355gat));
endmodule


