//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n824_, new_n825_,
    new_n826_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n841_, new_n843_, new_n844_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n881_,
    new_n883_, new_n884_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT82), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT82), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n206_), .B1(new_n202_), .B2(new_n203_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(new_n208_), .B(KEYINPUT31), .Z(new_n209_));
  INV_X1    g008(.A(G99gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT79), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(KEYINPUT24), .A3(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n212_), .B(KEYINPUT79), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT24), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT23), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT25), .B(G183gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT78), .ZN(new_n223_));
  INV_X1    g022(.A(G190gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT26), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n224_), .A2(KEYINPUT26), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n222_), .B(new_n225_), .C1(new_n226_), .C2(new_n223_), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n216_), .A2(new_n219_), .A3(new_n221_), .A4(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n221_), .B1(G183gat), .B2(G190gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n230_));
  OR3_X1    g029(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n229_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n228_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT80), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT80), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n228_), .A2(new_n235_), .A3(new_n232_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G15gat), .B(G43gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT81), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT30), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n237_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n234_), .A2(new_n236_), .A3(new_n240_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G227gat), .A2(G233gat), .ZN(new_n244_));
  INV_X1    g043(.A(G71gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n242_), .A2(new_n243_), .A3(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n247_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n249_));
  OR3_X1    g048(.A1(new_n211_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n211_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G1gat), .B(G29gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(G85gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT0), .B(G57gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G155gat), .A2(G162gat), .ZN(new_n258_));
  OR2_X1    g057(.A1(G155gat), .A2(G162gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT3), .ZN(new_n260_));
  INV_X1    g059(.A(G141gat), .ZN(new_n261_));
  INV_X1    g060(.A(G148gat), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G141gat), .A2(G148gat), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT84), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n263_), .B(new_n264_), .C1(new_n267_), .C2(KEYINPUT2), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n267_), .A2(KEYINPUT2), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n258_), .B(new_n259_), .C1(new_n268_), .C2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n261_), .A2(new_n262_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT83), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n272_), .B1(new_n258_), .B2(KEYINPUT1), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n258_), .A2(KEYINPUT1), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(new_n274_), .A3(new_n259_), .ZN(new_n275_));
  NOR3_X1   g074(.A1(new_n258_), .A2(new_n272_), .A3(KEYINPUT1), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n265_), .B(new_n271_), .C1(new_n275_), .C2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n270_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n278_), .A2(new_n205_), .A3(new_n207_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n270_), .A2(new_n277_), .A3(new_n204_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT4), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n279_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G225gat), .A2(G233gat), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n281_), .A2(new_n286_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n257_), .B1(new_n287_), .B2(new_n289_), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n256_), .B(new_n288_), .C1(new_n285_), .C2(new_n286_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT90), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G78gat), .B(G106gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT86), .B(G204gat), .ZN(new_n295_));
  INV_X1    g094(.A(G197gat), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT87), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT87), .B1(new_n296_), .B2(G204gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n299_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G211gat), .B(G218gat), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT21), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n298_), .A2(new_n300_), .A3(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(KEYINPUT21), .B1(new_n298_), .B2(new_n300_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n302_), .B1(G197gat), .B2(G204gat), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n306_), .B1(new_n295_), .B2(G197gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n301_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n304_), .B1(new_n305_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G228gat), .A2(G233gat), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n278_), .A2(KEYINPUT29), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n312_), .A2(KEYINPUT85), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(KEYINPUT85), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n311_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT88), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n311_), .A2(new_n313_), .A3(KEYINPUT88), .A4(new_n314_), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n310_), .B1(new_n309_), .B2(new_n312_), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n293_), .B(new_n294_), .C1(new_n319_), .C2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n320_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n294_), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT90), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n278_), .A2(KEYINPUT29), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT28), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G22gat), .B(G50gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n294_), .B(KEYINPUT89), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n328_), .B1(new_n322_), .B2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n321_), .A2(new_n324_), .A3(new_n330_), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n322_), .A2(new_n329_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n322_), .A2(new_n329_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n328_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n292_), .B1(new_n331_), .B2(new_n334_), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n305_), .A2(new_n308_), .ZN(new_n336_));
  AOI22_X1  g135(.A1(new_n234_), .A2(new_n236_), .B1(new_n336_), .B2(new_n304_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G226gat), .A2(G233gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT26), .B(G190gat), .ZN(new_n342_));
  AOI22_X1  g141(.A1(new_n222_), .A2(new_n342_), .B1(new_n218_), .B2(new_n212_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n216_), .A2(new_n221_), .A3(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT22), .B(G169gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT92), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n346_), .A2(G176gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n229_), .A2(new_n215_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n344_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  OAI211_X1 g148(.A(KEYINPUT20), .B(new_n341_), .C1(new_n349_), .C2(new_n309_), .ZN(new_n350_));
  OR3_X1    g149(.A1(new_n337_), .A2(new_n350_), .A3(KEYINPUT93), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n309_), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n352_), .B(KEYINPUT20), .C1(new_n237_), .C2(new_n309_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(new_n340_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT93), .B1(new_n337_), .B2(new_n350_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n351_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G8gat), .B(G36gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT18), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G64gat), .B(G92gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n358_), .B(new_n359_), .Z(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n356_), .A2(new_n361_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n351_), .A2(new_n354_), .A3(new_n360_), .A4(new_n355_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT95), .B(KEYINPUT27), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n363_), .A2(KEYINPUT27), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT94), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT20), .B1(new_n349_), .B2(new_n309_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n337_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n368_), .A2(new_n367_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n341_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n353_), .A2(new_n340_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n361_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n364_), .A2(new_n365_), .B1(new_n366_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n335_), .A2(new_n374_), .ZN(new_n375_));
  AOI22_X1  g174(.A1(new_n282_), .A2(new_n284_), .B1(G225gat), .B2(G233gat), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n256_), .B1(new_n281_), .B2(new_n286_), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT33), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n290_), .A2(new_n378_), .ZN(new_n379_));
  OAI211_X1 g178(.A(KEYINPUT33), .B(new_n257_), .C1(new_n287_), .C2(new_n289_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n362_), .A2(new_n379_), .A3(new_n363_), .A4(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n371_), .A2(new_n372_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n360_), .A2(KEYINPUT32), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n292_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n356_), .B1(KEYINPUT32), .B2(new_n360_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n381_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(new_n334_), .A3(new_n331_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n252_), .B1(new_n375_), .B2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n292_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n389_), .A2(new_n334_), .A3(new_n331_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT96), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n364_), .A2(new_n365_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n366_), .A2(new_n373_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n391_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n374_), .A2(new_n391_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n390_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n388_), .A2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G15gat), .B(G22gat), .ZN(new_n399_));
  INV_X1    g198(.A(G1gat), .ZN(new_n400_));
  INV_X1    g199(.A(G8gat), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT14), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n399_), .A2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G1gat), .B(G8gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G29gat), .B(G36gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G43gat), .B(G50gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n405_), .B(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n410_), .A2(G229gat), .A3(G233gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n408_), .B(KEYINPUT15), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n405_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G229gat), .A2(G233gat), .ZN(new_n414_));
  XOR2_X1   g213(.A(new_n414_), .B(KEYINPUT76), .Z(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n405_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n416_), .B1(new_n417_), .B2(new_n408_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n413_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n411_), .A2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G113gat), .B(G141gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G169gat), .B(G197gat), .ZN(new_n422_));
  XOR2_X1   g221(.A(new_n421_), .B(new_n422_), .Z(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n420_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT77), .ZN(new_n426_));
  INV_X1    g225(.A(new_n420_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n426_), .B1(new_n427_), .B2(new_n423_), .ZN(new_n428_));
  NOR3_X1   g227(.A1(new_n420_), .A2(KEYINPUT77), .A3(new_n424_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n425_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n398_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G57gat), .B(G64gat), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n433_), .A2(KEYINPUT11), .ZN(new_n434_));
  INV_X1    g233(.A(G64gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(G57gat), .ZN(new_n436_));
  INV_X1    g235(.A(G57gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(G64gat), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n438_), .A3(KEYINPUT11), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT67), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT67), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n433_), .A2(new_n441_), .A3(KEYINPUT11), .ZN(new_n442_));
  XOR2_X1   g241(.A(G71gat), .B(G78gat), .Z(new_n443_));
  NAND4_X1  g242(.A1(new_n434_), .A2(new_n440_), .A3(new_n442_), .A4(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n443_), .B1(KEYINPUT11), .B2(new_n433_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n439_), .A2(KEYINPUT67), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n441_), .B1(new_n433_), .B2(KEYINPUT11), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n445_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n444_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT68), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n444_), .A2(new_n448_), .A3(KEYINPUT68), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G231gat), .A2(G233gat), .ZN(new_n454_));
  XOR2_X1   g253(.A(new_n454_), .B(KEYINPUT75), .Z(new_n455_));
  XNOR2_X1  g254(.A(new_n405_), .B(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n453_), .B(new_n456_), .ZN(new_n457_));
  XOR2_X1   g256(.A(G127gat), .B(G155gat), .Z(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT16), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G183gat), .B(G211gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT17), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n461_), .A2(new_n462_), .ZN(new_n464_));
  NOR3_X1   g263(.A1(new_n457_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n456_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n463_), .B1(new_n466_), .B2(new_n449_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n467_), .B1(new_n449_), .B2(new_n466_), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n465_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT37), .ZN(new_n470_));
  INV_X1    g269(.A(G85gat), .ZN(new_n471_));
  INV_X1    g270(.A(G92gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G85gat), .A2(G92gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT9), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n474_), .A2(KEYINPUT9), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G99gat), .A2(G106gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT6), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT6), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(G99gat), .A3(G106gat), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n478_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT10), .B(G99gat), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n484_), .A2(G106gat), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT64), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NOR3_X1   g286(.A1(new_n484_), .A2(KEYINPUT64), .A3(G106gat), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n477_), .B(new_n483_), .C1(new_n487_), .C2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT65), .ZN(new_n490_));
  INV_X1    g289(.A(G106gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n210_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT7), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n480_), .A2(new_n482_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT7), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n490_), .A2(new_n495_), .A3(new_n210_), .A4(new_n491_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n493_), .A2(new_n494_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT8), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT66), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n498_), .B1(new_n475_), .B2(new_n499_), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n497_), .A2(new_n476_), .A3(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n500_), .B1(new_n497_), .B2(new_n476_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT69), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n501_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n497_), .A2(new_n476_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n500_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n497_), .A2(new_n500_), .A3(new_n476_), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT69), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n489_), .B1(new_n504_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(new_n412_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G232gat), .A2(G233gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT34), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT35), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n489_), .A2(new_n508_), .A3(new_n507_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n511_), .B(new_n516_), .C1(new_n409_), .C2(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n514_), .A2(new_n515_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT74), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n518_), .A2(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n520_), .A2(new_n521_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n524_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n518_), .A2(new_n526_), .A3(new_n522_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G190gat), .B(G218gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G134gat), .B(G162gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n530_), .B(KEYINPUT36), .Z(new_n531_));
  NAND3_X1  g330(.A1(new_n525_), .A2(new_n527_), .A3(new_n531_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n525_), .A2(new_n527_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n530_), .A2(KEYINPUT36), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n470_), .B(new_n532_), .C1(new_n533_), .C2(new_n535_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n525_), .A2(new_n527_), .A3(new_n531_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n535_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT37), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n469_), .B1(new_n536_), .B2(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n501_), .A2(new_n502_), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n444_), .A2(new_n448_), .A3(KEYINPUT68), .ZN(new_n542_));
  AOI21_X1  g341(.A(KEYINPUT68), .B1(new_n444_), .B2(new_n448_), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n541_), .B(new_n489_), .C1(new_n542_), .C2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n517_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G230gat), .A2(G233gat), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT71), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n544_), .A2(new_n550_), .A3(new_n547_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n550_), .B1(new_n544_), .B2(new_n547_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT12), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n449_), .A2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n510_), .A2(KEYINPUT70), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT70), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n477_), .A2(new_n483_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n487_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n488_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n558_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n503_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n507_), .A2(KEYINPUT69), .A3(new_n508_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n561_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n555_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n557_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n545_), .A2(new_n554_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n556_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n549_), .B1(new_n553_), .B2(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(G120gat), .B(G148gat), .Z(new_n570_));
  XNOR2_X1  g369(.A(G176gat), .B(G204gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n572_), .B(new_n573_), .Z(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n569_), .A2(new_n575_), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n549_), .B(new_n574_), .C1(new_n553_), .C2(new_n568_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n578_), .B1(KEYINPUT73), .B2(KEYINPUT13), .ZN(new_n579_));
  XOR2_X1   g378(.A(KEYINPUT73), .B(KEYINPUT13), .Z(new_n580_));
  OAI21_X1  g379(.A(new_n579_), .B1(new_n578_), .B2(new_n580_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n540_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n432_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT97), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT97), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n432_), .A2(new_n585_), .A3(new_n582_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n584_), .A2(new_n400_), .A3(new_n292_), .A4(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT38), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n537_), .A2(new_n538_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT98), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n398_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n581_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n593_), .A2(new_n431_), .A3(new_n469_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n292_), .ZN(new_n596_));
  OAI21_X1  g395(.A(G1gat), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n587_), .A2(new_n588_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n589_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT99), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n589_), .A2(KEYINPUT99), .A3(new_n597_), .A4(new_n598_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(G1324gat));
  XNOR2_X1  g402(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT39), .ZN(new_n605_));
  INV_X1    g404(.A(new_n595_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n392_), .A2(new_n393_), .A3(new_n391_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n607_), .A2(new_n394_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n605_), .B1(new_n609_), .B2(G8gat), .ZN(new_n610_));
  AOI211_X1 g409(.A(KEYINPUT39), .B(new_n401_), .C1(new_n606_), .C2(new_n608_), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n584_), .A2(new_n401_), .A3(new_n608_), .A4(new_n586_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n604_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  OAI211_X1 g413(.A(new_n613_), .B(new_n604_), .C1(new_n610_), .C2(new_n611_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n614_), .A2(new_n616_), .ZN(G1325gat));
  INV_X1    g416(.A(new_n252_), .ZN(new_n618_));
  OAI21_X1  g417(.A(G15gat), .B1(new_n595_), .B2(new_n618_), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n619_), .A2(KEYINPUT101), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(KEYINPUT101), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n620_), .A2(KEYINPUT41), .A3(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(KEYINPUT41), .B1(new_n620_), .B2(new_n621_), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n583_), .A2(G15gat), .A3(new_n618_), .ZN(new_n624_));
  OR3_X1    g423(.A1(new_n622_), .A2(new_n623_), .A3(new_n624_), .ZN(G1326gat));
  INV_X1    g424(.A(KEYINPUT42), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n331_), .A2(new_n334_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT102), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n606_), .A2(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n626_), .B1(new_n629_), .B2(G22gat), .ZN(new_n630_));
  INV_X1    g429(.A(G22gat), .ZN(new_n631_));
  AOI211_X1 g430(.A(KEYINPUT42), .B(new_n631_), .C1(new_n606_), .C2(new_n628_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n628_), .A2(new_n631_), .ZN(new_n633_));
  OAI22_X1  g432(.A1(new_n630_), .A2(new_n632_), .B1(new_n583_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT103), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(G1327gat));
  NAND3_X1  g435(.A1(new_n581_), .A2(new_n430_), .A3(new_n469_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n637_), .B(KEYINPUT104), .Z(new_n638_));
  AND2_X1   g437(.A1(new_n536_), .A2(new_n539_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n639_), .B1(new_n388_), .B2(new_n397_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT105), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n640_), .A2(new_n641_), .A3(KEYINPUT43), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT43), .B1(new_n640_), .B2(new_n641_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n638_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT44), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  OAI211_X1 g445(.A(new_n638_), .B(KEYINPUT44), .C1(new_n642_), .C2(new_n643_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n646_), .A2(new_n292_), .A3(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(G29gat), .ZN(new_n649_));
  INV_X1    g448(.A(new_n469_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n590_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n593_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n432_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n596_), .A2(G29gat), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT106), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n649_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(KEYINPUT107), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT107), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n649_), .A2(new_n660_), .A3(new_n657_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n661_), .ZN(G1328gat));
  NAND3_X1  g461(.A1(new_n646_), .A2(new_n608_), .A3(new_n647_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(G36gat), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n608_), .B(KEYINPUT108), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n653_), .A2(G36gat), .A3(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT45), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n666_), .B(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n664_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT46), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n664_), .A2(new_n668_), .A3(KEYINPUT46), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1329gat));
  NAND4_X1  g472(.A1(new_n646_), .A2(G43gat), .A3(new_n252_), .A4(new_n647_), .ZN(new_n674_));
  INV_X1    g473(.A(G43gat), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n675_), .B1(new_n653_), .B2(new_n618_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g477(.A(G50gat), .B1(new_n654_), .B2(new_n628_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n646_), .A2(new_n647_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n627_), .A2(G50gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n679_), .B1(new_n680_), .B2(new_n681_), .ZN(G1331gat));
  NOR2_X1   g481(.A1(new_n398_), .A2(new_n430_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n639_), .A2(new_n581_), .A3(new_n469_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n685_), .A2(KEYINPUT109), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n596_), .B1(new_n685_), .B2(KEYINPUT109), .ZN(new_n687_));
  AOI21_X1  g486(.A(G57gat), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n688_), .A2(KEYINPUT110), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(KEYINPUT110), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n581_), .A2(new_n430_), .A3(new_n469_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n591_), .ZN(new_n692_));
  OAI211_X1 g491(.A(new_n691_), .B(new_n692_), .C1(new_n388_), .C2(new_n397_), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n693_), .A2(KEYINPUT111), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(KEYINPUT111), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n596_), .A2(new_n437_), .ZN(new_n697_));
  AOI22_X1  g496(.A1(new_n689_), .A2(new_n690_), .B1(new_n696_), .B2(new_n697_), .ZN(G1332gat));
  INV_X1    g497(.A(new_n685_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n665_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(new_n435_), .A3(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n694_), .A2(new_n700_), .A3(new_n695_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n702_), .A2(G64gat), .A3(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n702_), .B2(G64gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n701_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT113), .ZN(G1333gat));
  NAND3_X1  g506(.A1(new_n699_), .A2(new_n245_), .A3(new_n252_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n696_), .A2(new_n252_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(G71gat), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n710_), .A2(KEYINPUT49), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(KEYINPUT49), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n708_), .B1(new_n711_), .B2(new_n712_), .ZN(G1334gat));
  INV_X1    g512(.A(new_n628_), .ZN(new_n714_));
  OR3_X1    g513(.A1(new_n685_), .A2(G78gat), .A3(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n696_), .A2(new_n628_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(G78gat), .ZN(new_n717_));
  XOR2_X1   g516(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n718_));
  AND2_X1   g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n717_), .A2(new_n718_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n715_), .B1(new_n719_), .B2(new_n720_), .ZN(G1335gat));
  NAND4_X1  g520(.A1(new_n683_), .A2(new_n593_), .A3(new_n469_), .A4(new_n590_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n723_), .A2(new_n471_), .A3(new_n292_), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n642_), .A2(new_n643_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n581_), .A2(new_n430_), .A3(new_n650_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n292_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n724_), .B1(new_n730_), .B2(new_n471_), .ZN(G1336gat));
  NAND3_X1  g530(.A1(new_n723_), .A2(new_n472_), .A3(new_n608_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n728_), .A2(new_n700_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n732_), .B1(new_n734_), .B2(new_n472_), .ZN(G1337gat));
  OAI21_X1  g534(.A(G99gat), .B1(new_n727_), .B2(new_n618_), .ZN(new_n736_));
  OR3_X1    g535(.A1(new_n722_), .A2(new_n618_), .A3(new_n484_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  AND2_X1   g537(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n738_), .B(new_n739_), .ZN(G1338gat));
  NAND3_X1  g539(.A1(new_n723_), .A2(new_n491_), .A3(new_n627_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT116), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n627_), .B(new_n726_), .C1(new_n642_), .C2(new_n643_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT52), .ZN(new_n744_));
  AND4_X1   g543(.A1(new_n742_), .A2(new_n743_), .A3(new_n744_), .A4(G106gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n491_), .B1(KEYINPUT116), .B2(KEYINPUT52), .ZN(new_n746_));
  AOI22_X1  g545(.A1(new_n743_), .A2(new_n746_), .B1(new_n742_), .B2(new_n744_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n741_), .B1(new_n745_), .B2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT53), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT53), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n750_), .B(new_n741_), .C1(new_n745_), .C2(new_n747_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(G1339gat));
  NAND3_X1  g551(.A1(new_n540_), .A2(new_n581_), .A3(new_n431_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT54), .Z(new_n754_));
  NAND2_X1  g553(.A1(new_n430_), .A2(new_n577_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT117), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT117), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n430_), .A2(new_n577_), .A3(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n556_), .A2(new_n566_), .A3(new_n544_), .A4(new_n567_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n548_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT118), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT118), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n760_), .A2(new_n763_), .A3(new_n548_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n765_), .B1(new_n553_), .B2(new_n568_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n544_), .A2(new_n547_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT71), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n544_), .A2(new_n550_), .A3(new_n547_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n564_), .A2(new_n565_), .ZN(new_n771_));
  AOI22_X1  g570(.A1(new_n771_), .A2(KEYINPUT70), .B1(new_n554_), .B2(new_n545_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n770_), .A2(new_n772_), .A3(KEYINPUT55), .A4(new_n566_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n762_), .A2(new_n764_), .A3(new_n766_), .A4(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n575_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT56), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n774_), .A2(KEYINPUT56), .A3(new_n575_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n759_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n428_), .A2(new_n429_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n413_), .B(new_n416_), .C1(new_n405_), .C2(new_n409_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n423_), .B1(new_n410_), .B2(new_n415_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n780_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n578_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n651_), .B1(new_n779_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT57), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n774_), .A2(KEYINPUT56), .A3(new_n575_), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT56), .B1(new_n774_), .B2(new_n575_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n756_), .B(new_n758_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n784_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n792_), .A2(KEYINPUT57), .A3(new_n651_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT119), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n783_), .A2(new_n577_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n794_), .B(new_n639_), .C1(new_n796_), .C2(KEYINPUT58), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(KEYINPUT58), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n783_), .A2(new_n577_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n800_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT58), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n794_), .B1(new_n803_), .B2(new_n639_), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n788_), .B(new_n793_), .C1(new_n799_), .C2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n754_), .B1(new_n805_), .B2(new_n469_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n806_), .A2(new_n627_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n608_), .A2(new_n596_), .A3(new_n618_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT59), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n807_), .A2(KEYINPUT59), .A3(new_n808_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n431_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(G113gat), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n430_), .A2(new_n814_), .ZN(new_n815_));
  OAI22_X1  g614(.A1(new_n813_), .A2(new_n814_), .B1(new_n809_), .B2(new_n815_), .ZN(G1340gat));
  AOI21_X1  g615(.A(new_n581_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n817_));
  INV_X1    g616(.A(G120gat), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n818_), .B1(new_n581_), .B2(KEYINPUT60), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(KEYINPUT60), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n819_), .B1(KEYINPUT120), .B2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n821_), .B1(KEYINPUT120), .B2(new_n819_), .ZN(new_n822_));
  OAI22_X1  g621(.A1(new_n817_), .A2(new_n818_), .B1(new_n809_), .B2(new_n822_), .ZN(G1341gat));
  AOI21_X1  g622(.A(new_n469_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n824_));
  INV_X1    g623(.A(G127gat), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n650_), .A2(new_n825_), .ZN(new_n826_));
  OAI22_X1  g625(.A1(new_n824_), .A2(new_n825_), .B1(new_n809_), .B2(new_n826_), .ZN(G1342gat));
  INV_X1    g626(.A(G134gat), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(new_n809_), .B2(new_n692_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT121), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT121), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n831_), .B(new_n828_), .C1(new_n809_), .C2(new_n692_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n811_), .A2(new_n812_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n639_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n834_), .A2(new_n828_), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n830_), .A2(new_n832_), .B1(new_n833_), .B2(new_n835_), .ZN(G1343gat));
  NAND4_X1  g635(.A1(new_n665_), .A2(new_n292_), .A3(new_n627_), .A4(new_n618_), .ZN(new_n837_));
  OR2_X1    g636(.A1(new_n806_), .A2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n838_), .A2(new_n431_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(new_n261_), .ZN(G1344gat));
  NOR2_X1   g639(.A1(new_n838_), .A2(new_n581_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(new_n262_), .ZN(G1345gat));
  NOR2_X1   g641(.A1(new_n838_), .A2(new_n469_), .ZN(new_n843_));
  XOR2_X1   g642(.A(KEYINPUT61), .B(G155gat), .Z(new_n844_));
  XNOR2_X1  g643(.A(new_n843_), .B(new_n844_), .ZN(G1346gat));
  OAI21_X1  g644(.A(G162gat), .B1(new_n838_), .B2(new_n834_), .ZN(new_n846_));
  OR2_X1    g645(.A1(new_n692_), .A2(G162gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n838_), .B2(new_n847_), .ZN(G1347gat));
  INV_X1    g647(.A(new_n806_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n389_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n665_), .A2(new_n850_), .A3(new_n628_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n849_), .A2(new_n430_), .A3(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT62), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n852_), .A2(new_n853_), .A3(G169gat), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n853_), .B1(new_n852_), .B2(G169gat), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT122), .ZN(new_n856_));
  INV_X1    g655(.A(new_n851_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n806_), .B2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(KEYINPUT57), .B1(new_n792_), .B2(new_n651_), .ZN(new_n859_));
  AOI211_X1 g658(.A(new_n787_), .B(new_n590_), .C1(new_n791_), .C2(new_n784_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n639_), .B1(new_n796_), .B2(KEYINPUT58), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT119), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n863_), .A2(new_n798_), .A3(new_n797_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n650_), .B1(new_n861_), .B2(new_n864_), .ZN(new_n865_));
  OAI211_X1 g664(.A(KEYINPUT122), .B(new_n851_), .C1(new_n865_), .C2(new_n754_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n858_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  OR2_X1    g667(.A1(new_n431_), .A2(new_n346_), .ZN(new_n869_));
  OAI22_X1  g668(.A1(new_n854_), .A2(new_n855_), .B1(new_n868_), .B2(new_n869_), .ZN(G1348gat));
  NOR2_X1   g669(.A1(new_n665_), .A2(new_n850_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n807_), .A2(G176gat), .A3(new_n593_), .A4(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n581_), .B1(new_n858_), .B2(new_n866_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(G176gat), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(KEYINPUT123), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT123), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n876_), .B(new_n872_), .C1(new_n873_), .C2(G176gat), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(G1349gat));
  NOR2_X1   g677(.A1(new_n469_), .A2(new_n222_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n807_), .A2(new_n650_), .A3(new_n871_), .ZN(new_n880_));
  INV_X1    g679(.A(G183gat), .ZN(new_n881_));
  AOI22_X1  g680(.A1(new_n867_), .A2(new_n879_), .B1(new_n880_), .B2(new_n881_), .ZN(G1350gat));
  OAI21_X1  g681(.A(G190gat), .B1(new_n868_), .B2(new_n834_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n867_), .A2(new_n342_), .A3(new_n591_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1351gat));
  AND3_X1   g684(.A1(new_n700_), .A2(new_n335_), .A3(new_n618_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n849_), .A2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n430_), .ZN(new_n888_));
  XOR2_X1   g687(.A(KEYINPUT124), .B(G197gat), .Z(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1352gat));
  NAND3_X1  g689(.A1(new_n849_), .A2(new_n593_), .A3(new_n886_), .ZN(new_n891_));
  INV_X1    g690(.A(G204gat), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT125), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n849_), .A2(new_n295_), .A3(new_n593_), .A4(new_n886_), .ZN(new_n895_));
  AND3_X1   g694(.A1(new_n893_), .A2(new_n894_), .A3(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n894_), .B1(new_n893_), .B2(new_n895_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1353gat));
  NAND3_X1  g697(.A1(new_n849_), .A2(new_n650_), .A3(new_n886_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n899_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT126), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT63), .B(G211gat), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n849_), .A2(new_n650_), .A3(new_n886_), .A4(new_n902_), .ZN(new_n903_));
  AND3_X1   g702(.A1(new_n900_), .A2(new_n901_), .A3(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n901_), .B1(new_n900_), .B2(new_n903_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1354gat));
  AOI21_X1  g705(.A(G218gat), .B1(new_n887_), .B2(new_n591_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n639_), .A2(G218gat), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(KEYINPUT127), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n907_), .B1(new_n887_), .B2(new_n909_), .ZN(G1355gat));
endmodule


