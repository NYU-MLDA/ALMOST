//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 0 1 1 0 1 0 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n638_, new_n639_, new_n640_, new_n641_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n813_, new_n814_,
    new_n815_, new_n817_, new_n818_, new_n819_, new_n821_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_;
  INV_X1    g000(.A(KEYINPUT12), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G85gat), .A2(G92gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT64), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n204_), .A2(KEYINPUT9), .ZN(new_n205_));
  INV_X1    g004(.A(G85gat), .ZN(new_n206_));
  INV_X1    g005(.A(G92gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n204_), .A2(KEYINPUT9), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n205_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n211_));
  AND3_X1   g010(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n212_));
  AOI21_X1  g011(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n211_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(KEYINPUT65), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n214_), .A2(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(KEYINPUT10), .B(G99gat), .Z(new_n221_));
  INV_X1    g020(.A(G106gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n210_), .A2(new_n220_), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n214_), .A2(new_n219_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G99gat), .A2(G106gat), .ZN(new_n227_));
  AND2_X1   g026(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n228_));
  NOR2_X1   g027(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n227_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  OAI22_X1  g029(.A1(KEYINPUT66), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT67), .B1(new_n226_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT8), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n208_), .A2(new_n203_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT68), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n208_), .A2(KEYINPUT68), .A3(new_n203_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n230_), .A2(new_n231_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(new_n241_), .A3(new_n220_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n233_), .A2(new_n234_), .A3(new_n239_), .A4(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT69), .B1(new_n212_), .B2(new_n213_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n217_), .A2(new_n245_), .A3(new_n218_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n239_), .B1(new_n247_), .B2(new_n232_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT8), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n225_), .B1(new_n243_), .B2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G57gat), .B(G64gat), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n251_), .A2(KEYINPUT11), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(KEYINPUT11), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G71gat), .B(G78gat), .ZN(new_n254_));
  OR3_X1    g053(.A1(new_n252_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n251_), .A2(new_n254_), .A3(KEYINPUT11), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n202_), .B1(new_n250_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n257_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n232_), .B1(new_n214_), .B2(new_n219_), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT8), .B1(new_n260_), .B2(new_n241_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n240_), .A2(new_n220_), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n262_), .A2(KEYINPUT67), .B1(new_n238_), .B2(new_n237_), .ZN(new_n263_));
  AOI22_X1  g062(.A1(new_n261_), .A2(new_n263_), .B1(KEYINPUT8), .B2(new_n248_), .ZN(new_n264_));
  OAI211_X1 g063(.A(KEYINPUT12), .B(new_n259_), .C1(new_n264_), .C2(new_n225_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n258_), .A2(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n239_), .B1(new_n260_), .B2(new_n241_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n242_), .A2(new_n234_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n249_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n269_), .A2(new_n224_), .A3(new_n257_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G230gat), .A2(G233gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n270_), .A2(KEYINPUT71), .A3(new_n271_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n266_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n270_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n250_), .A2(KEYINPUT70), .A3(new_n257_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n250_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n259_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n271_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT72), .B1(new_n276_), .B2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G120gat), .B(G148gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(G204gat), .ZN(new_n286_));
  XOR2_X1   g085(.A(KEYINPUT5), .B(G176gat), .Z(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n270_), .A2(new_n277_), .ZN(new_n289_));
  AOI21_X1  g088(.A(KEYINPUT70), .B1(new_n250_), .B2(new_n257_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n282_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n271_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  AOI211_X1 g092(.A(new_n273_), .B(new_n292_), .C1(new_n250_), .C2(new_n257_), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT71), .B1(new_n270_), .B2(new_n271_), .ZN(new_n295_));
  OAI211_X1 g094(.A(new_n258_), .B(new_n265_), .C1(new_n294_), .C2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT72), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n293_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n284_), .A2(new_n288_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT73), .ZN(new_n300_));
  OR3_X1    g099(.A1(new_n276_), .A2(new_n283_), .A3(new_n288_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n284_), .A2(new_n298_), .A3(new_n302_), .A4(new_n288_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n300_), .A2(new_n301_), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT74), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT74), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n300_), .A2(new_n306_), .A3(new_n301_), .A4(new_n303_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT13), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n305_), .A2(KEYINPUT13), .A3(new_n307_), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G113gat), .B(G141gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G169gat), .B(G197gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n316_), .A2(KEYINPUT83), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT78), .B(G8gat), .ZN(new_n318_));
  INV_X1    g117(.A(G1gat), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT14), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT79), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G15gat), .B(G22gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(G1gat), .B(G8gat), .Z(new_n325_));
  OR2_X1    g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(new_n325_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G29gat), .B(G36gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G43gat), .B(G50gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n328_), .A2(new_n331_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT81), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n328_), .A2(KEYINPUT81), .A3(new_n331_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n332_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G229gat), .A2(G233gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n331_), .B(KEYINPUT15), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n326_), .A2(new_n327_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n341_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n338_), .B(KEYINPUT82), .Z(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  OAI221_X1 g144(.A(new_n317_), .B1(new_n337_), .B2(new_n338_), .C1(new_n343_), .C2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n337_), .A2(new_n338_), .ZN(new_n347_));
  AOI211_X1 g146(.A(new_n341_), .B(new_n345_), .C1(new_n335_), .C2(new_n336_), .ZN(new_n348_));
  OAI22_X1  g147(.A1(new_n347_), .A2(new_n348_), .B1(KEYINPUT83), .B2(new_n316_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n346_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G231gat), .A2(G233gat), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n257_), .B(new_n352_), .Z(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(new_n328_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G183gat), .B(G211gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G127gat), .B(G155gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT17), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n360_), .A2(KEYINPUT17), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n355_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n354_), .B1(KEYINPUT17), .B2(new_n360_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n312_), .A2(new_n351_), .A3(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n281_), .A2(new_n339_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n250_), .A2(new_n331_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G232gat), .A2(G233gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT34), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n368_), .B(new_n369_), .C1(KEYINPUT35), .C2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(KEYINPUT35), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT77), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G134gat), .B(G162gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G190gat), .B(G218gat), .ZN(new_n379_));
  XOR2_X1   g178(.A(new_n378_), .B(new_n379_), .Z(new_n380_));
  NOR2_X1   g179(.A1(new_n380_), .A2(KEYINPUT36), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n375_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n374_), .A2(KEYINPUT77), .A3(new_n381_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT37), .ZN(new_n386_));
  INV_X1    g185(.A(new_n380_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n374_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT36), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n385_), .A2(new_n386_), .A3(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n386_), .B1(new_n385_), .B2(new_n389_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT94), .B(G197gat), .ZN(new_n394_));
  INV_X1    g193(.A(G204gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(G197gat), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n396_), .B(KEYINPUT21), .C1(new_n397_), .C2(new_n395_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT95), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G211gat), .B(G218gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT96), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n397_), .A2(G204gat), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n402_), .B1(new_n394_), .B2(G204gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n399_), .B(new_n401_), .C1(KEYINPUT21), .C2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT97), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n401_), .B1(new_n406_), .B2(new_n404_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n407_), .B(KEYINPUT21), .C1(new_n406_), .C2(new_n404_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n405_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G228gat), .A2(G233gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT93), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n409_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G141gat), .A2(G148gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT91), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT2), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT92), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n417_), .B1(new_n418_), .B2(new_n415_), .ZN(new_n419_));
  INV_X1    g218(.A(G141gat), .ZN(new_n420_));
  INV_X1    g219(.A(G148gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n422_), .A2(KEYINPUT3), .B1(new_n423_), .B2(KEYINPUT92), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n419_), .B(new_n424_), .C1(KEYINPUT3), .C2(new_n422_), .ZN(new_n425_));
  INV_X1    g224(.A(G155gat), .ZN(new_n426_));
  INV_X1    g225(.A(G162gat), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT88), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT88), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n429_), .A2(G155gat), .A3(G162gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n425_), .B(new_n431_), .C1(G155gat), .C2(G162gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(KEYINPUT1), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT89), .ZN(new_n434_));
  AOI22_X1  g233(.A1(new_n433_), .A2(new_n434_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n435_), .B1(new_n434_), .B2(new_n433_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n431_), .A2(KEYINPUT1), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT90), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n422_), .B(new_n415_), .C1(new_n436_), .C2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n414_), .B1(new_n432_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT99), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n442_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n413_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n432_), .A2(new_n440_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT29), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n412_), .B1(new_n447_), .B2(new_n409_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G78gat), .B(G106gat), .ZN(new_n449_));
  INV_X1    g248(.A(G22gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  OR3_X1    g250(.A1(new_n445_), .A2(new_n448_), .A3(new_n451_), .ZN(new_n452_));
  OR3_X1    g251(.A1(new_n446_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n453_));
  INV_X1    g252(.A(G50gat), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT28), .B1(new_n446_), .B2(KEYINPUT29), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n453_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n454_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n451_), .B1(new_n445_), .B2(new_n448_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n452_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n458_), .B1(new_n452_), .B2(new_n459_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G225gat), .A2(G233gat), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT4), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G127gat), .B(G134gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G113gat), .B(G120gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n446_), .A2(new_n466_), .A3(new_n470_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n446_), .A2(KEYINPUT104), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n446_), .A2(KEYINPUT104), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n469_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n470_), .B1(new_n446_), .B2(KEYINPUT104), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n465_), .B(new_n471_), .C1(new_n476_), .C2(new_n466_), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n474_), .A2(new_n475_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n464_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G1gat), .B(G29gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(new_n206_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(KEYINPUT0), .B(G57gat), .ZN(new_n482_));
  XOR2_X1   g281(.A(new_n481_), .B(new_n482_), .Z(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n477_), .A2(new_n479_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(KEYINPUT105), .A2(KEYINPUT33), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT86), .ZN(new_n488_));
  NOR2_X1   g287(.A1(G169gat), .A2(G176gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT85), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n490_), .A2(KEYINPUT24), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G183gat), .A2(G190gat), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT23), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n488_), .B1(new_n491_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT85), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n489_), .B(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT24), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n494_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT86), .ZN(new_n500_));
  NAND2_X1  g299(.A1(KEYINPUT84), .A2(G190gat), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n501_), .A2(KEYINPUT26), .ZN(new_n502_));
  XNOR2_X1  g301(.A(KEYINPUT25), .B(G183gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(KEYINPUT26), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(G169gat), .ZN(new_n506_));
  INV_X1    g305(.A(G176gat), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n490_), .B(KEYINPUT24), .C1(new_n506_), .C2(new_n507_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n495_), .A2(new_n500_), .A3(new_n505_), .A4(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n494_), .ZN(new_n510_));
  OR2_X1    g309(.A1(G183gat), .A2(G190gat), .ZN(new_n511_));
  AOI22_X1  g310(.A1(new_n510_), .A2(new_n511_), .B1(G169gat), .B2(G176gat), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n506_), .A2(KEYINPUT22), .ZN(new_n513_));
  OR2_X1    g312(.A1(new_n513_), .A2(KEYINPUT87), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(KEYINPUT87), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(new_n507_), .A3(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n506_), .A2(KEYINPUT22), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n512_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n509_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n409_), .A2(new_n519_), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n499_), .A2(KEYINPUT102), .ZN(new_n521_));
  XOR2_X1   g320(.A(KEYINPUT26), .B(G190gat), .Z(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT101), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n503_), .B(KEYINPUT100), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n499_), .A2(KEYINPUT102), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n521_), .A2(new_n525_), .A3(new_n508_), .A4(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n513_), .A2(new_n517_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT103), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n512_), .B1(new_n529_), .B2(G176gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n520_), .B(KEYINPUT20), .C1(new_n409_), .C2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G226gat), .A2(G233gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT19), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n532_), .A2(new_n535_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n409_), .A2(new_n519_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n409_), .A2(new_n531_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n537_), .A2(KEYINPUT20), .A3(new_n534_), .A4(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n536_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G8gat), .B(G36gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(G92gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT18), .B(G64gat), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n542_), .B(new_n543_), .Z(new_n544_));
  NOR2_X1   g343(.A1(new_n540_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n544_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n546_), .B1(new_n536_), .B2(new_n539_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n478_), .A2(new_n465_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n471_), .B1(new_n476_), .B2(new_n466_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n549_), .B(new_n483_), .C1(new_n550_), .C2(new_n465_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT105), .B(KEYINPUT33), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n477_), .A2(new_n479_), .A3(new_n484_), .A4(new_n552_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n487_), .A2(new_n548_), .A3(new_n551_), .A4(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(KEYINPUT106), .B1(new_n544_), .B2(KEYINPUT32), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n540_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT106), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n557_), .B1(new_n536_), .B2(new_n539_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n532_), .A2(new_n534_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n537_), .A2(KEYINPUT20), .A3(new_n538_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n559_), .B1(new_n534_), .B2(new_n560_), .ZN(new_n561_));
  OAI211_X1 g360(.A(KEYINPUT32), .B(new_n544_), .C1(new_n558_), .C2(new_n561_), .ZN(new_n562_));
  AND3_X1   g361(.A1(new_n477_), .A2(new_n479_), .A3(new_n484_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n484_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n556_), .B(new_n562_), .C1(new_n563_), .C2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n463_), .B1(new_n554_), .B2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G71gat), .B(G99gat), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G227gat), .A2(G233gat), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n567_), .B(new_n568_), .Z(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT30), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n519_), .B(new_n571_), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n572_), .A2(new_n469_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n469_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G15gat), .B(G43gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT31), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n573_), .A2(new_n574_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n577_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n570_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n580_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n582_), .A2(new_n569_), .A3(new_n578_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n462_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(new_n585_), .A3(new_n460_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n581_), .A2(new_n583_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n587_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n564_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(new_n485_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT27), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n592_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n561_), .A2(new_n546_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n547_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n594_), .A2(new_n595_), .A3(KEYINPUT27), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n593_), .A2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n591_), .A2(new_n597_), .ZN(new_n598_));
  AOI22_X1  g397(.A1(new_n566_), .A2(new_n584_), .B1(new_n589_), .B2(new_n598_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n367_), .A2(new_n393_), .A3(new_n599_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n600_), .A2(new_n319_), .A3(new_n591_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n601_), .A2(KEYINPUT38), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n602_), .A2(KEYINPUT107), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(KEYINPUT38), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(KEYINPUT107), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n554_), .A2(new_n565_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n463_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n606_), .A2(new_n584_), .A3(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n589_), .A2(new_n598_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n385_), .A2(new_n389_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n367_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n591_), .ZN(new_n616_));
  OAI21_X1  g415(.A(G1gat), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n603_), .A2(new_n604_), .A3(new_n605_), .A4(new_n617_), .ZN(G1324gat));
  INV_X1    g417(.A(new_n597_), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n367_), .A2(new_n619_), .A3(new_n613_), .ZN(new_n620_));
  INV_X1    g419(.A(G8gat), .ZN(new_n621_));
  OR3_X1    g420(.A1(new_n620_), .A2(KEYINPUT108), .A3(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(KEYINPUT108), .B1(new_n620_), .B2(new_n621_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(KEYINPUT39), .A3(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n600_), .A2(new_n318_), .A3(new_n597_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT39), .ZN(new_n626_));
  OAI211_X1 g425(.A(KEYINPUT108), .B(new_n626_), .C1(new_n620_), .C2(new_n621_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n624_), .A2(new_n625_), .A3(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(G1325gat));
  INV_X1    g429(.A(G15gat), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n600_), .A2(new_n631_), .A3(new_n587_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G15gat), .B1(new_n615_), .B2(new_n584_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT41), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n633_), .A2(new_n634_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n632_), .B1(new_n635_), .B2(new_n636_), .ZN(G1326gat));
  NAND3_X1  g436(.A1(new_n600_), .A2(new_n450_), .A3(new_n463_), .ZN(new_n638_));
  OAI21_X1  g437(.A(G22gat), .B1(new_n615_), .B2(new_n607_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n639_), .A2(KEYINPUT42), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n639_), .A2(KEYINPUT42), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n638_), .B1(new_n640_), .B2(new_n641_), .ZN(G1327gat));
  NAND3_X1  g441(.A1(new_n312_), .A2(new_n351_), .A3(new_n365_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n643_), .A2(new_n612_), .A3(new_n599_), .ZN(new_n644_));
  AOI21_X1  g443(.A(G29gat), .B1(new_n644_), .B2(new_n591_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT44), .ZN(new_n646_));
  OAI21_X1  g445(.A(KEYINPUT43), .B1(new_n599_), .B2(new_n392_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT43), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n610_), .A2(new_n648_), .A3(new_n393_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n646_), .B1(new_n651_), .B2(new_n643_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n643_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n650_), .A2(new_n653_), .A3(KEYINPUT44), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n591_), .A2(G29gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n645_), .B1(new_n655_), .B2(new_n656_), .ZN(G1328gat));
  INV_X1    g456(.A(G36gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n658_), .B1(new_n655_), .B2(new_n597_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n597_), .B(KEYINPUT110), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n644_), .A2(new_n658_), .A3(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT45), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT46), .ZN(new_n665_));
  OR3_X1    g464(.A1(new_n659_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n659_), .B2(new_n664_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1329gat));
  INV_X1    g467(.A(KEYINPUT111), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n655_), .A2(new_n669_), .A3(G43gat), .A4(new_n587_), .ZN(new_n670_));
  INV_X1    g469(.A(G43gat), .ZN(new_n671_));
  INV_X1    g470(.A(new_n644_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(new_n672_), .B2(new_n584_), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n652_), .A2(new_n654_), .A3(G43gat), .A4(new_n587_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT111), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n670_), .A2(new_n673_), .A3(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT47), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT47), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n670_), .A2(new_n678_), .A3(new_n673_), .A4(new_n675_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(G1330gat));
  AOI21_X1  g479(.A(G50gat), .B1(new_n644_), .B2(new_n463_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n607_), .A2(new_n454_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n655_), .B2(new_n682_), .ZN(G1331gat));
  INV_X1    g482(.A(new_n312_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n351_), .A2(new_n365_), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n684_), .A2(new_n612_), .A3(new_n610_), .A4(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(G57gat), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n686_), .A2(new_n687_), .A3(new_n616_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n599_), .A2(new_n393_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(G57gat), .B1(new_n691_), .B2(new_n591_), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n692_), .A2(KEYINPUT112), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(KEYINPUT112), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n688_), .B1(new_n693_), .B2(new_n694_), .ZN(G1332gat));
  OR3_X1    g494(.A1(new_n690_), .A2(G64gat), .A3(new_n660_), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n686_), .A2(new_n660_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT48), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n697_), .A2(new_n698_), .A3(G64gat), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n698_), .B1(new_n697_), .B2(G64gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n696_), .B1(new_n700_), .B2(new_n701_), .ZN(G1333gat));
  OR3_X1    g501(.A1(new_n690_), .A2(G71gat), .A3(new_n584_), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n686_), .A2(new_n584_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(KEYINPUT113), .B(KEYINPUT49), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(G71gat), .A3(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n705_), .B1(new_n704_), .B2(G71gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n703_), .B1(new_n707_), .B2(new_n708_), .ZN(G1334gat));
  OR3_X1    g508(.A1(new_n690_), .A2(G78gat), .A3(new_n607_), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n686_), .A2(new_n607_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT50), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(new_n712_), .A3(G78gat), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n712_), .B1(new_n711_), .B2(G78gat), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n710_), .B1(new_n714_), .B2(new_n715_), .ZN(G1335gat));
  NOR2_X1   g515(.A1(new_n312_), .A2(new_n351_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n599_), .A2(new_n612_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n717_), .A2(new_n365_), .A3(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT114), .ZN(new_n720_));
  AOI21_X1  g519(.A(G85gat), .B1(new_n720_), .B2(new_n591_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n650_), .A2(new_n365_), .A3(new_n717_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n723_), .A2(new_n206_), .A3(new_n616_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n721_), .A2(new_n724_), .ZN(G1336gat));
  AOI21_X1  g524(.A(G92gat), .B1(new_n720_), .B2(new_n597_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n723_), .A2(new_n207_), .A3(new_n660_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1337gat));
  NAND3_X1  g527(.A1(new_n720_), .A2(new_n221_), .A3(new_n587_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT115), .ZN(new_n730_));
  OAI21_X1  g529(.A(G99gat), .B1(new_n723_), .B2(new_n584_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT115), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n720_), .A2(new_n732_), .A3(new_n221_), .A4(new_n587_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n730_), .A2(new_n731_), .A3(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT51), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT51), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n730_), .A2(new_n736_), .A3(new_n731_), .A4(new_n733_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1338gat));
  NAND3_X1  g537(.A1(new_n720_), .A2(new_n222_), .A3(new_n463_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT52), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n722_), .A2(new_n463_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n741_), .B2(G106gat), .ZN(new_n742_));
  AOI211_X1 g541(.A(KEYINPUT52), .B(new_n222_), .C1(new_n722_), .C2(new_n463_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n739_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g544(.A1(new_n347_), .A2(new_n348_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n343_), .A2(new_n345_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n337_), .A2(new_n344_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  MUX2_X1   g548(.A(new_n746_), .B(new_n749_), .S(new_n315_), .Z(new_n750_));
  AOI21_X1  g549(.A(new_n750_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n276_), .A2(KEYINPUT55), .ZN(new_n752_));
  INV_X1    g551(.A(new_n280_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n292_), .B1(new_n753_), .B2(new_n266_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n276_), .A2(KEYINPUT55), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n752_), .A2(new_n754_), .A3(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n288_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT56), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT56), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n756_), .A2(new_n759_), .A3(new_n288_), .ZN(new_n760_));
  AND4_X1   g559(.A1(new_n351_), .A2(new_n758_), .A3(new_n301_), .A4(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n612_), .B1(new_n751_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT57), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n316_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n746_), .B2(new_n316_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n766_), .A2(new_n758_), .A3(new_n301_), .A4(new_n760_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT58), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n768_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n393_), .A3(new_n770_), .ZN(new_n771_));
  OAI211_X1 g570(.A(KEYINPUT57), .B(new_n612_), .C1(new_n751_), .C2(new_n761_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n764_), .A2(new_n771_), .A3(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n365_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT117), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n310_), .A2(new_n311_), .A3(new_n392_), .A4(new_n685_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT54), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT117), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n773_), .A2(new_n778_), .A3(new_n365_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n775_), .A2(new_n777_), .A3(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT59), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n616_), .A2(new_n588_), .A3(new_n597_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n780_), .A2(new_n781_), .A3(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n774_), .A2(new_n777_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n782_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT59), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n783_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(G113gat), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n787_), .A2(new_n788_), .A3(new_n350_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n785_), .A2(new_n350_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n790_), .A2(G113gat), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n791_), .A2(KEYINPUT116), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n790_), .A2(new_n793_), .A3(G113gat), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n789_), .A2(new_n792_), .A3(new_n794_), .ZN(G1340gat));
  NAND3_X1  g594(.A1(new_n783_), .A2(new_n684_), .A3(new_n786_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT118), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n783_), .A2(KEYINPUT118), .A3(new_n684_), .A4(new_n786_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(G120gat), .A3(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n785_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT60), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n802_), .B1(new_n312_), .B2(G120gat), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n801_), .B(new_n803_), .C1(new_n802_), .C2(G120gat), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n800_), .A2(new_n804_), .ZN(G1341gat));
  INV_X1    g604(.A(G127gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n806_), .B1(new_n785_), .B2(new_n365_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT119), .ZN(new_n808_));
  INV_X1    g607(.A(new_n787_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n365_), .A2(new_n806_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(KEYINPUT120), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n808_), .B1(new_n809_), .B2(new_n811_), .ZN(G1342gat));
  AOI21_X1  g611(.A(G134gat), .B1(new_n801_), .B2(new_n611_), .ZN(new_n813_));
  XOR2_X1   g612(.A(KEYINPUT121), .B(G134gat), .Z(new_n814_));
  NOR2_X1   g613(.A1(new_n392_), .A2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n813_), .B1(new_n809_), .B2(new_n815_), .ZN(G1343gat));
  INV_X1    g615(.A(new_n586_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n784_), .A2(new_n591_), .A3(new_n817_), .A4(new_n660_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n818_), .A2(new_n350_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(new_n420_), .ZN(G1344gat));
  NOR2_X1   g619(.A1(new_n818_), .A2(new_n312_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(new_n421_), .ZN(G1345gat));
  INV_X1    g621(.A(new_n818_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n823_), .A2(new_n426_), .A3(new_n366_), .ZN(new_n824_));
  OAI21_X1  g623(.A(G155gat), .B1(new_n818_), .B2(new_n365_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n824_), .A2(new_n827_), .A3(new_n825_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(G1346gat));
  AOI21_X1  g630(.A(G162gat), .B1(new_n823_), .B2(new_n611_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n392_), .A2(new_n427_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(KEYINPUT123), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n832_), .B1(new_n823_), .B2(new_n834_), .ZN(G1347gat));
  NOR2_X1   g634(.A1(new_n660_), .A2(new_n591_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n587_), .ZN(new_n837_));
  XOR2_X1   g636(.A(new_n837_), .B(KEYINPUT124), .Z(new_n838_));
  NOR2_X1   g637(.A1(new_n838_), .A2(new_n463_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n780_), .A2(new_n839_), .A3(new_n351_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(G169gat), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT62), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n841_), .A2(KEYINPUT125), .A3(new_n842_), .ZN(new_n843_));
  OR2_X1    g642(.A1(new_n842_), .A2(KEYINPUT125), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(KEYINPUT125), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n840_), .A2(G169gat), .A3(new_n844_), .A4(new_n845_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n843_), .B(new_n846_), .C1(new_n529_), .C2(new_n840_), .ZN(G1348gat));
  NAND3_X1  g646(.A1(new_n780_), .A2(new_n839_), .A3(new_n684_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n507_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT126), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n848_), .A2(KEYINPUT126), .A3(new_n507_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n774_), .A2(new_n777_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(new_n463_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n838_), .A2(new_n507_), .A3(new_n312_), .ZN(new_n855_));
  AOI22_X1  g654(.A1(new_n851_), .A2(new_n852_), .B1(new_n854_), .B2(new_n855_), .ZN(G1349gat));
  NOR2_X1   g655(.A1(new_n838_), .A2(new_n365_), .ZN(new_n857_));
  AOI21_X1  g656(.A(G183gat), .B1(new_n854_), .B2(new_n857_), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n780_), .A2(new_n839_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n365_), .A2(new_n524_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n858_), .B1(new_n859_), .B2(new_n860_), .ZN(G1350gat));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n393_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(G190gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n859_), .A2(new_n611_), .A3(new_n523_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(G1351gat));
  NOR2_X1   g664(.A1(new_n853_), .A2(new_n586_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n866_), .A2(new_n836_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n351_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n684_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g670(.A(new_n365_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT127), .ZN(new_n873_));
  OR2_X1    g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n873_), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n866_), .A2(new_n836_), .A3(new_n874_), .A4(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n877_));
  XOR2_X1   g676(.A(new_n876_), .B(new_n877_), .Z(G1354gat));
  AOI21_X1  g677(.A(G218gat), .B1(new_n867_), .B2(new_n611_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n393_), .A2(G218gat), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n867_), .B2(new_n880_), .ZN(G1355gat));
endmodule


