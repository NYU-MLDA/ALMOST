//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 1 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n593_,
    new_n594_, new_n595_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n801_, new_n803_,
    new_n804_, new_n806_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n841_, new_n843_, new_n844_, new_n845_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_;
  XNOR2_X1  g000(.A(G155gat), .B(G162gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT92), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT3), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT2), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(KEYINPUT91), .A3(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n203_), .A2(new_n208_), .ZN(new_n209_));
  AOI21_X1  g008(.A(KEYINPUT91), .B1(new_n205_), .B2(new_n207_), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n204_), .ZN(new_n212_));
  INV_X1    g011(.A(G155gat), .ZN(new_n213_));
  INV_X1    g012(.A(G162gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT1), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n215_), .B1(G155gat), .B2(G162gat), .ZN(new_n216_));
  NOR3_X1   g015(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT1), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n212_), .B(new_n206_), .C1(new_n216_), .C2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n211_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT93), .B(KEYINPUT28), .ZN(new_n220_));
  OR3_X1    g019(.A1(new_n219_), .A2(KEYINPUT29), .A3(new_n220_), .ZN(new_n221_));
  XOR2_X1   g020(.A(G22gat), .B(G50gat), .Z(new_n222_));
  OAI21_X1  g021(.A(new_n220_), .B1(new_n219_), .B2(KEYINPUT29), .ZN(new_n223_));
  AND3_X1   g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n222_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G78gat), .B(G106gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n219_), .A2(KEYINPUT29), .ZN(new_n230_));
  INV_X1    g029(.A(G204gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT95), .B1(new_n231_), .B2(G197gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT95), .ZN(new_n233_));
  INV_X1    g032(.A(G197gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(new_n234_), .A3(G204gat), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n232_), .B(new_n235_), .C1(new_n234_), .C2(G204gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT98), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G211gat), .B(G218gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT97), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT21), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n240_), .B1(new_n239_), .B2(new_n238_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n237_), .A2(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n231_), .A2(G197gat), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n234_), .A2(G204gat), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT21), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT96), .B(KEYINPUT21), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n245_), .B(new_n238_), .C1(new_n236_), .C2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n242_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n230_), .A2(KEYINPUT94), .A3(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G228gat), .A2(G233gat), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n230_), .A2(KEYINPUT94), .A3(new_n250_), .A4(new_n248_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n229_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n254_), .A2(KEYINPUT99), .ZN(new_n255_));
  OAI21_X1  g054(.A(KEYINPUT100), .B1(new_n227_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n252_), .A2(new_n253_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(new_n228_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT99), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT100), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(new_n261_), .A3(new_n226_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n257_), .A2(new_n228_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n263_), .A2(new_n254_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n256_), .A2(new_n262_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(G169gat), .ZN(new_n267_));
  INV_X1    g066(.A(G176gat), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(KEYINPUT86), .B(G176gat), .Z(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT85), .B1(new_n267_), .B2(KEYINPUT22), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT22), .B(G169gat), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n271_), .B(new_n272_), .C1(KEYINPUT85), .C2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT23), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n275_), .A2(G183gat), .A3(G190gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT87), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n275_), .B1(G183gat), .B2(G190gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(G183gat), .A2(G190gat), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n270_), .B(new_n274_), .C1(new_n279_), .C2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT25), .B(G183gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT26), .B(G190gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n284_), .B(KEYINPUT84), .Z(new_n285_));
  NOR3_X1   g084(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n286_));
  XOR2_X1   g085(.A(G169gat), .B(G176gat), .Z(new_n287_));
  AOI21_X1  g086(.A(new_n286_), .B1(new_n287_), .B2(KEYINPUT24), .ZN(new_n288_));
  INV_X1    g087(.A(new_n278_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(new_n276_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n281_), .B1(new_n285_), .B2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT88), .ZN(new_n293_));
  XOR2_X1   g092(.A(G71gat), .B(G99gat), .Z(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT89), .B(G43gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n293_), .B(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(G127gat), .B(G134gat), .Z(new_n298_));
  XOR2_X1   g097(.A(G113gat), .B(G120gat), .Z(new_n299_));
  AOI21_X1  g098(.A(KEYINPUT90), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n298_), .A2(new_n299_), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n300_), .B(new_n301_), .Z(new_n302_));
  OR2_X1    g101(.A1(new_n297_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G227gat), .A2(G233gat), .ZN(new_n304_));
  INV_X1    g103(.A(G15gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT30), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT31), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n297_), .A2(new_n302_), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n303_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n308_), .B1(new_n303_), .B2(new_n309_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n264_), .B1(new_n256_), .B2(new_n262_), .ZN(new_n313_));
  NOR3_X1   g112(.A1(new_n266_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n303_), .A2(new_n309_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n308_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n303_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n256_), .A2(new_n262_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n264_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n319_), .B1(new_n322_), .B2(new_n265_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n314_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G225gat), .A2(G233gat), .ZN(new_n325_));
  XOR2_X1   g124(.A(new_n325_), .B(KEYINPUT103), .Z(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n219_), .A2(new_n302_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n298_), .A2(new_n299_), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n211_), .B(new_n218_), .C1(new_n301_), .C2(new_n329_), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(KEYINPUT102), .B1(new_n331_), .B2(KEYINPUT4), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n328_), .A2(KEYINPUT4), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n331_), .A2(KEYINPUT102), .A3(KEYINPUT4), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n327_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G1gat), .B(G29gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(G85gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT0), .B(G57gat), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n338_), .B(new_n339_), .Z(new_n340_));
  NOR2_X1   g139(.A1(new_n331_), .A2(new_n326_), .ZN(new_n341_));
  OR3_X1    g140(.A1(new_n336_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n340_), .B1(new_n336_), .B2(new_n341_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  XOR2_X1   g144(.A(KEYINPUT105), .B(KEYINPUT27), .Z(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n248_), .ZN(new_n348_));
  XOR2_X1   g147(.A(KEYINPUT101), .B(KEYINPUT24), .Z(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n287_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n349_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n352_));
  AND3_X1   g151(.A1(new_n351_), .A2(new_n284_), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n279_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n290_), .B1(G183gat), .B2(G190gat), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n269_), .B1(new_n271_), .B2(new_n273_), .ZN(new_n356_));
  AOI22_X1  g155(.A1(new_n353_), .A2(new_n354_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT20), .B1(new_n348_), .B2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n358_), .B1(new_n293_), .B2(new_n348_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G226gat), .A2(G233gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT19), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  OR2_X1    g161(.A1(new_n359_), .A2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G8gat), .B(G36gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT18), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G64gat), .B(G92gat), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n365_), .B(new_n366_), .Z(new_n367_));
  OR2_X1    g166(.A1(new_n293_), .A2(new_n348_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT20), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n369_), .B1(new_n348_), .B2(new_n357_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n368_), .A2(new_n362_), .A3(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n363_), .A2(new_n367_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n367_), .B1(new_n363_), .B2(new_n371_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n347_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n362_), .B1(new_n368_), .B2(new_n370_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n359_), .A2(new_n362_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  OAI211_X1 g177(.A(KEYINPUT27), .B(new_n372_), .C1(new_n378_), .C2(new_n367_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n375_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n345_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n367_), .A2(KEYINPUT32), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n363_), .A2(new_n371_), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT104), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n363_), .A2(new_n371_), .A3(KEYINPUT104), .A4(new_n383_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n386_), .B(new_n387_), .C1(new_n378_), .C2(new_n383_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n388_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n374_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n334_), .A2(new_n327_), .A3(new_n335_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n340_), .B1(new_n331_), .B2(new_n326_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n390_), .A2(new_n393_), .A3(new_n372_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n343_), .A2(KEYINPUT33), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT33), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n396_), .B(new_n340_), .C1(new_n336_), .C2(new_n341_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n394_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n389_), .A2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n266_), .A2(new_n313_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n312_), .ZN(new_n401_));
  OAI22_X1  g200(.A1(new_n324_), .A2(new_n382_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n402_));
  XOR2_X1   g201(.A(KEYINPUT70), .B(KEYINPUT12), .Z(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(G85gat), .ZN(new_n405_));
  INV_X1    g204(.A(G92gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G85gat), .A2(G92gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT7), .ZN(new_n410_));
  INV_X1    g209(.A(G99gat), .ZN(new_n411_));
  INV_X1    g210(.A(G106gat), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n410_), .A2(new_n411_), .A3(new_n412_), .A4(KEYINPUT67), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT67), .ZN(new_n414_));
  OAI22_X1  g213(.A1(new_n414_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G99gat), .A2(G106gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT6), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n409_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT8), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT69), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n409_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT6), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n417_), .B(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n413_), .A2(new_n415_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n422_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT69), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n426_), .A2(new_n427_), .A3(KEYINPUT8), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT68), .B1(new_n426_), .B2(KEYINPUT8), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n416_), .A2(new_n418_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT68), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n430_), .A2(new_n431_), .A3(new_n420_), .A4(new_n422_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n421_), .A2(new_n428_), .A3(new_n429_), .A4(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT10), .B(G99gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT65), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n409_), .B1(KEYINPUT9), .B2(new_n406_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT9), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n407_), .A2(new_n437_), .A3(new_n408_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n436_), .A2(KEYINPUT66), .A3(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(KEYINPUT66), .B1(new_n436_), .B2(new_n438_), .ZN(new_n440_));
  OAI221_X1 g239(.A(new_n418_), .B1(new_n435_), .B2(G106gat), .C1(new_n439_), .C2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G57gat), .B(G64gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G71gat), .B(G78gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n443_), .A3(KEYINPUT11), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n442_), .A2(KEYINPUT11), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n445_), .A2(new_n443_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n442_), .A2(KEYINPUT11), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n444_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n433_), .A2(new_n441_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n448_), .B1(new_n433_), .B2(new_n441_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n404_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G230gat), .A2(G233gat), .ZN(new_n453_));
  XOR2_X1   g252(.A(new_n453_), .B(KEYINPUT64), .Z(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n433_), .A2(new_n441_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n448_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(KEYINPUT70), .A2(KEYINPUT12), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n452_), .A2(new_n455_), .A3(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n454_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(G120gat), .B(G148gat), .Z(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT72), .ZN(new_n465_));
  XOR2_X1   g264(.A(G176gat), .B(G204gat), .Z(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  OR2_X1    g268(.A1(new_n463_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n463_), .A2(new_n469_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(KEYINPUT73), .B(KEYINPUT13), .Z(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT13), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n475_), .A2(KEYINPUT73), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n474_), .B1(new_n472_), .B2(new_n476_), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n477_), .A2(KEYINPUT74), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(KEYINPUT74), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(G29gat), .B(G36gat), .Z(new_n481_));
  XOR2_X1   g280(.A(G43gat), .B(G50gat), .Z(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT15), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G15gat), .B(G22gat), .ZN(new_n485_));
  INV_X1    g284(.A(G1gat), .ZN(new_n486_));
  INV_X1    g285(.A(G8gat), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT14), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n485_), .B1(new_n488_), .B2(KEYINPUT79), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n488_), .A2(KEYINPUT79), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G1gat), .B(G8gat), .ZN(new_n491_));
  OR3_X1    g290(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n491_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n484_), .A2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n492_), .A2(new_n483_), .A3(new_n493_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G229gat), .A2(G233gat), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n495_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n483_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n494_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n496_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n497_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n499_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT82), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT83), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT83), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n505_), .A2(new_n506_), .A3(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G113gat), .B(G141gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G169gat), .B(G197gat), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n512_), .B(new_n513_), .Z(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n511_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n508_), .A2(new_n510_), .A3(new_n514_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n480_), .A2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G190gat), .B(G218gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT76), .ZN(new_n522_));
  XOR2_X1   g321(.A(G134gat), .B(G162gat), .Z(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT36), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT36), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n433_), .A2(new_n500_), .A3(new_n441_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n484_), .B1(new_n433_), .B2(new_n441_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT75), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT35), .ZN(new_n531_));
  INV_X1    g330(.A(new_n456_), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n531_), .B(new_n527_), .C1(new_n532_), .C2(new_n484_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G232gat), .A2(G233gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n530_), .A2(new_n533_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n536_), .ZN(new_n538_));
  OAI211_X1 g337(.A(KEYINPUT75), .B(new_n538_), .C1(new_n528_), .C2(new_n529_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n526_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n525_), .B1(new_n540_), .B2(new_n524_), .ZN(new_n541_));
  AOI21_X1  g340(.A(KEYINPUT77), .B1(new_n537_), .B2(new_n539_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n542_), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n544_), .B(new_n525_), .C1(new_n540_), .C2(new_n524_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(new_n545_), .A3(KEYINPUT78), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT37), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n543_), .A2(new_n545_), .A3(KEYINPUT78), .A4(KEYINPUT37), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT17), .ZN(new_n551_));
  XOR2_X1   g350(.A(G127gat), .B(G155gat), .Z(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT16), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G183gat), .B(G211gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G231gat), .A2(G233gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n494_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(new_n448_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT80), .ZN(new_n559_));
  AOI211_X1 g358(.A(new_n551_), .B(new_n555_), .C1(new_n558_), .C2(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n560_), .B1(new_n559_), .B2(new_n558_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n555_), .B(KEYINPUT17), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n558_), .A2(new_n562_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n563_), .A2(KEYINPUT81), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(KEYINPUT81), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n561_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n550_), .A2(new_n566_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n402_), .A2(new_n520_), .A3(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n344_), .B(KEYINPUT106), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n568_), .A2(new_n486_), .A3(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT107), .B(KEYINPUT38), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n571_), .B(new_n572_), .Z(new_n573_));
  NAND2_X1  g372(.A1(new_n543_), .A2(new_n545_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n402_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT109), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n478_), .A2(new_n479_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n566_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n578_), .A2(new_n518_), .A3(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT108), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n577_), .A2(new_n581_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n582_), .A2(new_n344_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n573_), .B1(new_n583_), .B2(new_n486_), .ZN(G1324gat));
  NAND3_X1  g383(.A1(new_n568_), .A2(new_n487_), .A3(new_n380_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n577_), .A2(new_n581_), .A3(new_n380_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT39), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n586_), .A2(new_n587_), .A3(G8gat), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n587_), .B1(new_n586_), .B2(G8gat), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n585_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT40), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(G1325gat));
  AOI21_X1  g391(.A(new_n305_), .B1(new_n582_), .B2(new_n319_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT41), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n568_), .A2(new_n305_), .A3(new_n319_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(G1326gat));
  INV_X1    g395(.A(G22gat), .ZN(new_n597_));
  INV_X1    g396(.A(new_n400_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n597_), .B1(new_n582_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT42), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n568_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(G1327gat));
  INV_X1    g402(.A(new_n520_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n402_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n574_), .A2(new_n579_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n604_), .A2(new_n605_), .A3(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(G29gat), .B1(new_n608_), .B2(new_n344_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT43), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n402_), .A2(new_n610_), .A3(new_n550_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT110), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n402_), .A2(KEYINPUT110), .A3(new_n610_), .A4(new_n550_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n402_), .A2(new_n550_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT43), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n613_), .A2(new_n614_), .A3(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n604_), .A2(new_n579_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT44), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n617_), .A2(KEYINPUT44), .A3(new_n618_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n570_), .A2(G29gat), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n609_), .B1(new_n623_), .B2(new_n624_), .ZN(G1328gat));
  OR2_X1    g424(.A1(new_n380_), .A2(KEYINPUT111), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n380_), .A2(KEYINPUT111), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n629_), .A2(G36gat), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n520_), .A2(new_n630_), .A3(new_n402_), .A4(new_n606_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT45), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT112), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n632_), .B1(new_n633_), .B2(KEYINPUT46), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n621_), .A2(new_n380_), .A3(new_n622_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n634_), .B1(new_n635_), .B2(G36gat), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT46), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n637_), .A2(KEYINPUT112), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n636_), .A2(new_n639_), .ZN(new_n640_));
  AOI211_X1 g439(.A(new_n638_), .B(new_n634_), .C1(new_n635_), .C2(G36gat), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1329gat));
  AND4_X1   g441(.A1(G43gat), .A2(new_n621_), .A3(new_n319_), .A4(new_n622_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT47), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n608_), .A2(new_n319_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n646_), .A2(G43gat), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n644_), .A2(new_n645_), .A3(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(KEYINPUT47), .B1(new_n643_), .B2(new_n647_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1330gat));
  AOI21_X1  g450(.A(G50gat), .B1(new_n608_), .B2(new_n598_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n598_), .A2(G50gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n652_), .B1(new_n623_), .B2(new_n653_), .ZN(G1331gat));
  AND4_X1   g453(.A1(new_n402_), .A2(new_n519_), .A3(new_n480_), .A4(new_n567_), .ZN(new_n655_));
  INV_X1    g454(.A(G57gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(new_n656_), .A3(new_n570_), .ZN(new_n657_));
  AND4_X1   g456(.A1(new_n577_), .A2(new_n519_), .A3(new_n480_), .A4(new_n579_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n658_), .A2(new_n344_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n657_), .B1(new_n659_), .B2(new_n656_), .ZN(G1332gat));
  INV_X1    g459(.A(G64gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n661_), .B1(new_n658_), .B2(new_n628_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT48), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n655_), .A2(new_n661_), .A3(new_n628_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1333gat));
  INV_X1    g465(.A(G71gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n667_), .B1(new_n658_), .B2(new_n319_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT49), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n668_), .B(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n655_), .A2(new_n667_), .A3(new_n319_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1334gat));
  INV_X1    g471(.A(G78gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n673_), .B1(new_n658_), .B2(new_n598_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT50), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n674_), .B(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n655_), .A2(new_n673_), .A3(new_n598_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1335gat));
  NAND2_X1  g477(.A1(new_n480_), .A2(new_n519_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n605_), .A2(new_n679_), .A3(new_n607_), .ZN(new_n680_));
  AOI21_X1  g479(.A(G85gat), .B1(new_n680_), .B2(new_n570_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT113), .Z(new_n682_));
  NOR2_X1   g481(.A1(new_n679_), .A2(new_n579_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n617_), .A2(new_n683_), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT114), .Z(new_n685_));
  NOR2_X1   g484(.A1(new_n345_), .A2(new_n405_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n682_), .B1(new_n685_), .B2(new_n686_), .ZN(G1336gat));
  NAND3_X1  g486(.A1(new_n680_), .A2(new_n406_), .A3(new_n380_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n685_), .A2(new_n628_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(new_n406_), .ZN(G1337gat));
  INV_X1    g489(.A(new_n435_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n680_), .A2(new_n691_), .A3(new_n319_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n617_), .A2(new_n319_), .A3(new_n683_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT115), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n693_), .A2(new_n694_), .A3(G99gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n693_), .B2(G99gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n692_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g497(.A1(new_n680_), .A2(new_n412_), .A3(new_n598_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n617_), .A2(new_n598_), .A3(new_n683_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT52), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n700_), .A2(new_n701_), .A3(G106gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n700_), .B2(G106gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n699_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g504(.A1(new_n314_), .A2(new_n381_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n569_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT59), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n567_), .A2(new_n519_), .A3(new_n477_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT54), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT54), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n567_), .A2(new_n712_), .A3(new_n519_), .A4(new_n477_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n495_), .A2(new_n496_), .A3(new_n503_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n502_), .A2(new_n497_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  MUX2_X1   g517(.A(new_n505_), .B(new_n718_), .S(new_n515_), .Z(new_n719_));
  NAND2_X1  g518(.A1(new_n470_), .A2(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n403_), .B1(new_n458_), .B2(new_n449_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n451_), .B1(KEYINPUT70), .B2(KEYINPUT12), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n454_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT116), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT55), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n461_), .A2(new_n726_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n452_), .A2(KEYINPUT55), .A3(new_n460_), .A4(new_n455_), .ZN(new_n728_));
  OAI211_X1 g527(.A(KEYINPUT116), .B(new_n454_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n725_), .A2(new_n727_), .A3(new_n728_), .A4(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(new_n469_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT56), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n730_), .A2(KEYINPUT56), .A3(new_n469_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n720_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT119), .ZN(new_n736_));
  OAI21_X1  g535(.A(KEYINPUT58), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n720_), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n730_), .A2(KEYINPUT56), .A3(new_n469_), .ZN(new_n739_));
  AOI21_X1  g538(.A(KEYINPUT56), .B1(new_n730_), .B2(new_n469_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n738_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT58), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(KEYINPUT119), .A3(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n737_), .A2(new_n550_), .A3(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n518_), .A2(new_n470_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n472_), .A2(new_n719_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n574_), .B1(new_n746_), .B2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n744_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT121), .ZN(new_n753_));
  INV_X1    g552(.A(new_n574_), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n518_), .B(new_n470_), .C1(new_n739_), .C2(new_n740_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n755_), .B2(new_n747_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT120), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(new_n757_), .A3(KEYINPUT57), .ZN(new_n758_));
  OAI211_X1 g557(.A(KEYINPUT57), .B(new_n574_), .C1(new_n746_), .C2(new_n748_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT120), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT121), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n744_), .A2(new_n762_), .A3(new_n751_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n753_), .A2(new_n761_), .A3(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n566_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT122), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n715_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  AOI22_X1  g566(.A1(new_n752_), .A2(KEYINPUT121), .B1(new_n760_), .B2(new_n758_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n579_), .B1(new_n768_), .B2(new_n763_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT122), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n709_), .B1(new_n767_), .B2(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n751_), .B(KEYINPUT118), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n761_), .A2(new_n744_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n566_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n714_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n708_), .B1(new_n775_), .B2(new_n707_), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT123), .B1(new_n771_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n709_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n714_), .B1(new_n769_), .B2(KEYINPUT122), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n765_), .A2(new_n766_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n778_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT123), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n775_), .A2(new_n707_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT59), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n781_), .A2(new_n782_), .A3(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n777_), .A2(new_n518_), .A3(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(G113gat), .ZN(new_n787_));
  OR3_X1    g586(.A1(new_n783_), .A2(G113gat), .A3(new_n519_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(G1340gat));
  NOR3_X1   g588(.A1(new_n771_), .A2(new_n578_), .A3(new_n776_), .ZN(new_n790_));
  INV_X1    g589(.A(G120gat), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(new_n578_), .B2(KEYINPUT60), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n792_), .B1(KEYINPUT60), .B2(new_n791_), .ZN(new_n793_));
  OAI22_X1  g592(.A1(new_n790_), .A2(new_n791_), .B1(new_n783_), .B2(new_n793_), .ZN(G1341gat));
  NAND3_X1  g593(.A1(new_n777_), .A2(new_n579_), .A3(new_n785_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(G127gat), .ZN(new_n796_));
  OR3_X1    g595(.A1(new_n783_), .A2(G127gat), .A3(new_n566_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(G1342gat));
  NAND3_X1  g597(.A1(new_n777_), .A2(new_n550_), .A3(new_n785_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(G134gat), .ZN(new_n800_));
  OR3_X1    g599(.A1(new_n783_), .A2(G134gat), .A3(new_n574_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(G1343gat));
  NAND4_X1  g601(.A1(new_n775_), .A2(new_n323_), .A3(new_n570_), .A4(new_n629_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n803_), .A2(new_n519_), .ZN(new_n804_));
  XOR2_X1   g603(.A(new_n804_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g604(.A1(new_n803_), .A2(new_n578_), .ZN(new_n806_));
  XOR2_X1   g605(.A(new_n806_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g606(.A1(new_n803_), .A2(new_n566_), .ZN(new_n808_));
  XOR2_X1   g607(.A(KEYINPUT61), .B(G155gat), .Z(new_n809_));
  XNOR2_X1  g608(.A(new_n808_), .B(new_n809_), .ZN(G1346gat));
  INV_X1    g609(.A(new_n550_), .ZN(new_n811_));
  OAI21_X1  g610(.A(G162gat), .B1(new_n803_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n754_), .A2(new_n214_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n803_), .B2(new_n813_), .ZN(G1347gat));
  INV_X1    g613(.A(KEYINPUT62), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n598_), .B1(new_n767_), .B2(new_n770_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n628_), .A2(new_n569_), .A3(new_n319_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n817_), .A2(new_n519_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(KEYINPUT124), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n816_), .A2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n815_), .B1(new_n820_), .B2(G169gat), .ZN(new_n821_));
  AOI211_X1 g620(.A(KEYINPUT62), .B(new_n267_), .C1(new_n816_), .C2(new_n819_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n817_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n400_), .B(new_n823_), .C1(new_n779_), .C2(new_n780_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n518_), .A2(new_n273_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(KEYINPUT125), .ZN(new_n826_));
  OAI22_X1  g625(.A1(new_n821_), .A2(new_n822_), .B1(new_n824_), .B2(new_n826_), .ZN(G1348gat));
  OAI21_X1  g626(.A(new_n271_), .B1(new_n824_), .B2(new_n578_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n598_), .B1(new_n774_), .B2(new_n714_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n829_), .A2(G176gat), .A3(new_n480_), .A4(new_n823_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT126), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n828_), .A2(KEYINPUT126), .A3(new_n830_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(G1349gat));
  NOR2_X1   g634(.A1(new_n817_), .A2(new_n566_), .ZN(new_n836_));
  AOI21_X1  g635(.A(G183gat), .B1(new_n829_), .B2(new_n836_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n817_), .A2(new_n282_), .A3(new_n566_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n837_), .B1(new_n816_), .B2(new_n838_), .ZN(G1350gat));
  OAI21_X1  g638(.A(G190gat), .B1(new_n824_), .B2(new_n811_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n754_), .A2(new_n283_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n824_), .B2(new_n841_), .ZN(G1351gat));
  NOR2_X1   g641(.A1(new_n629_), .A2(new_n344_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n775_), .A2(new_n323_), .A3(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n844_), .A2(new_n519_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(new_n234_), .ZN(G1352gat));
  NOR2_X1   g645(.A1(new_n844_), .A2(new_n578_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(new_n231_), .ZN(G1353gat));
  INV_X1    g647(.A(KEYINPUT63), .ZN(new_n849_));
  INV_X1    g648(.A(G211gat), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n579_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  OR3_X1    g650(.A1(new_n844_), .A2(KEYINPUT127), .A3(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(KEYINPUT127), .B1(new_n844_), .B2(new_n851_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n849_), .A2(new_n850_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n854_), .B(new_n855_), .ZN(G1354gat));
  OAI21_X1  g655(.A(G218gat), .B1(new_n844_), .B2(new_n811_), .ZN(new_n857_));
  OR2_X1    g656(.A1(new_n574_), .A2(G218gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n844_), .B2(new_n858_), .ZN(G1355gat));
endmodule


