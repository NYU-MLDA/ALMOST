//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 0 1 0 0 0 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n628_, new_n629_, new_n630_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n662_,
    new_n663_, new_n664_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n801_,
    new_n802_, new_n803_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n814_, new_n816_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n853_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G211gat), .B(G218gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT87), .B(G197gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(G204gat), .ZN(new_n205_));
  INV_X1    g004(.A(G197gat), .ZN(new_n206_));
  INV_X1    g005(.A(G204gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT21), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n207_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT88), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n210_), .B1(new_n206_), .B2(G204gat), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n209_), .B(new_n211_), .C1(new_n204_), .C2(new_n207_), .ZN(new_n212_));
  OAI221_X1 g011(.A(new_n203_), .B1(new_n205_), .B2(new_n208_), .C1(new_n212_), .C2(KEYINPUT21), .ZN(new_n213_));
  INV_X1    g012(.A(new_n203_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(KEYINPUT21), .A3(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT3), .ZN(new_n218_));
  INV_X1    g017(.A(G141gat), .ZN(new_n219_));
  INV_X1    g018(.A(G148gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G141gat), .A2(G148gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT2), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n221_), .A2(new_n224_), .A3(new_n225_), .A4(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G155gat), .A2(G162gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G155gat), .A2(G162gat), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n227_), .A2(new_n228_), .A3(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT83), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n219_), .A2(new_n220_), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT82), .B1(new_n228_), .B2(KEYINPUT1), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n228_), .A2(KEYINPUT1), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(new_n230_), .A3(new_n235_), .ZN(new_n236_));
  NOR3_X1   g035(.A1(new_n228_), .A2(KEYINPUT82), .A3(KEYINPUT1), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n222_), .B(new_n233_), .C1(new_n236_), .C2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n232_), .A2(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n217_), .B1(new_n239_), .B2(KEYINPUT29), .ZN(new_n240_));
  INV_X1    g039(.A(G78gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(KEYINPUT85), .B(G228gat), .Z(new_n243_));
  XOR2_X1   g042(.A(KEYINPUT86), .B(G233gat), .Z(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(G106gat), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n242_), .A2(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n242_), .A2(new_n246_), .ZN(new_n248_));
  XOR2_X1   g047(.A(KEYINPUT84), .B(KEYINPUT28), .Z(new_n249_));
  OR3_X1    g048(.A1(new_n239_), .A2(KEYINPUT29), .A3(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n249_), .B1(new_n239_), .B2(KEYINPUT29), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(G22gat), .B(G50gat), .Z(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT89), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n250_), .A2(new_n253_), .A3(new_n251_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  OR3_X1    g057(.A1(new_n247_), .A2(new_n248_), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n255_), .A2(new_n257_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT89), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n261_), .B(new_n258_), .C1(new_n247_), .C2(new_n248_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n259_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G183gat), .A2(G190gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT23), .ZN(new_n266_));
  XOR2_X1   g065(.A(KEYINPUT77), .B(G183gat), .Z(new_n267_));
  OAI21_X1  g066(.A(new_n266_), .B1(G190gat), .B2(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(G169gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(G169gat), .A2(G176gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT78), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n273_), .A2(KEYINPUT24), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT24), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n275_), .B1(G169gat), .B2(G176gat), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n274_), .B1(new_n273_), .B2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n265_), .B(KEYINPUT23), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(KEYINPUT26), .B(G190gat), .Z(new_n280_));
  NAND2_X1  g079(.A1(new_n267_), .A2(KEYINPUT25), .ZN(new_n281_));
  OR2_X1    g080(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n280_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n271_), .B1(new_n279_), .B2(new_n283_), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n284_), .A2(new_n216_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT20), .ZN(new_n286_));
  XOR2_X1   g085(.A(KEYINPUT25), .B(G183gat), .Z(new_n287_));
  OAI211_X1 g086(.A(new_n277_), .B(new_n278_), .C1(new_n280_), .C2(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n266_), .B1(G183gat), .B2(G190gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(new_n270_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n286_), .B1(new_n291_), .B2(new_n216_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n285_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G226gat), .A2(G233gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT19), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(G8gat), .B(G36gat), .Z(new_n297_));
  XNOR2_X1  g096(.A(G64gat), .B(G92gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n299_), .B(new_n300_), .Z(new_n301_));
  NAND2_X1  g100(.A1(new_n284_), .A2(new_n216_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n295_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n288_), .A2(new_n217_), .A3(new_n290_), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n302_), .A2(KEYINPUT20), .A3(new_n303_), .A4(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n296_), .A2(new_n301_), .A3(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(KEYINPUT92), .B(KEYINPUT20), .Z(new_n307_));
  NAND3_X1  g106(.A1(new_n302_), .A2(new_n304_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n295_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n285_), .A2(new_n292_), .A3(new_n303_), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n306_), .B(KEYINPUT27), .C1(new_n311_), .C2(new_n301_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n301_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n303_), .B1(new_n285_), .B2(new_n292_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n305_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n313_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n306_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT27), .ZN(new_n318_));
  AOI21_X1  g117(.A(KEYINPUT93), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT93), .ZN(new_n320_));
  AOI211_X1 g119(.A(new_n320_), .B(KEYINPUT27), .C1(new_n306_), .C2(new_n316_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n312_), .B1(new_n319_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT94), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  OAI211_X1 g123(.A(KEYINPUT94), .B(new_n312_), .C1(new_n319_), .C2(new_n321_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n264_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G127gat), .B(G134gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT79), .ZN(new_n328_));
  XOR2_X1   g127(.A(G113gat), .B(G120gat), .Z(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT80), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G71gat), .B(G99gat), .ZN(new_n332_));
  INV_X1    g131(.A(G43gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT31), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n331_), .B(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G227gat), .A2(G233gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(G15gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT30), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n336_), .B(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n284_), .B(KEYINPUT81), .Z(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n340_), .A2(new_n342_), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G225gat), .A2(G233gat), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  XOR2_X1   g146(.A(KEYINPUT91), .B(KEYINPUT4), .Z(new_n348_));
  NAND3_X1  g147(.A1(new_n331_), .A2(new_n239_), .A3(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n331_), .A2(new_n239_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n330_), .A2(new_n232_), .A3(new_n238_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT4), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n347_), .B(new_n349_), .C1(new_n352_), .C2(new_n353_), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n350_), .A2(new_n351_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(new_n346_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G1gat), .B(G29gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(G85gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT0), .B(G57gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n358_), .B(new_n359_), .Z(new_n360_));
  NAND3_X1  g159(.A1(new_n354_), .A2(new_n356_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n360_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n345_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT33), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n361_), .A2(new_n367_), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n306_), .A2(new_n316_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n354_), .A2(new_n356_), .A3(KEYINPUT33), .A4(new_n360_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n360_), .B1(new_n355_), .B2(new_n347_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n349_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n371_), .B1(new_n347_), .B2(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n368_), .A2(new_n369_), .A3(new_n370_), .A4(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n301_), .A2(KEYINPUT32), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n375_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n314_), .A2(new_n315_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n376_), .B1(new_n377_), .B2(new_n375_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n378_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n374_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n364_), .A2(new_n259_), .A3(new_n262_), .ZN(new_n381_));
  OAI22_X1  g180(.A1(new_n380_), .A2(new_n264_), .B1(new_n322_), .B2(new_n381_), .ZN(new_n382_));
  AOI22_X1  g181(.A1(new_n326_), .A2(new_n366_), .B1(new_n382_), .B2(new_n345_), .ZN(new_n383_));
  XOR2_X1   g182(.A(G134gat), .B(G162gat), .Z(new_n384_));
  XNOR2_X1  g183(.A(G190gat), .B(G218gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G232gat), .A2(G233gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT34), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n390_), .A2(KEYINPUT35), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G29gat), .B(G36gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G43gat), .B(G50gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT15), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT64), .ZN(new_n396_));
  OR2_X1    g195(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n397_));
  INV_X1    g196(.A(G106gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(G85gat), .ZN(new_n401_));
  INV_X1    g200(.A(G92gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G85gat), .A2(G92gat), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(KEYINPUT9), .A3(new_n404_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n400_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G99gat), .A2(G106gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT6), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT6), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n409_), .A2(G99gat), .A3(G106gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n404_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT9), .ZN(new_n412_));
  AOI22_X1  g211(.A1(new_n408_), .A2(new_n410_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n396_), .B1(new_n406_), .B2(new_n413_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n413_), .A2(new_n396_), .A3(new_n405_), .A4(new_n400_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT65), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n403_), .A2(new_n417_), .A3(new_n404_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT7), .ZN(new_n419_));
  INV_X1    g218(.A(G99gat), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(new_n420_), .A3(new_n398_), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n408_), .A2(new_n410_), .ZN(new_n424_));
  AOI211_X1 g223(.A(KEYINPUT8), .B(new_n418_), .C1(new_n423_), .C2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT8), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n424_), .A2(new_n422_), .A3(new_n421_), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n403_), .A2(new_n417_), .A3(new_n404_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n426_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  OAI22_X1  g228(.A1(new_n414_), .A2(new_n416_), .B1(new_n425_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n395_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n391_), .B1(new_n432_), .B2(KEYINPUT71), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT66), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n430_), .A2(new_n434_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n408_), .A2(new_n410_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n421_), .A2(new_n422_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n428_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT8), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n427_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n400_), .A2(new_n405_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n411_), .A2(new_n412_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n424_), .A2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT64), .B1(new_n442_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(new_n415_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n441_), .A2(new_n446_), .A3(KEYINPUT66), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n435_), .A2(new_n394_), .A3(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n431_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n390_), .A2(KEYINPUT35), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n433_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n448_), .A2(KEYINPUT71), .A3(new_n431_), .A4(new_n391_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n388_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT73), .B(KEYINPUT36), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n386_), .B(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n451_), .A2(new_n452_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT74), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n451_), .A2(KEYINPUT74), .A3(new_n452_), .A4(new_n455_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n453_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n460_), .B(KEYINPUT97), .Z(new_n461_));
  NOR2_X1   g260(.A1(new_n383_), .A2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G15gat), .B(G22gat), .ZN(new_n463_));
  INV_X1    g262(.A(G8gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G1gat), .B(G8gat), .ZN(new_n467_));
  XOR2_X1   g266(.A(new_n466_), .B(new_n467_), .Z(new_n468_));
  NAND2_X1  g267(.A1(G231gat), .A2(G233gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G57gat), .B(G64gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT11), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT67), .B(G71gat), .ZN(new_n474_));
  AOI22_X1  g273(.A1(new_n472_), .A2(new_n473_), .B1(new_n474_), .B2(new_n241_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n241_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT68), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n479_), .B1(new_n471_), .B2(KEYINPUT11), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n471_), .A2(KEYINPUT11), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n481_), .A2(KEYINPUT68), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n478_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(KEYINPUT68), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n471_), .A2(new_n479_), .A3(KEYINPUT11), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n475_), .A2(new_n484_), .A3(new_n477_), .A4(new_n485_), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n483_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n470_), .B(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT17), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G127gat), .B(G155gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT16), .ZN(new_n491_));
  XOR2_X1   g290(.A(G183gat), .B(G211gat), .Z(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  NOR3_X1   g292(.A1(new_n488_), .A2(new_n489_), .A3(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(KEYINPUT17), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n488_), .A2(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n441_), .A2(KEYINPUT66), .A3(new_n446_), .ZN(new_n498_));
  AOI21_X1  g297(.A(KEYINPUT66), .B1(new_n441_), .B2(new_n446_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n483_), .A2(new_n486_), .ZN(new_n501_));
  OR3_X1    g300(.A1(new_n500_), .A2(KEYINPUT69), .A3(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(G230gat), .ZN(new_n503_));
  INV_X1    g302(.A(G233gat), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n487_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n435_), .A2(new_n447_), .A3(new_n501_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(new_n507_), .A3(KEYINPUT69), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n502_), .A2(new_n505_), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n430_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n483_), .A2(new_n486_), .A3(KEYINPUT12), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT12), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n512_), .B1(new_n506_), .B2(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n505_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n509_), .A2(new_n516_), .ZN(new_n517_));
  XOR2_X1   g316(.A(G120gat), .B(G148gat), .Z(new_n518_));
  XNOR2_X1  g317(.A(G176gat), .B(G204gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n517_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n509_), .A2(new_n516_), .A3(new_n522_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT13), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n524_), .A2(KEYINPUT13), .A3(new_n525_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(KEYINPUT75), .B1(new_n468_), .B2(new_n394_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n468_), .A2(new_n394_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n533_), .A2(G229gat), .A3(G233gat), .ZN(new_n534_));
  INV_X1    g333(.A(new_n468_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n395_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G229gat), .A2(G233gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n468_), .A2(new_n394_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n534_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G113gat), .B(G141gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G169gat), .B(G197gat), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n541_), .B(new_n542_), .Z(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n540_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n534_), .A2(new_n539_), .A3(new_n543_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n530_), .A2(new_n548_), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n462_), .A2(new_n497_), .A3(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n202_), .B1(new_n550_), .B2(new_n365_), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n551_), .B(KEYINPUT98), .Z(new_n552_));
  XOR2_X1   g351(.A(new_n547_), .B(KEYINPUT76), .Z(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n383_), .A2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n528_), .A2(new_n497_), .A3(new_n529_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT37), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n453_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n456_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n559_), .B1(new_n460_), .B2(KEYINPUT37), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n556_), .A2(new_n560_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n555_), .A2(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(KEYINPUT95), .B(KEYINPUT38), .Z(new_n563_));
  AOI21_X1  g362(.A(G1gat), .B1(new_n563_), .B2(KEYINPUT96), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n562_), .A2(new_n365_), .A3(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n563_), .A2(KEYINPUT96), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n552_), .A2(new_n567_), .ZN(G1324gat));
  NAND2_X1  g367(.A1(new_n324_), .A2(new_n325_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n562_), .A2(new_n464_), .A3(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT39), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n550_), .A2(new_n570_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n572_), .B1(new_n573_), .B2(G8gat), .ZN(new_n574_));
  AOI211_X1 g373(.A(KEYINPUT39), .B(new_n464_), .C1(new_n550_), .C2(new_n570_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n571_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n576_), .B(new_n578_), .ZN(G1325gat));
  INV_X1    g378(.A(G15gat), .ZN(new_n580_));
  INV_X1    g379(.A(new_n345_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n580_), .B1(new_n550_), .B2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT41), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n562_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(G1326gat));
  INV_X1    g384(.A(G22gat), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n586_), .B1(new_n550_), .B2(new_n264_), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n587_), .B(KEYINPUT42), .Z(new_n588_));
  NAND3_X1  g387(.A1(new_n562_), .A2(new_n586_), .A3(new_n264_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(G1327gat));
  INV_X1    g389(.A(new_n497_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n460_), .A2(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n530_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n555_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(G29gat), .B1(new_n595_), .B2(new_n365_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n549_), .A2(new_n591_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT100), .ZN(new_n598_));
  INV_X1    g397(.A(new_n560_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n383_), .A2(KEYINPUT43), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT43), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n326_), .A2(new_n366_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n264_), .B1(new_n374_), .B2(new_n379_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n322_), .A2(new_n381_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n345_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n601_), .B1(new_n606_), .B2(new_n560_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n598_), .B1(new_n600_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT44), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT43), .B1(new_n383_), .B2(new_n599_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n606_), .A2(new_n601_), .A3(new_n560_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n613_), .A2(KEYINPUT44), .A3(new_n598_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n610_), .A2(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n365_), .A2(G29gat), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n596_), .B1(new_n615_), .B2(new_n616_), .ZN(G1328gat));
  NAND3_X1  g416(.A1(new_n610_), .A2(new_n570_), .A3(new_n614_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(G36gat), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n594_), .A2(G36gat), .A3(new_n569_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT45), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n619_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT46), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n619_), .A2(new_n622_), .A3(KEYINPUT46), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(G1329gat));
  NAND4_X1  g426(.A1(new_n610_), .A2(G43gat), .A3(new_n581_), .A4(new_n614_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n333_), .B1(new_n594_), .B2(new_n345_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g430(.A1(new_n594_), .A2(G50gat), .A3(new_n263_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n610_), .A2(new_n264_), .A3(new_n614_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n633_), .A2(KEYINPUT101), .ZN(new_n634_));
  OAI21_X1  g433(.A(G50gat), .B1(new_n633_), .B2(KEYINPUT101), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n632_), .B1(new_n634_), .B2(new_n635_), .ZN(G1331gat));
  NAND2_X1  g435(.A1(new_n530_), .A2(new_n497_), .ZN(new_n637_));
  NOR4_X1   g436(.A1(new_n383_), .A2(new_n461_), .A3(new_n553_), .A4(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(new_n365_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n637_), .A2(new_n560_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n641_), .A2(KEYINPUT102), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(KEYINPUT102), .ZN(new_n643_));
  NOR4_X1   g442(.A1(new_n383_), .A2(new_n642_), .A3(new_n643_), .A4(new_n547_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n364_), .A2(G57gat), .ZN(new_n645_));
  AOI22_X1  g444(.A1(new_n639_), .A2(G57gat), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT103), .ZN(G1332gat));
  INV_X1    g446(.A(G64gat), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n648_), .B1(new_n638_), .B2(new_n570_), .ZN(new_n649_));
  XOR2_X1   g448(.A(KEYINPUT104), .B(KEYINPUT48), .Z(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n644_), .A2(new_n648_), .A3(new_n570_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(G1333gat));
  INV_X1    g452(.A(G71gat), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n644_), .A2(new_n654_), .A3(new_n581_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT49), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n638_), .A2(new_n581_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n656_), .B1(new_n657_), .B2(G71gat), .ZN(new_n658_));
  AOI211_X1 g457(.A(KEYINPUT49), .B(new_n654_), .C1(new_n638_), .C2(new_n581_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n655_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT105), .Z(G1334gat));
  AOI21_X1  g460(.A(new_n241_), .B1(new_n638_), .B2(new_n264_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT50), .Z(new_n663_));
  NAND3_X1  g462(.A1(new_n644_), .A2(new_n241_), .A3(new_n264_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1335gat));
  NOR2_X1   g464(.A1(new_n383_), .A2(new_n547_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n530_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n667_), .A2(new_n592_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n401_), .B1(new_n669_), .B2(new_n364_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT106), .Z(new_n671_));
  NAND3_X1  g470(.A1(new_n530_), .A2(new_n591_), .A3(new_n548_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT107), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n673_), .B1(new_n600_), .B2(new_n607_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n611_), .A2(new_n612_), .A3(KEYINPUT107), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n672_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n364_), .A2(new_n401_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n671_), .B1(new_n676_), .B2(new_n677_), .ZN(G1336gat));
  OAI21_X1  g477(.A(new_n402_), .B1(new_n669_), .B2(new_n569_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT108), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n569_), .A2(new_n402_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n676_), .B2(new_n681_), .ZN(G1337gat));
  NAND2_X1  g481(.A1(new_n674_), .A2(new_n675_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n672_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n683_), .A2(new_n581_), .A3(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(G99gat), .ZN(new_n686_));
  INV_X1    g485(.A(new_n669_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n687_), .A2(new_n581_), .A3(new_n397_), .A4(new_n399_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n686_), .A2(KEYINPUT109), .A3(KEYINPUT51), .A4(new_n688_), .ZN(new_n689_));
  OR2_X1    g488(.A1(KEYINPUT109), .A2(KEYINPUT51), .ZN(new_n690_));
  NAND2_X1  g489(.A1(KEYINPUT109), .A2(KEYINPUT51), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n420_), .B1(new_n676_), .B2(new_n581_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n688_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n690_), .B(new_n691_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n689_), .A2(new_n694_), .ZN(G1338gat));
  NAND3_X1  g494(.A1(new_n687_), .A2(new_n398_), .A3(new_n264_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT110), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n672_), .A2(new_n263_), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n697_), .B(new_n698_), .C1(new_n600_), .C2(new_n607_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(G106gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n697_), .B1(new_n613_), .B2(new_n698_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n700_), .A2(new_n701_), .A3(KEYINPUT52), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT52), .ZN(new_n703_));
  INV_X1    g502(.A(new_n698_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n704_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n398_), .B1(new_n705_), .B2(new_n697_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n698_), .B1(new_n600_), .B2(new_n607_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT110), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n703_), .B1(new_n706_), .B2(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n696_), .B1(new_n702_), .B2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT53), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT53), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n712_), .B(new_n696_), .C1(new_n702_), .C2(new_n709_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1339gat));
  INV_X1    g513(.A(KEYINPUT54), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n561_), .B2(new_n554_), .ZN(new_n716_));
  NOR4_X1   g515(.A1(new_n556_), .A2(new_n553_), .A3(new_n560_), .A4(KEYINPUT54), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n533_), .A2(new_n537_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n537_), .B1(new_n468_), .B2(new_n394_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n543_), .B1(new_n536_), .B2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n546_), .A2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n525_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n514_), .A2(KEYINPUT55), .A3(new_n515_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n487_), .A2(KEYINPUT12), .A3(new_n430_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n501_), .B1(new_n435_), .B2(new_n447_), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n726_), .B(new_n507_), .C1(new_n727_), .C2(KEYINPUT12), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n505_), .ZN(new_n729_));
  AOI21_X1  g528(.A(KEYINPUT55), .B1(new_n514_), .B2(new_n515_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT111), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n725_), .B(new_n729_), .C1(new_n730_), .C2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT55), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n726_), .B1(new_n727_), .B2(KEYINPUT12), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n507_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n733_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n736_), .A2(KEYINPUT111), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n523_), .B1(new_n732_), .B2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT56), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  OAI211_X1 g539(.A(KEYINPUT56), .B(new_n523_), .C1(new_n732_), .C2(new_n737_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n724_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n599_), .B1(new_n742_), .B2(KEYINPUT58), .ZN(new_n743_));
  XNOR2_X1  g542(.A(KEYINPUT113), .B(KEYINPUT58), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n744_), .B1(new_n742_), .B2(KEYINPUT112), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n746_));
  AOI211_X1 g545(.A(new_n746_), .B(new_n724_), .C1(new_n740_), .C2(new_n741_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n743_), .B1(new_n745_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n460_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n547_), .A2(new_n525_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n750_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n526_), .A2(new_n723_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n749_), .B1(new_n751_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT57), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n750_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n741_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n736_), .A2(KEYINPUT111), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n516_), .A2(new_n731_), .A3(new_n733_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n759_), .A2(new_n760_), .A3(new_n725_), .A4(new_n729_), .ZN(new_n761_));
  AOI21_X1  g560(.A(KEYINPUT56), .B1(new_n761_), .B2(new_n523_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n757_), .B1(new_n758_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n752_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n764_), .A2(KEYINPUT57), .A3(new_n749_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n748_), .A2(new_n756_), .A3(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n718_), .B1(new_n766_), .B2(new_n591_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n326_), .A2(new_n365_), .A3(new_n581_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(G113gat), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n770_), .A3(new_n547_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT59), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n772_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n768_), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT57), .B1(new_n764_), .B2(new_n749_), .ZN(new_n775_));
  AOI211_X1 g574(.A(new_n755_), .B(new_n460_), .C1(new_n763_), .C2(new_n752_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n497_), .B1(new_n777_), .B2(new_n748_), .ZN(new_n778_));
  OAI211_X1 g577(.A(KEYINPUT59), .B(new_n774_), .C1(new_n778_), .C2(new_n718_), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n773_), .A2(KEYINPUT114), .A3(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT114), .B1(new_n773_), .B2(new_n779_), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n780_), .A2(new_n781_), .A3(new_n554_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n771_), .B1(new_n782_), .B2(new_n770_), .ZN(G1340gat));
  NOR2_X1   g582(.A1(new_n667_), .A2(KEYINPUT60), .ZN(new_n784_));
  INV_X1    g583(.A(G120gat), .ZN(new_n785_));
  MUX2_X1   g584(.A(KEYINPUT60), .B(new_n784_), .S(new_n785_), .Z(new_n786_));
  NAND2_X1  g585(.A1(new_n769_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n769_), .A2(KEYINPUT115), .A3(new_n786_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n667_), .B1(new_n773_), .B2(new_n779_), .ZN(new_n792_));
  OAI21_X1  g591(.A(G120gat), .B1(new_n792_), .B2(KEYINPUT116), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n794_));
  AOI211_X1 g593(.A(new_n794_), .B(new_n667_), .C1(new_n773_), .C2(new_n779_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n791_), .B1(new_n793_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT117), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  OAI211_X1 g597(.A(KEYINPUT117), .B(new_n791_), .C1(new_n793_), .C2(new_n795_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(G1341gat));
  INV_X1    g599(.A(G127gat), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n769_), .A2(new_n801_), .A3(new_n497_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n780_), .A2(new_n781_), .A3(new_n591_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n803_), .B2(new_n801_), .ZN(G1342gat));
  AOI21_X1  g603(.A(G134gat), .B1(new_n769_), .B2(new_n461_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n780_), .A2(new_n781_), .ZN(new_n806_));
  XOR2_X1   g605(.A(KEYINPUT118), .B(G134gat), .Z(new_n807_));
  NAND2_X1  g606(.A1(new_n560_), .A2(new_n807_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT119), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n805_), .B1(new_n806_), .B2(new_n809_), .ZN(G1343gat));
  INV_X1    g609(.A(new_n767_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n581_), .A2(new_n364_), .A3(new_n263_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(new_n569_), .A3(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(new_n548_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(new_n219_), .ZN(G1344gat));
  NOR2_X1   g614(.A1(new_n813_), .A2(new_n667_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(new_n220_), .ZN(G1345gat));
  NOR2_X1   g616(.A1(new_n813_), .A2(new_n591_), .ZN(new_n818_));
  XOR2_X1   g617(.A(KEYINPUT61), .B(G155gat), .Z(new_n819_));
  XNOR2_X1  g618(.A(new_n818_), .B(new_n819_), .ZN(G1346gat));
  INV_X1    g619(.A(G162gat), .ZN(new_n821_));
  INV_X1    g620(.A(new_n461_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n813_), .B2(new_n822_), .ZN(new_n823_));
  XOR2_X1   g622(.A(new_n823_), .B(KEYINPUT120), .Z(new_n824_));
  NAND2_X1  g623(.A1(new_n560_), .A2(G162gat), .ZN(new_n825_));
  XOR2_X1   g624(.A(new_n825_), .B(KEYINPUT121), .Z(new_n826_));
  NOR2_X1   g625(.A1(new_n813_), .A2(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n824_), .A2(new_n827_), .ZN(G1347gat));
  INV_X1    g627(.A(KEYINPUT122), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n767_), .A2(new_n264_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n570_), .A2(new_n366_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n830_), .A2(new_n547_), .A3(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n829_), .B1(new_n833_), .B2(G169gat), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT62), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n833_), .A2(new_n829_), .A3(G169gat), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n834_), .A2(new_n835_), .ZN(new_n839_));
  XOR2_X1   g638(.A(KEYINPUT22), .B(G169gat), .Z(new_n840_));
  OAI211_X1 g639(.A(new_n838_), .B(new_n839_), .C1(new_n833_), .C2(new_n840_), .ZN(G1348gat));
  NAND2_X1  g640(.A1(new_n830_), .A2(new_n832_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(G176gat), .B1(new_n843_), .B2(new_n530_), .ZN(new_n844_));
  XOR2_X1   g643(.A(new_n830_), .B(KEYINPUT123), .Z(new_n845_));
  AND3_X1   g644(.A1(new_n832_), .A2(G176gat), .A3(new_n530_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n844_), .B1(new_n845_), .B2(new_n846_), .ZN(G1349gat));
  AND3_X1   g646(.A1(new_n843_), .A2(new_n287_), .A3(new_n497_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n845_), .A2(new_n497_), .A3(new_n832_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n267_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n848_), .B1(new_n849_), .B2(new_n850_), .ZN(G1350gat));
  OAI21_X1  g650(.A(G190gat), .B1(new_n842_), .B2(new_n599_), .ZN(new_n852_));
  OR2_X1    g651(.A1(new_n822_), .A2(new_n280_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n842_), .B2(new_n853_), .ZN(G1351gat));
  INV_X1    g653(.A(KEYINPUT125), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n345_), .A2(new_n364_), .A3(new_n264_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(KEYINPUT124), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n569_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n855_), .B1(new_n767_), .B2(new_n859_), .ZN(new_n860_));
  OAI211_X1 g659(.A(KEYINPUT125), .B(new_n858_), .C1(new_n778_), .C2(new_n718_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n547_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n530_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g665(.A(new_n591_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n862_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(KEYINPUT126), .ZN(new_n869_));
  NOR2_X1   g668(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT126), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n862_), .A2(new_n871_), .A3(new_n867_), .ZN(new_n872_));
  AND3_X1   g671(.A1(new_n869_), .A2(new_n870_), .A3(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n870_), .B1(new_n869_), .B2(new_n872_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1354gat));
  NAND2_X1  g674(.A1(new_n862_), .A2(new_n461_), .ZN(new_n876_));
  XOR2_X1   g675(.A(KEYINPUT127), .B(G218gat), .Z(new_n877_));
  NOR2_X1   g676(.A1(new_n599_), .A2(new_n877_), .ZN(new_n878_));
  AOI22_X1  g677(.A1(new_n876_), .A2(new_n877_), .B1(new_n862_), .B2(new_n878_), .ZN(G1355gat));
endmodule


