//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 0 1 0 0 0 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n626_, new_n627_, new_n628_, new_n629_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n866_, new_n868_, new_n869_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n904_, new_n905_,
    new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n915_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  NOR2_X1   g001(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G169gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G183gat), .A2(G190gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT81), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n205_), .A2(KEYINPUT23), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  AOI21_X1  g012(.A(KEYINPUT92), .B1(new_n211_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT92), .ZN(new_n215_));
  AOI211_X1 g014(.A(new_n215_), .B(new_n212_), .C1(new_n209_), .C2(new_n210_), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n204_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n205_), .A2(new_n208_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n205_), .B(KEYINPUT81), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n218_), .B1(new_n219_), .B2(new_n208_), .ZN(new_n220_));
  NOR3_X1   g019(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT25), .B(G183gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT26), .B(G190gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  AND3_X1   g028(.A1(new_n225_), .A2(new_n229_), .A3(KEYINPUT90), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT90), .B1(new_n225_), .B2(new_n229_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n222_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT91), .ZN(new_n233_));
  XOR2_X1   g032(.A(G197gat), .B(G204gat), .Z(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT21), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G211gat), .B(G218gat), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G197gat), .B(G204gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT21), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n235_), .A2(new_n240_), .A3(new_n236_), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n237_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT91), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n222_), .B(new_n243_), .C1(new_n230_), .C2(new_n231_), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n217_), .A2(new_n233_), .A3(new_n242_), .A4(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G226gat), .A2(G233gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT19), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT20), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT79), .ZN(new_n250_));
  INV_X1    g049(.A(G183gat), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n250_), .B1(new_n251_), .B2(KEYINPUT25), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n224_), .B(new_n252_), .C1(new_n223_), .C2(new_n250_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT80), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n221_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(new_n254_), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n255_), .A2(new_n211_), .A3(new_n256_), .A4(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n204_), .B1(new_n220_), .B2(new_n212_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n242_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n249_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  AND3_X1   g061(.A1(new_n245_), .A2(new_n248_), .A3(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n217_), .A2(new_n233_), .A3(new_n244_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(new_n261_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n258_), .A2(new_n242_), .A3(new_n259_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT20), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT89), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n266_), .A2(KEYINPUT89), .A3(KEYINPUT20), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n265_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n263_), .B1(new_n271_), .B2(new_n247_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G8gat), .B(G36gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT18), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G64gat), .B(G92gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n272_), .A2(new_n277_), .ZN(new_n278_));
  AOI22_X1  g077(.A1(new_n261_), .A2(new_n264_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n248_), .B1(new_n279_), .B2(new_n270_), .ZN(new_n280_));
  NOR3_X1   g079(.A1(new_n280_), .A2(new_n276_), .A3(new_n263_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n202_), .B1(new_n278_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n272_), .A2(new_n277_), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n265_), .A2(new_n269_), .A3(new_n248_), .A4(new_n270_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n217_), .A2(new_n242_), .A3(new_n232_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n262_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(new_n247_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n284_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n276_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n283_), .A2(KEYINPUT27), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n282_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G78gat), .B(G106gat), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(G155gat), .A2(G162gat), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G155gat), .A2(G162gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NOR3_X1   g096(.A1(KEYINPUT86), .A2(G141gat), .A3(G148gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT3), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G141gat), .A2(G148gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT87), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT2), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n297_), .B1(new_n299_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n296_), .A2(KEYINPUT84), .A3(KEYINPUT1), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT84), .B1(new_n296_), .B2(KEYINPUT1), .ZN(new_n307_));
  OAI221_X1 g106(.A(new_n295_), .B1(KEYINPUT1), .B2(new_n296_), .C1(new_n306_), .C2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT85), .ZN(new_n309_));
  XOR2_X1   g108(.A(G141gat), .B(G148gat), .Z(new_n310_));
  NAND3_X1  g109(.A1(new_n308_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n309_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n305_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT29), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n261_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(G228gat), .A3(G233gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G228gat), .A2(G233gat), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n315_), .A2(new_n318_), .A3(new_n261_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n293_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n317_), .A2(new_n319_), .A3(new_n293_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n314_), .A2(KEYINPUT29), .ZN(new_n324_));
  XOR2_X1   g123(.A(G22gat), .B(G50gat), .Z(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT28), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n324_), .B(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n327_), .B1(new_n320_), .B2(KEYINPUT88), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n323_), .A2(new_n328_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n321_), .A2(KEYINPUT88), .A3(new_n322_), .A4(new_n327_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G127gat), .B(G134gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G113gat), .B(G120gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n334_), .B(new_n305_), .C1(new_n312_), .C2(new_n313_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n313_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n304_), .B1(new_n336_), .B2(new_n311_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n334_), .A2(KEYINPUT83), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT83), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n339_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n335_), .B(KEYINPUT4), .C1(new_n337_), .C2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n341_), .ZN(new_n343_));
  XOR2_X1   g142(.A(KEYINPUT93), .B(KEYINPUT4), .Z(new_n344_));
  NAND3_X1  g143(.A1(new_n314_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n342_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G225gat), .A2(G233gat), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G1gat), .B(G29gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(G85gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT0), .B(G57gat), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n351_), .B(new_n352_), .Z(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n314_), .A2(new_n343_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n348_), .B1(new_n355_), .B2(new_n335_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n349_), .A2(new_n354_), .A3(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n347_), .B1(new_n342_), .B2(new_n345_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n353_), .B1(new_n359_), .B2(new_n356_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G227gat), .A2(G233gat), .ZN(new_n362_));
  INV_X1    g161(.A(G15gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT30), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n260_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT82), .B(G43gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n341_), .B(KEYINPUT31), .ZN(new_n369_));
  XOR2_X1   g168(.A(G71gat), .B(G99gat), .Z(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n368_), .B(new_n371_), .ZN(new_n372_));
  NOR4_X1   g171(.A1(new_n291_), .A2(new_n331_), .A3(new_n361_), .A4(new_n372_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n282_), .A2(new_n290_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n361_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n276_), .B1(new_n280_), .B2(new_n263_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n355_), .A2(new_n348_), .A3(new_n335_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n354_), .B(new_n378_), .C1(new_n346_), .C2(new_n348_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n377_), .A2(new_n283_), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT33), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n360_), .A2(new_n381_), .ZN(new_n382_));
  OAI211_X1 g181(.A(KEYINPUT33), .B(new_n353_), .C1(new_n359_), .C2(new_n356_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n380_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT95), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n277_), .A2(KEYINPUT32), .ZN(new_n387_));
  XOR2_X1   g186(.A(new_n387_), .B(KEYINPUT94), .Z(new_n388_));
  NAND2_X1  g187(.A1(new_n272_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n288_), .A2(new_n387_), .ZN(new_n390_));
  AND4_X1   g189(.A1(new_n386_), .A2(new_n389_), .A3(new_n361_), .A4(new_n390_), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n272_), .A2(new_n388_), .B1(new_n288_), .B2(new_n387_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n386_), .B1(new_n392_), .B2(new_n361_), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n385_), .A2(new_n391_), .A3(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n376_), .B1(new_n394_), .B2(new_n331_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n373_), .B1(new_n395_), .B2(new_n372_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT13), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G57gat), .B(G64gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT11), .ZN(new_n399_));
  XOR2_X1   g198(.A(G71gat), .B(G78gat), .Z(new_n400_));
  OR2_X1    g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n398_), .A2(KEYINPUT11), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n399_), .A2(new_n400_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n401_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  XOR2_X1   g203(.A(KEYINPUT10), .B(G99gat), .Z(new_n405_));
  XOR2_X1   g204(.A(KEYINPUT64), .B(G106gat), .Z(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G99gat), .A2(G106gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT6), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT6), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n410_), .A2(G99gat), .A3(G106gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT9), .ZN(new_n413_));
  INV_X1    g212(.A(G85gat), .ZN(new_n414_));
  INV_X1    g213(.A(G92gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G85gat), .A2(G92gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n413_), .B(new_n416_), .C1(new_n418_), .C2(KEYINPUT65), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT65), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n416_), .A2(new_n420_), .A3(KEYINPUT9), .A4(new_n417_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n407_), .A2(new_n412_), .A3(new_n419_), .A4(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT66), .B1(G99gat), .B2(G106gat), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT7), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NOR3_X1   g224(.A1(KEYINPUT66), .A2(G99gat), .A3(G106gat), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT67), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT66), .ZN(new_n428_));
  INV_X1    g227(.A(G99gat), .ZN(new_n429_));
  INV_X1    g228(.A(G106gat), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT67), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n431_), .A2(new_n432_), .A3(new_n424_), .A4(new_n423_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n429_), .A2(new_n430_), .ZN(new_n434_));
  AOI22_X1  g233(.A1(new_n409_), .A2(new_n411_), .B1(new_n434_), .B2(KEYINPUT7), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n427_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT8), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n416_), .A2(new_n417_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n437_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n404_), .B(new_n422_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT68), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n436_), .A2(new_n438_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT8), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n447_), .A2(KEYINPUT68), .A3(new_n404_), .A4(new_n422_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n422_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n404_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n443_), .A2(new_n448_), .A3(new_n451_), .ZN(new_n452_));
  AND2_X1   g251(.A1(G230gat), .A2(G233gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  XOR2_X1   g253(.A(KEYINPUT70), .B(KEYINPUT12), .Z(new_n455_));
  INV_X1    g254(.A(new_n422_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n456_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n455_), .B1(new_n457_), .B2(new_n404_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n453_), .B1(new_n457_), .B2(new_n404_), .ZN(new_n459_));
  OR2_X1    g258(.A1(new_n403_), .A2(new_n402_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(KEYINPUT12), .A3(new_n401_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n439_), .A2(new_n440_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n422_), .B(KEYINPUT69), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n462_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n458_), .A2(new_n459_), .A3(new_n465_), .ZN(new_n466_));
  XOR2_X1   g265(.A(G120gat), .B(G148gat), .Z(new_n467_));
  XNOR2_X1  g266(.A(G176gat), .B(G204gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n470_));
  XOR2_X1   g269(.A(new_n469_), .B(new_n470_), .Z(new_n471_));
  AND3_X1   g270(.A1(new_n454_), .A2(new_n466_), .A3(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n471_), .B1(new_n454_), .B2(new_n466_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n397_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n454_), .A2(new_n466_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n471_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n454_), .A2(new_n466_), .A3(new_n471_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(KEYINPUT13), .A3(new_n478_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n474_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G113gat), .B(G141gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G169gat), .B(G197gat), .ZN(new_n482_));
  XOR2_X1   g281(.A(new_n481_), .B(new_n482_), .Z(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(KEYINPUT75), .B(G8gat), .Z(new_n485_));
  INV_X1    g284(.A(G1gat), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT14), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G15gat), .B(G22gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G1gat), .B(G8gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G29gat), .B(G36gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G43gat), .B(G50gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT15), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n491_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n490_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n489_), .B(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n494_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G229gat), .A2(G233gat), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n496_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n494_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n491_), .A2(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n500_), .B1(new_n504_), .B2(new_n499_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n484_), .B1(new_n502_), .B2(new_n505_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n499_), .A2(new_n504_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n501_), .B(new_n483_), .C1(new_n507_), .C2(new_n500_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n480_), .A2(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n396_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT74), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G232gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT34), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT35), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  OAI22_X1  g316(.A1(new_n449_), .A2(new_n503_), .B1(KEYINPUT35), .B2(new_n514_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT15), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n494_), .B(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT69), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n422_), .B(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n520_), .B1(new_n522_), .B2(new_n447_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n517_), .B1(new_n518_), .B2(new_n523_), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n457_), .A2(new_n494_), .B1(new_n516_), .B2(new_n515_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n517_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n495_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(G190gat), .B(G218gat), .Z(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT72), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G134gat), .B(G162gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT73), .B(KEYINPUT36), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n524_), .A2(new_n528_), .A3(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n532_), .B(KEYINPUT36), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n536_), .B1(new_n524_), .B2(new_n528_), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n512_), .B(KEYINPUT37), .C1(new_n535_), .C2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n524_), .A2(new_n528_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n536_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n524_), .A2(new_n528_), .A3(new_n534_), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n512_), .A2(KEYINPUT37), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n512_), .A2(KEYINPUT37), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .A4(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n538_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G231gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n404_), .B(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(new_n498_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n450_), .A2(new_n547_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n460_), .A2(new_n547_), .A3(new_n401_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n491_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G183gat), .B(G211gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G127gat), .B(G155gat), .Z(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n558_), .A2(new_n559_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n555_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n562_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n564_), .A2(new_n554_), .A3(new_n560_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  AOI22_X1  g365(.A1(new_n549_), .A2(new_n553_), .B1(new_n566_), .B2(KEYINPUT17), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(KEYINPUT17), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n549_), .A2(new_n553_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n567_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n546_), .A2(new_n570_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n511_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n361_), .B(KEYINPUT96), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n572_), .A2(new_n486_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT38), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n535_), .A2(new_n537_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT98), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n396_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n510_), .A2(KEYINPUT97), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n474_), .A2(new_n479_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n509_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT97), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n570_), .B1(new_n582_), .B2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n581_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n361_), .ZN(new_n590_));
  OAI21_X1  g389(.A(G1gat), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n575_), .A2(new_n576_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n577_), .A2(new_n591_), .A3(new_n592_), .ZN(G1324gat));
  NAND3_X1  g392(.A1(new_n572_), .A2(new_n485_), .A3(new_n291_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n373_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n389_), .A2(new_n361_), .A3(new_n390_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT95), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n392_), .A2(new_n386_), .A3(new_n361_), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n597_), .B(new_n598_), .C1(new_n380_), .C2(new_n384_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n331_), .ZN(new_n600_));
  AOI22_X1  g399(.A1(new_n599_), .A2(new_n600_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n372_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n595_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  AND4_X1   g402(.A1(new_n291_), .A2(new_n603_), .A3(new_n579_), .A4(new_n588_), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n604_), .A2(KEYINPUT99), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT39), .ZN(new_n606_));
  INV_X1    g405(.A(G8gat), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n607_), .B1(new_n604_), .B2(KEYINPUT99), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n605_), .A2(new_n606_), .A3(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n606_), .B1(new_n605_), .B2(new_n608_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n594_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT40), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  OAI211_X1 g412(.A(KEYINPUT40), .B(new_n594_), .C1(new_n609_), .C2(new_n610_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(G1325gat));
  NAND3_X1  g414(.A1(new_n572_), .A2(new_n363_), .A3(new_n602_), .ZN(new_n616_));
  OAI21_X1  g415(.A(G15gat), .B1(new_n589_), .B2(new_n372_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT41), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n617_), .A2(new_n618_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n616_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT100), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  OAI211_X1 g422(.A(KEYINPUT100), .B(new_n616_), .C1(new_n619_), .C2(new_n620_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1326gat));
  OAI21_X1  g424(.A(G22gat), .B1(new_n589_), .B2(new_n600_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT42), .ZN(new_n627_));
  INV_X1    g426(.A(G22gat), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n572_), .A2(new_n628_), .A3(new_n331_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(G1327gat));
  INV_X1    g429(.A(new_n570_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n578_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n603_), .A2(new_n585_), .A3(new_n632_), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n633_), .A2(KEYINPUT102), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(KEYINPUT102), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(G29gat), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(new_n637_), .A3(new_n361_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT43), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n538_), .A2(new_n545_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n639_), .B1(new_n396_), .B2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n582_), .A2(new_n587_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n603_), .A2(KEYINPUT43), .A3(new_n546_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n641_), .A2(new_n570_), .A3(new_n642_), .A4(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT44), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n603_), .A2(new_n546_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n631_), .B1(new_n647_), .B2(new_n639_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n648_), .A2(KEYINPUT44), .A3(new_n642_), .A4(new_n643_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n646_), .A2(new_n649_), .A3(new_n574_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n650_), .A2(KEYINPUT101), .ZN(new_n651_));
  OAI21_X1  g450(.A(G29gat), .B1(new_n650_), .B2(KEYINPUT101), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n638_), .B1(new_n651_), .B2(new_n652_), .ZN(G1328gat));
  NAND3_X1  g452(.A1(new_n646_), .A2(new_n649_), .A3(new_n291_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(G36gat), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n374_), .A2(G36gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n634_), .A2(new_n635_), .A3(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT45), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT45), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n634_), .A2(new_n659_), .A3(new_n635_), .A4(new_n656_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n655_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT46), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n655_), .A2(new_n661_), .A3(KEYINPUT46), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1329gat));
  NAND4_X1  g465(.A1(new_n646_), .A2(new_n649_), .A3(G43gat), .A4(new_n602_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n634_), .A2(new_n602_), .A3(new_n635_), .ZN(new_n668_));
  INV_X1    g467(.A(G43gat), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n667_), .A2(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g471(.A(G50gat), .B1(new_n636_), .B2(new_n331_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n646_), .A2(new_n649_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n331_), .A2(G50gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n673_), .B1(new_n674_), .B2(new_n675_), .ZN(G1331gat));
  NOR2_X1   g475(.A1(new_n509_), .A2(new_n570_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n583_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n581_), .A2(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(G57gat), .B1(new_n679_), .B2(new_n590_), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n396_), .A2(KEYINPUT103), .A3(new_n509_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n603_), .B2(new_n584_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n681_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(new_n571_), .A3(new_n583_), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n573_), .A2(G57gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n680_), .B1(new_n685_), .B2(new_n686_), .ZN(G1332gat));
  NOR3_X1   g486(.A1(new_n685_), .A2(G64gat), .A3(new_n374_), .ZN(new_n688_));
  OAI21_X1  g487(.A(G64gat), .B1(new_n679_), .B2(new_n374_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(KEYINPUT104), .B(KEYINPUT48), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n688_), .A2(new_n691_), .ZN(G1333gat));
  OR2_X1    g491(.A1(new_n372_), .A2(G71gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n581_), .A2(new_n602_), .A3(new_n678_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT49), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n694_), .A2(new_n695_), .A3(G71gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n694_), .B2(G71gat), .ZN(new_n697_));
  OAI22_X1  g496(.A1(new_n685_), .A2(new_n693_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT105), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n698_), .B(new_n699_), .ZN(G1334gat));
  OAI21_X1  g499(.A(G78gat), .B1(new_n679_), .B2(new_n600_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT50), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n600_), .A2(G78gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n685_), .B2(new_n703_), .ZN(G1335gat));
  NOR2_X1   g503(.A1(new_n480_), .A2(new_n509_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n648_), .A2(new_n643_), .A3(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(G85gat), .B1(new_n706_), .B2(new_n590_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n583_), .B(new_n632_), .C1(new_n681_), .C2(new_n683_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n708_), .A2(KEYINPUT106), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n708_), .A2(KEYINPUT106), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n574_), .A2(new_n414_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n707_), .B1(new_n711_), .B2(new_n712_), .ZN(G1336gat));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n648_), .A2(new_n291_), .A3(new_n643_), .A4(new_n705_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(G92gat), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n291_), .A2(new_n415_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n714_), .B(new_n716_), .C1(new_n711_), .C2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n684_), .A2(new_n719_), .A3(new_n583_), .A4(new_n632_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n708_), .A2(KEYINPUT106), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n716_), .ZN(new_n723_));
  OAI21_X1  g522(.A(KEYINPUT107), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n718_), .A2(new_n724_), .ZN(G1337gat));
  INV_X1    g524(.A(KEYINPUT51), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n648_), .A2(new_n602_), .A3(new_n643_), .A4(new_n705_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(G99gat), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n602_), .A2(new_n405_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n726_), .B(new_n728_), .C1(new_n711_), .C2(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n728_), .ZN(new_n732_));
  OAI21_X1  g531(.A(KEYINPUT51), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n730_), .A2(new_n733_), .ZN(G1338gat));
  NAND4_X1  g533(.A1(new_n648_), .A2(new_n331_), .A3(new_n643_), .A4(new_n705_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT52), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n735_), .A2(new_n736_), .A3(G106gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n735_), .B2(G106gat), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n331_), .A2(new_n406_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n741_));
  OAI21_X1  g540(.A(KEYINPUT53), .B1(new_n739_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n740_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n743_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT53), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n744_), .B(new_n745_), .C1(new_n738_), .C2(new_n737_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n742_), .A2(new_n746_), .ZN(G1339gat));
  INV_X1    g546(.A(KEYINPUT114), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n480_), .A2(new_n640_), .A3(new_n677_), .ZN(new_n749_));
  AOI21_X1  g548(.A(KEYINPUT109), .B1(new_n749_), .B2(KEYINPUT54), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n474_), .A2(new_n479_), .A3(new_n677_), .ZN(new_n751_));
  OAI211_X1 g550(.A(KEYINPUT109), .B(KEYINPUT54), .C1(new_n751_), .C2(new_n546_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n751_), .A2(new_n546_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT54), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT108), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT108), .ZN(new_n757_));
  NOR4_X1   g556(.A1(new_n751_), .A2(new_n546_), .A3(new_n757_), .A4(KEYINPUT54), .ZN(new_n758_));
  OAI22_X1  g557(.A1(new_n750_), .A2(new_n753_), .B1(new_n756_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n480_), .A2(new_n640_), .A3(new_n755_), .A4(new_n677_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n757_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n754_), .A2(KEYINPUT108), .A3(new_n755_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(KEYINPUT54), .B1(new_n751_), .B2(new_n546_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n752_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n765_), .A2(new_n769_), .A3(KEYINPUT110), .ZN(new_n770_));
  INV_X1    g569(.A(new_n500_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n496_), .A2(new_n499_), .A3(new_n771_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n484_), .B(new_n772_), .C1(new_n507_), .C2(new_n771_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n508_), .A2(new_n773_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n472_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n466_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n458_), .A2(new_n465_), .A3(new_n441_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n453_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n458_), .A2(new_n459_), .A3(KEYINPUT55), .A4(new_n465_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n777_), .A2(new_n779_), .A3(new_n780_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n781_), .A2(KEYINPUT56), .A3(new_n476_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT56), .B1(new_n781_), .B2(new_n476_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n775_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT58), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n640_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n781_), .A2(new_n476_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT56), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n781_), .A2(KEYINPUT56), .A3(new_n476_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n791_), .A2(new_n792_), .A3(KEYINPUT58), .A4(new_n775_), .ZN(new_n793_));
  OAI211_X1 g592(.A(KEYINPUT58), .B(new_n775_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT113), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n786_), .A2(new_n793_), .A3(new_n795_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n578_), .A2(KEYINPUT57), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n584_), .A2(new_n472_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n800_), .B1(KEYINPUT111), .B2(new_n788_), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n781_), .A2(new_n476_), .A3(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n788_), .A2(KEYINPUT111), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n803_), .B1(new_n781_), .B2(new_n476_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n802_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n790_), .A2(new_n800_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n799_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n472_), .A2(new_n473_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n808_), .A2(new_n774_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n797_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n578_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n781_), .A2(new_n476_), .A3(new_n801_), .ZN(new_n812_));
  AOI22_X1  g611(.A1(new_n776_), .A2(new_n466_), .B1(new_n778_), .B2(new_n453_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n471_), .B1(new_n813_), .B2(new_n780_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n812_), .B1(new_n814_), .B2(new_n803_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT112), .B1(new_n814_), .B2(KEYINPUT56), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n798_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n809_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n811_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n796_), .B(new_n810_), .C1(new_n819_), .C2(KEYINPUT57), .ZN(new_n820_));
  AOI22_X1  g619(.A1(new_n761_), .A2(new_n770_), .B1(new_n570_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT59), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n291_), .A2(new_n331_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n823_), .A2(new_n602_), .A3(new_n574_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n821_), .A2(new_n822_), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n820_), .A2(new_n570_), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n765_), .A2(KEYINPUT110), .A3(new_n769_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT110), .B1(new_n765_), .B2(new_n769_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n826_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n824_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT59), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n748_), .B1(new_n825_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n822_), .B1(new_n821_), .B2(new_n824_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n829_), .A2(KEYINPUT59), .A3(new_n830_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(KEYINPUT114), .A3(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n509_), .A2(new_n836_), .A3(G113gat), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(new_n836_), .B2(G113gat), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n832_), .A2(new_n835_), .A3(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(G113gat), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n821_), .A2(new_n824_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n840_), .B1(new_n842_), .B2(new_n584_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n839_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT116), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n839_), .A2(new_n846_), .A3(new_n843_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(G1340gat));
  INV_X1    g647(.A(G120gat), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n480_), .B2(KEYINPUT60), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n841_), .B(new_n850_), .C1(KEYINPUT60), .C2(new_n849_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n480_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n852_), .B2(new_n849_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT117), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n853_), .B(new_n854_), .ZN(G1341gat));
  NAND3_X1  g654(.A1(new_n832_), .A2(new_n631_), .A3(new_n835_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(G127gat), .ZN(new_n857_));
  OR2_X1    g656(.A1(new_n570_), .A2(G127gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n842_), .B2(new_n858_), .ZN(G1342gat));
  XNOR2_X1  g658(.A(KEYINPUT118), .B(G134gat), .ZN(new_n860_));
  AND4_X1   g659(.A1(new_n546_), .A2(new_n832_), .A3(new_n835_), .A4(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(G134gat), .B1(new_n841_), .B2(new_n580_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1343gat));
  NAND4_X1  g662(.A1(new_n374_), .A2(new_n574_), .A3(new_n331_), .A4(new_n372_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n821_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n509_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n583_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(KEYINPUT119), .B(G148gat), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n868_), .B(new_n869_), .ZN(G1345gat));
  NAND2_X1  g669(.A1(new_n865_), .A2(new_n631_), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n871_), .A2(KEYINPUT120), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(KEYINPUT120), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT61), .B(G155gat), .ZN(new_n874_));
  AND3_X1   g673(.A1(new_n872_), .A2(new_n873_), .A3(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1346gat));
  INV_X1    g676(.A(G162gat), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n865_), .A2(new_n878_), .A3(new_n580_), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n821_), .A2(new_n640_), .A3(new_n864_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n878_), .B2(new_n880_), .ZN(G1347gat));
  NAND3_X1  g680(.A1(new_n600_), .A2(new_n291_), .A3(new_n602_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n821_), .A2(new_n574_), .A3(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n509_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n883_), .A2(KEYINPUT121), .A3(new_n509_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n886_), .A2(G169gat), .A3(new_n887_), .ZN(new_n888_));
  AND2_X1   g687(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n889_));
  NOR2_X1   g688(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n888_), .A2(new_n891_), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n886_), .A2(G169gat), .A3(new_n887_), .A4(new_n889_), .ZN(new_n893_));
  XOR2_X1   g692(.A(KEYINPUT22), .B(G169gat), .Z(new_n894_));
  NOR2_X1   g693(.A1(new_n584_), .A2(new_n894_), .ZN(new_n895_));
  XOR2_X1   g694(.A(new_n895_), .B(KEYINPUT123), .Z(new_n896_));
  NAND2_X1  g695(.A1(new_n883_), .A2(new_n896_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n892_), .A2(new_n893_), .A3(new_n897_), .ZN(G1348gat));
  AND2_X1   g697(.A1(KEYINPUT124), .A2(G176gat), .ZN(new_n899_));
  NOR2_X1   g698(.A1(KEYINPUT124), .A2(G176gat), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n883_), .A2(new_n583_), .ZN(new_n902_));
  MUX2_X1   g701(.A(new_n901_), .B(new_n899_), .S(new_n902_), .Z(G1349gat));
  NAND2_X1  g702(.A1(new_n883_), .A2(new_n631_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n223_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n905_), .B1(new_n251_), .B2(new_n904_), .ZN(G1350gat));
  NAND2_X1  g705(.A1(new_n883_), .A2(new_n546_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(G190gat), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT125), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n883_), .A2(new_n224_), .A3(new_n580_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1351gat));
  NAND3_X1  g711(.A1(new_n291_), .A2(new_n375_), .A3(new_n372_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n821_), .A2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(new_n509_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n583_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g717(.A1(new_n914_), .A2(new_n631_), .ZN(new_n919_));
  OR2_X1    g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  XOR2_X1   g720(.A(KEYINPUT63), .B(G211gat), .Z(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n919_), .B2(new_n922_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(KEYINPUT126), .ZN(G1354gat));
  AOI21_X1  g723(.A(G218gat), .B1(new_n914_), .B2(new_n580_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n546_), .A2(G218gat), .ZN(new_n926_));
  XOR2_X1   g725(.A(new_n926_), .B(KEYINPUT127), .Z(new_n927_));
  AOI21_X1  g726(.A(new_n925_), .B1(new_n914_), .B2(new_n927_), .ZN(G1355gat));
endmodule


