//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 1 0 0 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n839_, new_n840_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n849_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n876_,
    new_n877_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_;
  XNOR2_X1  g000(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n202_));
  AND2_X1   g001(.A1(KEYINPUT77), .A2(KEYINPUT22), .ZN(new_n203_));
  OAI21_X1  g002(.A(G169gat), .B1(new_n203_), .B2(G176gat), .ZN(new_n204_));
  INV_X1    g003(.A(G169gat), .ZN(new_n205_));
  INV_X1    g004(.A(G176gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT23), .ZN(new_n209_));
  INV_X1    g008(.A(G183gat), .ZN(new_n210_));
  INV_X1    g009(.A(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  AND3_X1   g011(.A1(new_n209_), .A2(KEYINPUT78), .A3(new_n212_), .ZN(new_n213_));
  AOI21_X1  g012(.A(KEYINPUT78), .B1(new_n209_), .B2(new_n212_), .ZN(new_n214_));
  OAI221_X1 g013(.A(new_n204_), .B1(new_n203_), .B2(new_n207_), .C1(new_n213_), .C2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT30), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT25), .B(G183gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT26), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT75), .B1(new_n218_), .B2(G190gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT26), .B(G190gat), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n217_), .B(new_n219_), .C1(new_n220_), .C2(KEYINPUT75), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n221_), .A2(KEYINPUT76), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n207_), .A2(KEYINPUT24), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n207_), .A2(KEYINPUT24), .A3(new_n224_), .ZN(new_n225_));
  AND3_X1   g024(.A1(new_n209_), .A2(new_n223_), .A3(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n221_), .A2(KEYINPUT76), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n222_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n215_), .A2(new_n216_), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n216_), .B1(new_n215_), .B2(new_n228_), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT79), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G127gat), .B(G134gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G113gat), .B(G120gat), .ZN(new_n234_));
  XOR2_X1   g033(.A(new_n233_), .B(new_n234_), .Z(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT80), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT80), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n233_), .A2(new_n234_), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G15gat), .B(G43gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G227gat), .A2(G233gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G71gat), .B(G99gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n232_), .A2(new_n239_), .A3(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n239_), .B1(new_n232_), .B2(new_n244_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n202_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT79), .ZN(new_n248_));
  INV_X1    g047(.A(new_n231_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n248_), .B1(new_n249_), .B2(new_n229_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n244_), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n238_), .B(new_n236_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n202_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n232_), .A2(new_n239_), .A3(new_n244_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  NOR3_X1   g054(.A1(new_n230_), .A2(new_n231_), .A3(KEYINPUT79), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n247_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n256_), .B1(new_n247_), .B2(new_n255_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G211gat), .B(G218gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT88), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT21), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  OR2_X1    g063(.A1(new_n261_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n261_), .A2(new_n264_), .ZN(new_n266_));
  INV_X1    g065(.A(G197gat), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n267_), .A2(G204gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT87), .B(G204gat), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n269_), .A2(new_n267_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n265_), .B(new_n266_), .C1(new_n268_), .C2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n267_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n267_), .A2(G204gat), .ZN(new_n273_));
  OR2_X1    g072(.A1(new_n273_), .A2(KEYINPUT86), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n263_), .B1(new_n273_), .B2(KEYINPUT86), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n272_), .A2(new_n274_), .A3(new_n261_), .A4(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n271_), .A2(new_n276_), .ZN(new_n277_));
  AND2_X1   g076(.A1(G155gat), .A2(G162gat), .ZN(new_n278_));
  NOR2_X1   g077(.A1(G155gat), .A2(G162gat), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT1), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  OR2_X1    g081(.A1(G141gat), .A2(G148gat), .ZN(new_n283_));
  AOI22_X1  g082(.A1(new_n278_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT82), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n282_), .A2(KEYINPUT82), .A3(new_n283_), .A4(new_n284_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT2), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n283_), .A2(KEYINPUT3), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n283_), .A2(KEYINPUT3), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  AOI22_X1  g092(.A1(new_n287_), .A2(new_n288_), .B1(new_n280_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT29), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n277_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G78gat), .B(G106gat), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n277_), .B(new_n297_), .C1(new_n294_), .C2(new_n295_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n277_), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n302_), .A2(KEYINPUT84), .ZN(new_n303_));
  XOR2_X1   g102(.A(KEYINPUT85), .B(G233gat), .Z(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(G228gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n301_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT83), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n299_), .A2(new_n303_), .A3(new_n305_), .A4(new_n300_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n287_), .A2(new_n288_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n293_), .A2(new_n280_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  OR3_X1    g112(.A1(new_n313_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n314_));
  XOR2_X1   g113(.A(G22gat), .B(G50gat), .Z(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT28), .B1(new_n313_), .B2(KEYINPUT29), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n314_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n315_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n310_), .B(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G225gat), .A2(G233gat), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n313_), .A2(new_n239_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT4), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n235_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n294_), .A2(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n324_), .B1(new_n323_), .B2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n322_), .B1(new_n326_), .B2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n323_), .A2(new_n321_), .A3(new_n328_), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n331_), .A2(KEYINPUT92), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(KEYINPUT92), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n330_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT93), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G1gat), .B(G29gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(G85gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT0), .B(G57gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n335_), .A2(new_n336_), .A3(KEYINPUT33), .A4(new_n341_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n330_), .A2(new_n332_), .A3(new_n333_), .A4(new_n341_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT33), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT93), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n342_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n215_), .A2(new_n228_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n277_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT91), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n224_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT22), .B(G169gat), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT89), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n351_), .B1(new_n354_), .B2(new_n206_), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n209_), .A2(KEYINPUT90), .A3(new_n212_), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT90), .B1(new_n209_), .B2(new_n212_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n217_), .A2(new_n220_), .ZN(new_n359_));
  AOI22_X1  g158(.A1(new_n355_), .A2(new_n358_), .B1(new_n226_), .B2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n302_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n347_), .A2(KEYINPUT91), .A3(new_n277_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n350_), .A2(new_n361_), .A3(KEYINPUT20), .A4(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G226gat), .A2(G233gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT19), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n363_), .A2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT20), .B1(new_n360_), .B2(new_n302_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n302_), .A2(new_n215_), .A3(new_n228_), .ZN(new_n369_));
  NOR3_X1   g168(.A1(new_n368_), .A2(new_n369_), .A3(new_n366_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n367_), .A2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G8gat), .B(G36gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(G92gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT18), .B(G64gat), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n374_), .B(new_n375_), .Z(new_n376_));
  NAND2_X1  g175(.A1(new_n372_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n323_), .A2(new_n328_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT4), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n322_), .B1(new_n379_), .B2(new_n325_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n323_), .A2(new_n322_), .A3(new_n328_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT94), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n381_), .A2(new_n382_), .A3(new_n340_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n382_), .B1(new_n381_), .B2(new_n340_), .ZN(new_n384_));
  NOR3_X1   g183(.A1(new_n380_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n376_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n367_), .A2(new_n371_), .A3(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n377_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n343_), .A2(new_n344_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n346_), .A2(new_n389_), .A3(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n334_), .A2(new_n340_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n343_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT32), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n372_), .B1(new_n395_), .B2(new_n387_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n363_), .A2(new_n365_), .ZN(new_n397_));
  OR3_X1    g196(.A1(new_n368_), .A2(new_n369_), .A3(new_n365_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n399_), .A2(KEYINPUT32), .A3(new_n376_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n394_), .A2(new_n396_), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n260_), .B(new_n320_), .C1(new_n392_), .C2(new_n402_), .ZN(new_n403_));
  XOR2_X1   g202(.A(new_n310_), .B(new_n319_), .Z(new_n404_));
  OAI21_X1  g203(.A(new_n404_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n256_), .ZN(new_n406_));
  NOR3_X1   g205(.A1(new_n245_), .A2(new_n246_), .A3(new_n202_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n253_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n406_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n247_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(new_n320_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n405_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n394_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n399_), .A2(new_n387_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n377_), .A2(new_n414_), .A3(KEYINPUT27), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT27), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n387_), .B1(new_n367_), .B2(new_n371_), .ZN(new_n417_));
  AOI211_X1 g216(.A(new_n376_), .B(new_n370_), .C1(new_n363_), .C2(new_n366_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n416_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n415_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n412_), .A2(new_n413_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n403_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G230gat), .A2(G233gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT7), .ZN(new_n426_));
  INV_X1    g225(.A(G99gat), .ZN(new_n427_));
  INV_X1    g226(.A(G106gat), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n426_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G99gat), .A2(G106gat), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT6), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n429_), .A2(new_n432_), .A3(new_n433_), .A4(new_n434_), .ZN(new_n435_));
  AND2_X1   g234(.A1(G85gat), .A2(G92gat), .ZN(new_n436_));
  NOR2_X1   g235(.A1(G85gat), .A2(G92gat), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n435_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n427_), .A2(KEYINPUT10), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT10), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(G99gat), .ZN(new_n445_));
  AOI21_X1  g244(.A(G106gat), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n432_), .A2(new_n433_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT9), .B1(new_n436_), .B2(new_n437_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT64), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT9), .ZN(new_n451_));
  INV_X1    g250(.A(G85gat), .ZN(new_n452_));
  INV_X1    g251(.A(G92gat), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n451_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n449_), .A2(new_n450_), .A3(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n436_), .A2(KEYINPUT64), .A3(KEYINPUT9), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n448_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n441_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n435_), .A2(new_n438_), .A3(new_n439_), .A4(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n442_), .A2(new_n457_), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(G57gat), .ZN(new_n461_));
  INV_X1    g260(.A(G64gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G57gat), .A2(G64gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT11), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G71gat), .B(G78gat), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT11), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n463_), .A2(new_n469_), .A3(new_n464_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n466_), .A2(new_n468_), .A3(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n465_), .A2(new_n467_), .A3(KEYINPUT11), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n460_), .A2(new_n474_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n473_), .A2(new_n442_), .A3(new_n457_), .A4(new_n459_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n475_), .A2(KEYINPUT12), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT12), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n460_), .A2(new_n478_), .A3(new_n474_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n425_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n424_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G176gat), .B(G204gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G120gat), .B(G148gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT66), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n482_), .B(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n489_), .B(KEYINPUT13), .Z(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  XOR2_X1   g290(.A(G15gat), .B(G22gat), .Z(new_n492_));
  NAND2_X1  g291(.A1(G1gat), .A2(G8gat), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n492_), .B1(KEYINPUT14), .B2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT72), .ZN(new_n495_));
  XOR2_X1   g294(.A(G1gat), .B(G8gat), .Z(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT72), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n494_), .B(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n496_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n497_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G29gat), .B(G36gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G43gat), .B(G50gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  XOR2_X1   g305(.A(G29gat), .B(G36gat), .Z(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(new_n504_), .ZN(new_n508_));
  XOR2_X1   g307(.A(G43gat), .B(G50gat), .Z(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n503_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n497_), .A2(new_n501_), .A3(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n506_), .A2(KEYINPUT74), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G229gat), .A2(G233gat), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT74), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n497_), .A2(new_n501_), .A3(new_n516_), .A4(new_n511_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n513_), .A2(new_n515_), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n505_), .A2(KEYINPUT15), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT15), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n511_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n506_), .B(new_n514_), .C1(new_n502_), .C2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G113gat), .B(G141gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G169gat), .B(G197gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n518_), .A2(new_n524_), .A3(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n528_), .B1(new_n518_), .B2(new_n524_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n491_), .A2(new_n531_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n423_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G231gat), .A2(G233gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n473_), .B(new_n534_), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n502_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G127gat), .B(G155gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(G211gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT16), .B(G183gat), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n538_), .B(new_n539_), .Z(new_n540_));
  INV_X1    g339(.A(KEYINPUT17), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n502_), .A2(new_n535_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n536_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n540_), .A2(new_n541_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n546_), .B1(new_n536_), .B2(new_n543_), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT73), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT73), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n536_), .A2(new_n543_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n549_), .B(new_n544_), .C1(new_n550_), .C2(new_n546_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n548_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT36), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G190gat), .B(G218gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(G162gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(KEYINPUT71), .B(G134gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G232gat), .A2(G233gat), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n558_), .B(KEYINPUT34), .Z(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT68), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n522_), .A2(new_n460_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT69), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n442_), .A2(new_n457_), .A3(new_n505_), .A4(new_n459_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n562_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(new_n563_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n561_), .B1(new_n568_), .B2(KEYINPUT70), .ZN(new_n569_));
  AOI21_X1  g368(.A(KEYINPUT69), .B1(new_n522_), .B2(new_n460_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n566_), .B1(new_n570_), .B2(new_n564_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT70), .ZN(new_n572_));
  NOR3_X1   g371(.A1(new_n571_), .A2(KEYINPUT68), .A3(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n560_), .B1(new_n569_), .B2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n568_), .A2(new_n561_), .A3(KEYINPUT70), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT68), .B1(new_n571_), .B2(new_n572_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n575_), .A2(new_n576_), .A3(new_n559_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT35), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n568_), .A2(new_n578_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n574_), .A2(new_n577_), .A3(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(KEYINPUT35), .B1(new_n574_), .B2(new_n577_), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n553_), .B(new_n557_), .C1(new_n580_), .C2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n574_), .A2(new_n577_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n578_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n557_), .A2(new_n553_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n574_), .A2(new_n577_), .A3(new_n579_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n557_), .A2(new_n553_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n584_), .A2(new_n585_), .A3(new_n586_), .A4(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n582_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT37), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n582_), .A2(new_n588_), .A3(KEYINPUT37), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  AND3_X1   g392(.A1(new_n533_), .A2(new_n552_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(G1gat), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n594_), .A2(new_n595_), .A3(new_n394_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT38), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n545_), .A2(new_n547_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n533_), .A2(new_n599_), .A3(new_n589_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT95), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n601_), .A2(new_n394_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n597_), .B1(new_n602_), .B2(new_n595_), .ZN(G1324gat));
  INV_X1    g402(.A(G8gat), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n604_), .B1(new_n600_), .B2(new_n420_), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n605_), .B(KEYINPUT39), .Z(new_n606_));
  NAND3_X1  g405(.A1(new_n594_), .A2(new_n604_), .A3(new_n420_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g408(.A(G15gat), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n610_), .B1(new_n601_), .B2(new_n259_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT41), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n594_), .A2(new_n610_), .A3(new_n259_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT96), .Z(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(G1326gat));
  INV_X1    g414(.A(G22gat), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n616_), .B1(new_n601_), .B2(new_n404_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT42), .Z(new_n618_));
  NAND3_X1  g417(.A1(new_n594_), .A2(new_n616_), .A3(new_n404_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(G1327gat));
  AND2_X1   g419(.A1(new_n582_), .A2(new_n588_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n552_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT101), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n533_), .A2(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT102), .Z(new_n626_));
  AOI21_X1  g425(.A(G29gat), .B1(new_n626_), .B2(new_n394_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n532_), .A2(new_n622_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT97), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n591_), .A2(new_n592_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT98), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT43), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n423_), .B(new_n630_), .C1(new_n631_), .C2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n630_), .A2(new_n631_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n417_), .A2(new_n418_), .A3(new_n385_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n635_), .A2(new_n390_), .A3(new_n345_), .A4(new_n342_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n259_), .B1(new_n636_), .B2(new_n401_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n420_), .B1(new_n405_), .B2(new_n411_), .ZN(new_n638_));
  AOI22_X1  g437(.A1(new_n637_), .A2(new_n320_), .B1(new_n638_), .B2(new_n413_), .ZN(new_n639_));
  OAI211_X1 g438(.A(KEYINPUT43), .B(new_n634_), .C1(new_n639_), .C2(new_n593_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n629_), .B1(new_n633_), .B2(new_n640_), .ZN(new_n641_));
  OR3_X1    g440(.A1(new_n641_), .A2(KEYINPUT99), .A3(KEYINPUT44), .ZN(new_n642_));
  OAI21_X1  g441(.A(KEYINPUT99), .B1(new_n641_), .B2(KEYINPUT44), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n644_), .A2(G29gat), .A3(new_n394_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n641_), .A2(KEYINPUT44), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n641_), .A2(KEYINPUT100), .A3(KEYINPUT44), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n627_), .B1(new_n645_), .B2(new_n650_), .ZN(G1328gat));
  INV_X1    g450(.A(G36gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n626_), .A2(new_n652_), .A3(new_n420_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT45), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n421_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n652_), .B1(new_n656_), .B2(new_n644_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(KEYINPUT46), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT46), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n660_), .B1(new_n655_), .B2(new_n657_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n661_), .ZN(G1329gat));
  NAND4_X1  g461(.A1(new_n644_), .A2(new_n650_), .A3(G43gat), .A4(new_n259_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(KEYINPUT103), .B(G43gat), .ZN(new_n664_));
  INV_X1    g463(.A(new_n626_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n664_), .B1(new_n665_), .B2(new_n260_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n663_), .A2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g467(.A(G50gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n669_), .B1(new_n665_), .B2(new_n320_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n650_), .A2(G50gat), .A3(new_n404_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n644_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n670_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(G1331gat));
  NAND2_X1  g474(.A1(new_n518_), .A2(new_n524_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(new_n527_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n518_), .A2(new_n524_), .A3(new_n528_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n490_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n639_), .A2(new_n622_), .A3(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n683_), .A2(new_n630_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n413_), .B1(new_n685_), .B2(KEYINPUT105), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n683_), .A2(new_n621_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n413_), .A2(new_n461_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n687_), .B1(KEYINPUT106), .B2(new_n688_), .ZN(new_n689_));
  OAI211_X1 g488(.A(new_n686_), .B(new_n689_), .C1(KEYINPUT105), .C2(new_n685_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G57gat), .B1(new_n689_), .B2(KEYINPUT106), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1332gat));
  AOI21_X1  g491(.A(new_n462_), .B1(new_n687_), .B2(new_n420_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT48), .Z(new_n694_));
  NAND2_X1  g493(.A1(new_n420_), .A2(new_n462_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT107), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n694_), .B1(new_n685_), .B2(new_n696_), .ZN(G1333gat));
  OR3_X1    g496(.A1(new_n685_), .A2(G71gat), .A3(new_n260_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n687_), .ZN(new_n699_));
  OAI21_X1  g498(.A(G71gat), .B1(new_n699_), .B2(new_n260_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT108), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n701_), .A2(KEYINPUT49), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(KEYINPUT49), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n698_), .B1(new_n702_), .B2(new_n703_), .ZN(G1334gat));
  OAI21_X1  g503(.A(G78gat), .B1(new_n699_), .B2(new_n320_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT50), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n320_), .A2(G78gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n706_), .B1(new_n685_), .B2(new_n707_), .ZN(G1335gat));
  AND3_X1   g507(.A1(new_n624_), .A2(new_n423_), .A3(new_n680_), .ZN(new_n709_));
  AOI21_X1  g508(.A(G85gat), .B1(new_n709_), .B2(new_n394_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n681_), .B1(new_n640_), .B2(new_n633_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n711_), .A2(new_n622_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n413_), .A2(new_n452_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n710_), .B1(new_n712_), .B2(new_n713_), .ZN(G1336gat));
  AOI21_X1  g513(.A(new_n453_), .B1(new_n712_), .B2(new_n420_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n421_), .A2(G92gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n709_), .B2(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT109), .ZN(G1337gat));
  AOI21_X1  g517(.A(new_n427_), .B1(new_n712_), .B2(new_n259_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n260_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n709_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT51), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(KEYINPUT110), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(KEYINPUT110), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n723_), .B(new_n724_), .ZN(G1338gat));
  NAND2_X1  g524(.A1(new_n640_), .A2(new_n633_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n726_), .A2(new_n404_), .A3(new_n622_), .A4(new_n680_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT112), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n711_), .A2(KEYINPUT112), .A3(new_n404_), .A4(new_n622_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n729_), .A2(G106gat), .A3(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT113), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT113), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n729_), .A2(new_n733_), .A3(G106gat), .A4(new_n730_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT52), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n732_), .A2(KEYINPUT52), .A3(new_n734_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n709_), .A2(new_n428_), .A3(new_n404_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT111), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n737_), .A2(new_n738_), .A3(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT53), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT53), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n737_), .A2(new_n743_), .A3(new_n738_), .A4(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1339gat));
  INV_X1    g544(.A(KEYINPUT114), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n746_), .B1(new_n622_), .B2(new_n679_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n531_), .A2(KEYINPUT114), .A3(new_n552_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n591_), .A2(new_n749_), .A3(new_n490_), .A4(new_n592_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT54), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n750_), .B(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n477_), .A2(new_n425_), .A3(new_n479_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n480_), .B1(KEYINPUT55), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT55), .ZN(new_n756_));
  AOI211_X1 g555(.A(new_n756_), .B(new_n425_), .C1(new_n477_), .C2(new_n479_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n754_), .A2(new_n755_), .A3(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n755_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(KEYINPUT117), .B1(new_n758_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT117), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n753_), .A2(KEYINPUT55), .ZN(new_n763_));
  OAI21_X1  g562(.A(KEYINPUT116), .B1(new_n763_), .B2(new_n480_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n762_), .B(new_n759_), .C1(new_n764_), .C2(new_n757_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n761_), .A2(new_n487_), .A3(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT56), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT118), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n679_), .B(new_n770_), .C1(new_n482_), .C2(new_n487_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n768_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n761_), .A2(new_n487_), .A3(new_n765_), .A4(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n482_), .A2(new_n487_), .ZN(new_n774_));
  OAI21_X1  g573(.A(KEYINPUT115), .B1(new_n531_), .B2(new_n774_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n769_), .A2(new_n771_), .A3(new_n773_), .A4(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n513_), .A2(new_n514_), .A3(new_n517_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n506_), .B1(new_n502_), .B2(new_n523_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n777_), .B(new_n527_), .C1(new_n514_), .C2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n678_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT119), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT119), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n779_), .A2(new_n782_), .A3(new_n678_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n489_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n776_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n589_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT57), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n761_), .A2(new_n765_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n767_), .A2(KEYINPUT120), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT120), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT56), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n791_), .A2(new_n487_), .A3(new_n792_), .A4(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n774_), .B1(new_n781_), .B2(new_n783_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n766_), .A2(new_n793_), .A3(KEYINPUT56), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n795_), .A2(new_n796_), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT58), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n795_), .A2(KEYINPUT58), .A3(new_n796_), .A4(new_n797_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n800_), .A2(new_n630_), .A3(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n787_), .A2(KEYINPUT57), .A3(new_n589_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n790_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n752_), .B1(new_n804_), .B2(new_n598_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n420_), .A2(new_n413_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(new_n259_), .A3(new_n320_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n805_), .A2(new_n807_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT121), .ZN(new_n809_));
  AOI21_X1  g608(.A(G113gat), .B1(new_n809_), .B2(new_n679_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n752_), .B1(new_n804_), .B2(new_n622_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n807_), .A2(KEYINPUT59), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT122), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT122), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT57), .B1(new_n787_), .B2(new_n589_), .ZN(new_n816_));
  AOI211_X1 g615(.A(new_n789_), .B(new_n621_), .C1(new_n776_), .C2(new_n786_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n552_), .B1(new_n818_), .B2(new_n802_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n815_), .B(new_n812_), .C1(new_n819_), .C2(new_n752_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n814_), .A2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT59), .B1(new_n805_), .B2(new_n807_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n679_), .A2(G113gat), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n810_), .B1(new_n823_), .B2(new_n824_), .ZN(G1340gat));
  NAND4_X1  g624(.A1(new_n821_), .A2(KEYINPUT123), .A3(new_n491_), .A4(new_n822_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n822_), .A2(new_n814_), .A3(new_n491_), .A4(new_n820_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT123), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n826_), .A2(G120gat), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT60), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n490_), .B2(G120gat), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n809_), .B(new_n832_), .C1(new_n831_), .C2(G120gat), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n830_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(KEYINPUT124), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT124), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n830_), .A2(new_n836_), .A3(new_n833_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(G1341gat));
  AOI21_X1  g637(.A(G127gat), .B1(new_n809_), .B2(new_n552_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n599_), .A2(G127gat), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n839_), .B1(new_n823_), .B2(new_n840_), .ZN(G1342gat));
  AOI21_X1  g640(.A(G134gat), .B1(new_n809_), .B2(new_n621_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n630_), .A2(G134gat), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n842_), .B1(new_n823_), .B2(new_n843_), .ZN(G1343gat));
  NOR2_X1   g643(.A1(new_n805_), .A2(new_n405_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n806_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n846_), .A2(new_n531_), .ZN(new_n847_));
  XOR2_X1   g646(.A(new_n847_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g647(.A1(new_n846_), .A2(new_n490_), .ZN(new_n849_));
  XOR2_X1   g648(.A(new_n849_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g649(.A1(new_n846_), .A2(new_n622_), .ZN(new_n851_));
  XOR2_X1   g650(.A(KEYINPUT61), .B(G155gat), .Z(new_n852_));
  XNOR2_X1  g651(.A(new_n851_), .B(new_n852_), .ZN(G1346gat));
  INV_X1    g652(.A(G162gat), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n846_), .B2(new_n589_), .ZN(new_n855_));
  XOR2_X1   g654(.A(new_n855_), .B(KEYINPUT125), .Z(new_n856_));
  NOR3_X1   g655(.A1(new_n846_), .A2(new_n854_), .A3(new_n593_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(G1347gat));
  INV_X1    g657(.A(KEYINPUT62), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n421_), .A2(new_n394_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n259_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n811_), .A2(new_n404_), .A3(new_n861_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n862_), .A2(new_n679_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n859_), .B1(new_n863_), .B2(new_n205_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n863_), .A2(new_n205_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n865_), .B1(new_n354_), .B2(new_n863_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n864_), .B1(new_n866_), .B2(new_n859_), .ZN(G1348gat));
  AOI21_X1  g666(.A(G176gat), .B1(new_n862_), .B2(new_n491_), .ZN(new_n868_));
  OR2_X1    g667(.A1(new_n805_), .A2(new_n404_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n869_), .A2(new_n206_), .A3(new_n490_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n861_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n868_), .B1(new_n870_), .B2(new_n871_), .ZN(G1349gat));
  OR3_X1    g671(.A1(new_n869_), .A2(new_n622_), .A3(new_n861_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n598_), .A2(new_n217_), .ZN(new_n874_));
  AOI22_X1  g673(.A1(new_n873_), .A2(new_n210_), .B1(new_n862_), .B2(new_n874_), .ZN(G1350gat));
  NAND3_X1  g674(.A1(new_n862_), .A2(new_n220_), .A3(new_n621_), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n862_), .A2(new_n630_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n877_), .B2(new_n211_), .ZN(G1351gat));
  NAND2_X1  g677(.A1(new_n845_), .A2(new_n860_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(new_n531_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(new_n267_), .ZN(G1352gat));
  INV_X1    g680(.A(new_n879_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n491_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(G204gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(new_n883_), .B2(new_n269_), .ZN(G1353gat));
  NOR2_X1   g684(.A1(new_n879_), .A2(new_n598_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n886_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n887_), .A2(KEYINPUT126), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(KEYINPUT126), .ZN(new_n889_));
  XOR2_X1   g688(.A(KEYINPUT63), .B(G211gat), .Z(new_n890_));
  AOI22_X1  g689(.A1(new_n888_), .A2(new_n889_), .B1(new_n886_), .B2(new_n890_), .ZN(G1354gat));
  AOI21_X1  g690(.A(G218gat), .B1(new_n882_), .B2(new_n621_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n630_), .A2(G218gat), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(KEYINPUT127), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n892_), .B1(new_n882_), .B2(new_n894_), .ZN(G1355gat));
endmodule


