//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n887_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n913_, new_n914_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_, new_n938_;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(new_n202_), .A2(KEYINPUT94), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT93), .ZN(new_n204_));
  INV_X1    g003(.A(G204gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n204_), .B1(new_n205_), .B2(G197gat), .ZN(new_n206_));
  INV_X1    g005(.A(G197gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(KEYINPUT93), .A3(G204gat), .ZN(new_n208_));
  OAI211_X1 g007(.A(new_n206_), .B(new_n208_), .C1(new_n207_), .C2(G204gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n202_), .A2(KEYINPUT94), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n203_), .A2(KEYINPUT21), .A3(new_n209_), .A4(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n205_), .A2(G197gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n207_), .A2(G204gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT21), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n214_), .B(new_n202_), .C1(new_n209_), .C2(KEYINPUT21), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n211_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G228gat), .ZN(new_n217_));
  INV_X1    g016(.A(G233gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT91), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT90), .ZN(new_n225_));
  AOI21_X1  g024(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT89), .ZN(new_n227_));
  AND3_X1   g026(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n230_));
  NOR3_X1   g029(.A1(new_n230_), .A2(G141gat), .A3(G148gat), .ZN(new_n231_));
  INV_X1    g030(.A(G141gat), .ZN(new_n232_));
  INV_X1    g031(.A(G148gat), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT3), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n229_), .B1(new_n231_), .B2(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n225_), .B1(new_n227_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G141gat), .A2(G148gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT2), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT89), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT89), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n226_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(G141gat), .A2(G148gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT3), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n230_), .B1(G141gat), .B2(G148gat), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n228_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n243_), .A2(new_n247_), .A3(KEYINPUT90), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n224_), .B1(new_n236_), .B2(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n222_), .B1(KEYINPUT1), .B2(new_n220_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n250_), .B1(KEYINPUT1), .B2(new_n220_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n244_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n251_), .A2(new_n237_), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n219_), .B1(new_n249_), .B2(new_n254_), .ZN(new_n255_));
  AND3_X1   g054(.A1(new_n243_), .A2(KEYINPUT90), .A3(new_n247_), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT90), .B1(new_n243_), .B2(new_n247_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n223_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(KEYINPUT91), .A3(new_n253_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n255_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT29), .ZN(new_n261_));
  OAI221_X1 g060(.A(new_n216_), .B1(new_n217_), .B2(new_n218_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT29), .B1(new_n249_), .B2(new_n254_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(new_n216_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n217_), .A2(new_n218_), .ZN(new_n265_));
  AOI21_X1  g064(.A(KEYINPUT95), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n264_), .A2(KEYINPUT95), .A3(new_n265_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n262_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT97), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G78gat), .B(G106gat), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n268_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n270_), .ZN(new_n272_));
  OAI221_X1 g071(.A(new_n262_), .B1(KEYINPUT97), .B2(new_n272_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n260_), .A2(new_n261_), .ZN(new_n274_));
  XOR2_X1   g073(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(G22gat), .B(G50gat), .Z(new_n277_));
  INV_X1    g076(.A(new_n275_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n260_), .A2(new_n261_), .A3(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n276_), .A2(new_n277_), .A3(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n276_), .A2(new_n279_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n277_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n271_), .A2(new_n273_), .A3(new_n280_), .A4(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n280_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n268_), .A2(KEYINPUT96), .A3(new_n272_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n270_), .B(KEYINPUT96), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n262_), .B(new_n287_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n285_), .A2(new_n286_), .A3(new_n288_), .ZN(new_n289_));
  AND2_X1   g088(.A1(new_n284_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT85), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT85), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(G183gat), .A3(G190gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT23), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT23), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n291_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  NOR3_X1   g098(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT24), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n301_), .B1(G169gat), .B2(G176gat), .ZN(new_n302_));
  INV_X1    g101(.A(G169gat), .ZN(new_n303_));
  INV_X1    g102(.A(G176gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n300_), .B1(new_n302_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT26), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(G190gat), .ZN(new_n308_));
  INV_X1    g107(.A(G190gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT26), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT25), .ZN(new_n311_));
  INV_X1    g110(.A(G183gat), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n308_), .B(new_n310_), .C1(new_n313_), .C2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n306_), .A2(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT98), .B1(new_n299_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n298_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n318_), .B1(new_n295_), .B2(KEYINPUT23), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT98), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n319_), .A2(new_n320_), .A3(new_n306_), .A4(new_n315_), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n317_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT22), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(G169gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n303_), .A2(KEYINPUT22), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT99), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT22), .B(G169gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT99), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n327_), .A2(new_n330_), .A3(new_n304_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G169gat), .A2(G176gat), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n295_), .A2(new_n297_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n291_), .A2(KEYINPUT23), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n312_), .A2(new_n309_), .ZN(new_n337_));
  AOI21_X1  g136(.A(KEYINPUT100), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(KEYINPUT23), .B1(new_n292_), .B2(new_n294_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n335_), .ZN(new_n340_));
  OAI211_X1 g139(.A(KEYINPUT100), .B(new_n337_), .C1(new_n339_), .C2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n333_), .B1(new_n338_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n216_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n322_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G226gat), .A2(G233gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT19), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT20), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT83), .B(G183gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n309_), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n296_), .A2(new_n298_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT86), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n328_), .A2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(G176gat), .B1(new_n324_), .B2(new_n353_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n332_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT26), .B1(new_n309_), .B2(KEYINPUT84), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n358_), .B1(KEYINPUT84), .B2(new_n308_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n312_), .A2(KEYINPUT83), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n312_), .A2(KEYINPUT83), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT25), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n314_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n359_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n306_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n365_));
  OAI22_X1  g164(.A1(new_n352_), .A2(new_n357_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n349_), .B1(new_n366_), .B2(new_n216_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n345_), .A2(new_n348_), .A3(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G8gat), .B(G36gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT18), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G64gat), .B(G92gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT20), .B1(new_n366_), .B2(new_n216_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n322_), .A2(new_n343_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n374_), .B1(new_n375_), .B2(new_n216_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n368_), .B(new_n373_), .C1(new_n376_), .C2(new_n348_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n348_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n367_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n331_), .A2(new_n332_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT100), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n339_), .A2(new_n340_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n337_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n381_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n380_), .B1(new_n384_), .B2(new_n341_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n299_), .A2(new_n316_), .ZN(new_n386_));
  NOR3_X1   g185(.A1(new_n385_), .A2(new_n216_), .A3(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n347_), .B1(new_n379_), .B2(new_n387_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n378_), .A2(new_n388_), .ZN(new_n389_));
  OAI211_X1 g188(.A(KEYINPUT27), .B(new_n377_), .C1(new_n389_), .C2(new_n373_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n317_), .A2(new_n321_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n385_), .A2(new_n391_), .A3(new_n216_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n364_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n365_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n319_), .A2(new_n351_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n326_), .A2(KEYINPUT86), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n396_), .A2(new_n355_), .B1(G169gat), .B2(G176gat), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n393_), .A2(new_n394_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  OAI211_X1 g197(.A(KEYINPUT20), .B(new_n348_), .C1(new_n398_), .C2(new_n344_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n392_), .A2(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n216_), .B1(new_n385_), .B2(new_n391_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n349_), .B1(new_n398_), .B2(new_n344_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n348_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n372_), .B1(new_n400_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(new_n377_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT27), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n390_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n290_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G227gat), .A2(G233gat), .ZN(new_n411_));
  INV_X1    g210(.A(G15gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(G71gat), .ZN(new_n414_));
  INV_X1    g213(.A(G99gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT87), .B(G43gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n366_), .B(KEYINPUT30), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT88), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n418_), .A2(new_n420_), .ZN(new_n421_));
  XOR2_X1   g220(.A(new_n419_), .B(KEYINPUT88), .Z(new_n422_));
  OAI21_X1  g221(.A(new_n421_), .B1(new_n422_), .B2(new_n418_), .ZN(new_n423_));
  XOR2_X1   g222(.A(G127gat), .B(G134gat), .Z(new_n424_));
  XNOR2_X1  g223(.A(G113gat), .B(G120gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT31), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  OR2_X1    g227(.A1(new_n423_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n423_), .A2(new_n428_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  XOR2_X1   g230(.A(G1gat), .B(G29gat), .Z(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G57gat), .B(G85gat), .ZN(new_n435_));
  XOR2_X1   g234(.A(new_n434_), .B(new_n435_), .Z(new_n436_));
  NAND2_X1  g235(.A1(G225gat), .A2(G233gat), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n255_), .A2(new_n259_), .A3(new_n426_), .ZN(new_n438_));
  OR3_X1    g237(.A1(new_n249_), .A2(new_n254_), .A3(new_n426_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT4), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT4), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n438_), .A2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n437_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n438_), .A2(new_n437_), .A3(new_n439_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT102), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT102), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n438_), .A2(new_n447_), .A3(new_n437_), .A4(new_n439_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n436_), .B1(new_n444_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n437_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n438_), .A2(new_n442_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n442_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n451_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n436_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n454_), .A2(new_n455_), .A3(new_n446_), .A4(new_n448_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n450_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n431_), .A2(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n410_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT33), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n456_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n449_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n462_), .A2(KEYINPUT33), .A3(new_n455_), .A4(new_n454_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n437_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n440_), .A2(new_n437_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n465_), .A2(new_n455_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n405_), .B1(new_n464_), .B2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n461_), .A2(new_n463_), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT103), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n373_), .A2(KEYINPUT32), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n368_), .B(new_n470_), .C1(new_n376_), .C2(new_n348_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n471_), .B1(new_n389_), .B2(new_n470_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n472_), .B1(new_n450_), .B2(new_n456_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n468_), .B1(new_n469_), .B2(new_n473_), .ZN(new_n474_));
  AOI211_X1 g273(.A(KEYINPUT103), .B(new_n472_), .C1(new_n456_), .C2(new_n450_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n290_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n284_), .A2(new_n289_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n477_), .A2(new_n457_), .A3(new_n409_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n431_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n459_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G29gat), .B(G36gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G43gat), .B(G50gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT15), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G15gat), .B(G22gat), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT76), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(G1gat), .ZN(new_n492_));
  INV_X1    g291(.A(G8gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT14), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT77), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n491_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G1gat), .B(G8gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n488_), .A2(new_n498_), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n498_), .A2(new_n486_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G229gat), .A2(G233gat), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n498_), .B(new_n486_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n501_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  XOR2_X1   g305(.A(G113gat), .B(G141gat), .Z(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT80), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G169gat), .B(G197gat), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n508_), .B(new_n509_), .Z(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT82), .B1(new_n506_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT82), .ZN(new_n512_));
  INV_X1    g311(.A(new_n510_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n502_), .A2(new_n505_), .A3(new_n512_), .A4(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n511_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT79), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n506_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT81), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n502_), .A2(new_n505_), .A3(KEYINPUT79), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .A4(new_n510_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n515_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n517_), .A2(new_n519_), .A3(new_n510_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT81), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n481_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G231gat), .A2(G233gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n498_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G57gat), .B(G64gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT11), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G71gat), .B(G78gat), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n530_), .A2(new_n532_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n529_), .A2(KEYINPUT11), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n534_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n528_), .B(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT78), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G127gat), .B(G155gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT16), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G183gat), .B(G211gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT17), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n540_), .B(new_n545_), .ZN(new_n546_));
  OR3_X1    g345(.A1(new_n539_), .A2(KEYINPUT17), .A3(new_n544_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(G190gat), .B(G218gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT73), .ZN(new_n550_));
  XOR2_X1   g349(.A(G134gat), .B(G162gat), .Z(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT36), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(KEYINPUT10), .B(G99gat), .Z(new_n555_));
  XOR2_X1   g354(.A(KEYINPUT64), .B(G106gat), .Z(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT65), .ZN(new_n558_));
  INV_X1    g357(.A(G85gat), .ZN(new_n559_));
  INV_X1    g358(.A(G92gat), .ZN(new_n560_));
  NOR3_X1   g359(.A1(new_n559_), .A2(new_n560_), .A3(KEYINPUT9), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G99gat), .A2(G106gat), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT6), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G85gat), .B(G92gat), .Z(new_n565_));
  AOI211_X1 g364(.A(new_n561_), .B(new_n564_), .C1(KEYINPUT9), .C2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n558_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT66), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n558_), .A2(KEYINPUT66), .A3(new_n566_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(G106gat), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n415_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT7), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n565_), .B1(new_n574_), .B2(new_n564_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT67), .ZN(new_n576_));
  AOI21_X1  g375(.A(KEYINPUT8), .B1(new_n565_), .B2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n575_), .B(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n571_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n488_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n578_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n486_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G232gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT34), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT35), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n581_), .A2(new_n584_), .A3(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(KEYINPUT72), .B1(new_n590_), .B2(KEYINPUT74), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n587_), .A2(new_n588_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n591_), .B(new_n592_), .C1(KEYINPUT72), .C2(new_n590_), .ZN(new_n593_));
  OAI221_X1 g392(.A(KEYINPUT72), .B1(new_n588_), .B2(new_n587_), .C1(new_n590_), .C2(KEYINPUT74), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n554_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n593_), .A2(new_n594_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n552_), .B(KEYINPUT36), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n596_), .B(KEYINPUT37), .C1(new_n597_), .C2(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n599_), .B1(new_n597_), .B2(KEYINPUT75), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT75), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n593_), .A2(new_n602_), .A3(new_n594_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n595_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n604_));
  OAI211_X1 g403(.A(new_n548_), .B(new_n600_), .C1(new_n604_), .C2(KEYINPUT37), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n571_), .A2(new_n537_), .A3(new_n579_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT68), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n580_), .A2(new_n538_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT68), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n582_), .A2(new_n609_), .A3(new_n537_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n607_), .A2(new_n608_), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G230gat), .A2(G233gat), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT69), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT69), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n611_), .A2(new_n616_), .A3(new_n613_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n608_), .A2(KEYINPUT12), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n582_), .A2(new_n537_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT12), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n618_), .A2(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n613_), .B1(new_n582_), .B2(new_n537_), .ZN(new_n623_));
  AOI22_X1  g422(.A1(new_n615_), .A2(new_n617_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G120gat), .B(G148gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT5), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G176gat), .B(G204gat), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n626_), .B(new_n627_), .Z(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n624_), .B(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT13), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n624_), .A2(new_n629_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n608_), .A2(KEYINPUT12), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n619_), .A2(new_n620_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n623_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n617_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n616_), .B1(new_n611_), .B2(new_n613_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n636_), .B(new_n629_), .C1(new_n637_), .C2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n633_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT13), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n632_), .A2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n605_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n526_), .A2(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT104), .Z(new_n646_));
  INV_X1    g445(.A(new_n457_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n646_), .A2(new_n492_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT38), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n481_), .A2(new_n604_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n548_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n643_), .A2(new_n525_), .A3(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(G1gat), .B1(new_n654_), .B2(new_n457_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n648_), .A2(new_n649_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n650_), .A2(new_n655_), .A3(new_n656_), .ZN(G1324gat));
  OAI21_X1  g456(.A(G8gat), .B1(new_n654_), .B2(new_n409_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT105), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n659_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n660_), .A2(KEYINPUT39), .A3(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n646_), .A2(new_n493_), .A3(new_n408_), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n661_), .A2(KEYINPUT39), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n662_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT40), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n662_), .A2(new_n663_), .A3(KEYINPUT40), .A4(new_n664_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1325gat));
  NAND4_X1  g468(.A1(new_n526_), .A2(new_n644_), .A3(new_n412_), .A4(new_n431_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n671_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G15gat), .B1(new_n654_), .B2(new_n480_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT41), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n675_), .A2(KEYINPUT41), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n674_), .A2(new_n676_), .A3(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT107), .ZN(G1326gat));
  OAI21_X1  g478(.A(G22gat), .B1(new_n654_), .B2(new_n290_), .ZN(new_n680_));
  XOR2_X1   g479(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n290_), .A2(G22gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n682_), .B1(new_n645_), .B2(new_n683_), .ZN(G1327gat));
  NOR2_X1   g483(.A1(new_n597_), .A2(new_n599_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT37), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n685_), .A2(new_n686_), .A3(new_n595_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n597_), .A2(KEYINPUT75), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n688_), .A2(new_n603_), .A3(new_n598_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n596_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n687_), .B1(new_n690_), .B2(new_n686_), .ZN(new_n691_));
  OAI21_X1  g490(.A(KEYINPUT43), .B1(new_n481_), .B2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n600_), .B1(new_n604_), .B2(KEYINPUT37), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n431_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n693_), .B(new_n694_), .C1(new_n695_), .C2(new_n459_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n692_), .A2(new_n696_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n643_), .A2(new_n525_), .A3(new_n548_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n697_), .A2(KEYINPUT44), .A3(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(KEYINPUT44), .B1(new_n697_), .B2(new_n698_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n699_), .A2(new_n700_), .A3(new_n457_), .ZN(new_n701_));
  INV_X1    g500(.A(G29gat), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n604_), .A2(new_n652_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n643_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n526_), .A2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n647_), .A2(new_n702_), .ZN(new_n706_));
  OAI22_X1  g505(.A1(new_n701_), .A2(new_n702_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT109), .ZN(G1328gat));
  INV_X1    g507(.A(new_n705_), .ZN(new_n709_));
  INV_X1    g508(.A(G36gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n709_), .A2(new_n710_), .A3(new_n408_), .ZN(new_n711_));
  XOR2_X1   g510(.A(KEYINPUT111), .B(KEYINPUT45), .Z(new_n712_));
  XNOR2_X1  g511(.A(KEYINPUT110), .B(KEYINPUT112), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n712_), .B(new_n713_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n711_), .B(new_n714_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n699_), .A2(new_n700_), .A3(new_n409_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n715_), .B1(new_n710_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT46), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n715_), .B(KEYINPUT46), .C1(new_n710_), .C2(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1329gat));
  AOI21_X1  g520(.A(G43gat), .B1(new_n709_), .B2(new_n431_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n699_), .A2(new_n700_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n431_), .A2(G43gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n722_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n725_), .B(new_n726_), .ZN(G1330gat));
  AOI21_X1  g526(.A(G50gat), .B1(new_n709_), .B2(new_n477_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n477_), .A2(G50gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n723_), .B2(new_n729_), .ZN(G1331gat));
  NAND2_X1  g529(.A1(new_n643_), .A2(new_n525_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n731_), .A2(new_n652_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n732_), .A2(new_n651_), .A3(G57gat), .A4(new_n647_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT115), .Z(new_n734_));
  NOR2_X1   g533(.A1(new_n481_), .A2(new_n524_), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n735_), .A2(new_n643_), .A3(new_n548_), .A4(new_n691_), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n736_), .A2(KEYINPUT114), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n457_), .B1(new_n736_), .B2(KEYINPUT114), .ZN(new_n738_));
  AOI21_X1  g537(.A(G57gat), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n734_), .A2(new_n739_), .ZN(G1332gat));
  NAND2_X1  g539(.A1(new_n732_), .A2(new_n651_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G64gat), .B1(new_n741_), .B2(new_n409_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT48), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n409_), .A2(G64gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n736_), .B2(new_n744_), .ZN(G1333gat));
  OAI21_X1  g544(.A(G71gat), .B1(new_n741_), .B2(new_n480_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT49), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n480_), .A2(G71gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n736_), .B2(new_n748_), .ZN(G1334gat));
  OAI21_X1  g548(.A(G78gat), .B1(new_n741_), .B2(new_n290_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n750_), .B(new_n751_), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n290_), .A2(G78gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n752_), .B1(new_n736_), .B2(new_n753_), .ZN(G1335gat));
  INV_X1    g553(.A(new_n643_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n755_), .A2(new_n703_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n735_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(new_n559_), .A3(new_n647_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n643_), .A2(new_n525_), .A3(new_n652_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n692_), .B2(new_n696_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n761_), .A2(new_n647_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n759_), .B1(new_n762_), .B2(new_n559_), .ZN(G1336gat));
  NAND3_X1  g562(.A1(new_n758_), .A2(new_n560_), .A3(new_n408_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n761_), .A2(new_n408_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(new_n560_), .ZN(G1337gat));
  AOI21_X1  g565(.A(new_n415_), .B1(new_n761_), .B2(new_n431_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n431_), .A2(new_n555_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n758_), .B2(new_n768_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT51), .Z(G1338gat));
  XNOR2_X1  g569(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT118), .ZN(new_n773_));
  AOI211_X1 g572(.A(new_n290_), .B(new_n760_), .C1(new_n692_), .C2(new_n696_), .ZN(new_n774_));
  OAI21_X1  g573(.A(KEYINPUT52), .B1(new_n774_), .B2(new_n572_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n760_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n697_), .A2(new_n477_), .A3(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n777_), .A2(new_n778_), .A3(G106gat), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n775_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n556_), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n757_), .A2(new_n290_), .A3(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n773_), .B1(new_n780_), .B2(new_n783_), .ZN(new_n784_));
  AOI211_X1 g583(.A(KEYINPUT118), .B(new_n782_), .C1(new_n775_), .C2(new_n779_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n772_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n774_), .A2(KEYINPUT52), .A3(new_n572_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n778_), .B1(new_n777_), .B2(G106gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n783_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT118), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n780_), .A2(new_n773_), .A3(new_n783_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n791_), .A3(new_n771_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n786_), .A2(new_n792_), .ZN(G1339gat));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n636_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n622_), .A2(KEYINPUT55), .A3(new_n623_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n607_), .A2(new_n610_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n612_), .B1(new_n622_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT119), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n795_), .B(new_n796_), .C1(new_n798_), .C2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n799_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n628_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n640_), .B1(new_n523_), .B2(new_n521_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n628_), .B(new_n804_), .C1(new_n800_), .C2(new_n802_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n806_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n503_), .A2(new_n501_), .ZN(new_n810_));
  OR3_X1    g609(.A1(new_n810_), .A2(KEYINPUT121), .A3(new_n513_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n499_), .A2(new_n500_), .A3(new_n504_), .ZN(new_n812_));
  OAI21_X1  g611(.A(KEYINPUT121), .B1(new_n810_), .B2(new_n513_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n811_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n814_), .A2(new_n515_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n633_), .B2(new_n640_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT122), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n630_), .A2(KEYINPUT122), .A3(new_n815_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n809_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n820_), .A2(KEYINPUT57), .A3(new_n690_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT57), .B1(new_n820_), .B2(new_n690_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT58), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT56), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n825_), .B(new_n628_), .C1(new_n800_), .C2(new_n802_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n826_), .A2(new_n639_), .A3(new_n815_), .ZN(new_n827_));
  OR2_X1    g626(.A1(new_n798_), .A2(new_n799_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n828_), .A2(new_n801_), .A3(new_n795_), .A4(new_n796_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n825_), .B1(new_n829_), .B2(new_n628_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n824_), .B1(new_n827_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n693_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT123), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  OR3_X1    g633(.A1(new_n827_), .A2(new_n830_), .A3(new_n824_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n831_), .A2(new_n693_), .A3(KEYINPUT123), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n834_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n548_), .B1(new_n823_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n839_), .B1(new_n644_), .B2(new_n525_), .ZN(new_n840_));
  NOR4_X1   g639(.A1(new_n605_), .A2(new_n643_), .A3(KEYINPUT54), .A4(new_n524_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n838_), .A2(new_n842_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n410_), .A2(new_n480_), .A3(new_n457_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n843_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(G113gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(new_n847_), .A3(new_n524_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT59), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n843_), .B2(new_n845_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n820_), .A2(new_n690_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n820_), .A2(KEYINPUT57), .A3(new_n690_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n836_), .A2(new_n835_), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT123), .B1(new_n831_), .B2(new_n693_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n853_), .B(new_n854_), .C1(new_n855_), .C2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n652_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n842_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n860_), .A2(KEYINPUT59), .A3(new_n844_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n525_), .B1(new_n850_), .B2(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n848_), .B1(new_n862_), .B2(new_n847_), .ZN(G1340gat));
  INV_X1    g662(.A(KEYINPUT60), .ZN(new_n864_));
  AOI21_X1  g663(.A(G120gat), .B1(new_n643_), .B2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT124), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT124), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n867_), .B1(new_n864_), .B2(G120gat), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n846_), .B(new_n866_), .C1(new_n865_), .C2(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n755_), .B1(new_n850_), .B2(new_n861_), .ZN(new_n870_));
  INV_X1    g669(.A(G120gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n869_), .B1(new_n870_), .B2(new_n871_), .ZN(G1341gat));
  INV_X1    g671(.A(G127gat), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n846_), .A2(new_n873_), .A3(new_n548_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n652_), .B1(new_n850_), .B2(new_n861_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(new_n873_), .ZN(G1342gat));
  INV_X1    g675(.A(G134gat), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n846_), .A2(new_n877_), .A3(new_n604_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n691_), .B1(new_n850_), .B2(new_n861_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n879_), .B2(new_n877_), .ZN(G1343gat));
  NOR2_X1   g679(.A1(new_n290_), .A2(new_n408_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n882_), .A2(new_n457_), .A3(new_n431_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n843_), .A2(new_n525_), .A3(new_n884_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(new_n232_), .ZN(G1344gat));
  NOR3_X1   g685(.A1(new_n843_), .A2(new_n755_), .A3(new_n884_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(new_n233_), .ZN(G1345gat));
  OAI211_X1 g687(.A(new_n548_), .B(new_n883_), .C1(new_n838_), .C2(new_n842_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(KEYINPUT125), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT125), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n860_), .A2(new_n891_), .A3(new_n548_), .A4(new_n883_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(KEYINPUT61), .B(G155gat), .ZN(new_n893_));
  AND3_X1   g692(.A1(new_n890_), .A2(new_n892_), .A3(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n893_), .B1(new_n890_), .B2(new_n892_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1346gat));
  INV_X1    g695(.A(G162gat), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n860_), .A2(new_n897_), .A3(new_n604_), .A4(new_n883_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n843_), .A2(new_n691_), .A3(new_n884_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n897_), .ZN(G1347gat));
  NOR3_X1   g699(.A1(new_n458_), .A2(new_n477_), .A3(new_n409_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n860_), .A2(new_n524_), .A3(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(G169gat), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n901_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n843_), .A2(new_n906_), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n907_), .A2(new_n327_), .A3(new_n330_), .A4(new_n524_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n902_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n905_), .A2(new_n908_), .A3(new_n909_), .ZN(G1348gat));
  NOR3_X1   g709(.A1(new_n843_), .A2(new_n755_), .A3(new_n906_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(new_n304_), .ZN(G1349gat));
  INV_X1    g711(.A(new_n350_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n913_), .B1(new_n907_), .B2(new_n548_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n313_), .A2(new_n314_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n843_), .A2(new_n652_), .A3(new_n906_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n914_), .B1(new_n915_), .B2(new_n916_), .ZN(G1350gat));
  NAND4_X1  g716(.A1(new_n907_), .A2(new_n308_), .A3(new_n310_), .A4(new_n604_), .ZN(new_n918_));
  NOR3_X1   g717(.A1(new_n843_), .A2(new_n691_), .A3(new_n906_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n309_), .B2(new_n919_), .ZN(G1351gat));
  NOR4_X1   g719(.A1(new_n290_), .A2(new_n431_), .A3(new_n647_), .A4(new_n409_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n860_), .A2(new_n524_), .A3(new_n921_), .ZN(new_n922_));
  OAI21_X1  g721(.A(KEYINPUT126), .B1(new_n922_), .B2(new_n207_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n207_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n921_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n925_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n927_));
  NAND4_X1  g726(.A1(new_n926_), .A2(new_n927_), .A3(G197gat), .A4(new_n524_), .ZN(new_n928_));
  AND3_X1   g727(.A1(new_n923_), .A2(new_n924_), .A3(new_n928_), .ZN(G1352gat));
  NAND2_X1  g728(.A1(new_n926_), .A2(new_n643_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g730(.A(KEYINPUT63), .B(G211gat), .C1(new_n926_), .C2(new_n548_), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n843_), .A2(new_n652_), .A3(new_n925_), .ZN(new_n933_));
  XOR2_X1   g732(.A(KEYINPUT63), .B(G211gat), .Z(new_n934_));
  AOI21_X1  g733(.A(new_n932_), .B1(new_n933_), .B2(new_n934_), .ZN(G1354gat));
  AOI21_X1  g734(.A(G218gat), .B1(new_n926_), .B2(new_n604_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n693_), .A2(G218gat), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(KEYINPUT127), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n936_), .B1(new_n926_), .B2(new_n938_), .ZN(G1355gat));
endmodule


