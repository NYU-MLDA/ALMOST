//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n623_,
    new_n624_, new_n625_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n855_, new_n856_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n884_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n905_;
  XOR2_X1   g000(.A(KEYINPUT10), .B(G99gat), .Z(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT6), .ZN(new_n206_));
  AND2_X1   g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G92gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G85gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT9), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(KEYINPUT66), .A3(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(G85gat), .ZN(new_n212_));
  INV_X1    g011(.A(G92gat), .ZN(new_n213_));
  NOR3_X1   g012(.A1(new_n210_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n214_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n211_), .A2(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(KEYINPUT66), .B1(new_n209_), .B2(new_n210_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n207_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  XOR2_X1   g017(.A(G85gat), .B(G92gat), .Z(new_n219_));
  OR3_X1    g018(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n206_), .A2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(KEYINPUT67), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n219_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT8), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  OAI211_X1 g025(.A(KEYINPUT8), .B(new_n219_), .C1(new_n221_), .C2(new_n223_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n218_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G29gat), .B(G36gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G43gat), .B(G50gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT73), .B(KEYINPUT15), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT72), .B(KEYINPUT35), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G232gat), .A2(G233gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  AOI22_X1  g036(.A1(new_n228_), .A2(new_n233_), .B1(new_n234_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n231_), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT74), .B1(new_n228_), .B2(new_n239_), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT75), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n237_), .A2(new_n234_), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n226_), .A2(new_n227_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT74), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n244_), .A2(new_n245_), .A3(new_n231_), .A4(new_n218_), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .A4(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n238_), .A2(new_n240_), .A3(new_n246_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n243_), .A2(new_n242_), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT75), .B1(new_n237_), .B2(new_n234_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n247_), .A2(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(G190gat), .B(G218gat), .Z(new_n253_));
  XNOR2_X1  g052(.A(G134gat), .B(G162gat), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n254_), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n257_), .A2(KEYINPUT36), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n258_), .B(KEYINPUT76), .Z(new_n259_));
  NAND2_X1  g058(.A1(new_n252_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT77), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n252_), .A2(KEYINPUT77), .A3(new_n259_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n257_), .A2(KEYINPUT36), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n247_), .A2(new_n251_), .A3(new_n258_), .A4(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n262_), .A2(new_n263_), .A3(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT78), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n266_), .A2(new_n267_), .A3(KEYINPUT37), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n266_), .A2(KEYINPUT37), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n260_), .A2(new_n265_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT78), .B1(new_n270_), .B2(KEYINPUT37), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n268_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G127gat), .B(G155gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT16), .ZN(new_n275_));
  XOR2_X1   g074(.A(G183gat), .B(G211gat), .Z(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT17), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G15gat), .B(G22gat), .ZN(new_n280_));
  INV_X1    g079(.A(G1gat), .ZN(new_n281_));
  INV_X1    g080(.A(G8gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT14), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G1gat), .B(G8gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G231gat), .A2(G233gat), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n286_), .B(new_n287_), .Z(new_n288_));
  XNOR2_X1  g087(.A(G57gat), .B(G64gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT11), .ZN(new_n290_));
  XOR2_X1   g089(.A(G71gat), .B(G78gat), .Z(new_n291_));
  OR2_X1    g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n289_), .A2(KEYINPUT11), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n290_), .A2(new_n291_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n292_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT68), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n279_), .B1(new_n288_), .B2(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n297_), .B1(new_n288_), .B2(new_n296_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n295_), .ZN(new_n299_));
  AOI211_X1 g098(.A(new_n278_), .B(new_n277_), .C1(new_n288_), .C2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n300_), .B1(new_n299_), .B2(new_n288_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n273_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT79), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G226gat), .A2(G233gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT19), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT20), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT21), .ZN(new_n310_));
  INV_X1    g109(.A(G204gat), .ZN(new_n311_));
  INV_X1    g110(.A(G197gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT87), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT87), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(G197gat), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n311_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(G197gat), .A2(G204gat), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n310_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(G218gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(G211gat), .ZN(new_n320_));
  INV_X1    g119(.A(G211gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(G218gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n313_), .A2(new_n315_), .A3(new_n311_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n310_), .B1(G197gat), .B2(G204gat), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n323_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n313_), .A2(new_n315_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n317_), .B1(new_n327_), .B2(G204gat), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n310_), .B1(new_n320_), .B2(new_n322_), .ZN(new_n329_));
  AOI22_X1  g128(.A1(new_n318_), .A2(new_n326_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT24), .ZN(new_n331_));
  INV_X1    g130(.A(G169gat), .ZN(new_n332_));
  INV_X1    g131(.A(G176gat), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n331_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G183gat), .A2(G190gat), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT23), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n334_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G169gat), .A2(G176gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(KEYINPUT24), .ZN(new_n341_));
  NOR2_X1   g140(.A1(G169gat), .A2(G176gat), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n339_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT26), .B(G190gat), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT81), .ZN(new_n346_));
  INV_X1    g145(.A(G183gat), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n346_), .B1(new_n347_), .B2(KEYINPUT25), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT25), .B(G183gat), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n345_), .B(new_n348_), .C1(new_n349_), .C2(new_n346_), .ZN(new_n350_));
  AND3_X1   g149(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  OR2_X1    g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT22), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n356_), .A2(new_n333_), .A3(G169gat), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n332_), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  AOI22_X1  g158(.A1(new_n344_), .A2(new_n350_), .B1(new_n355_), .B2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n309_), .B1(new_n330_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n318_), .A2(new_n326_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n328_), .A2(new_n329_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n341_), .A2(KEYINPUT88), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT88), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n340_), .A2(new_n366_), .A3(KEYINPUT24), .ZN(new_n367_));
  INV_X1    g166(.A(new_n342_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n365_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n339_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n349_), .A2(new_n345_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  AOI22_X1  g171(.A1(new_n353_), .A2(new_n354_), .B1(new_n358_), .B2(new_n357_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n364_), .A2(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n308_), .B1(new_n361_), .B2(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT20), .B1(new_n364_), .B2(new_n375_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n330_), .A2(new_n360_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n377_), .B1(new_n308_), .B2(new_n380_), .ZN(new_n381_));
  XOR2_X1   g180(.A(G8gat), .B(G36gat), .Z(new_n382_));
  XNOR2_X1  g181(.A(G64gat), .B(G92gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n381_), .A2(new_n387_), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n361_), .A2(new_n376_), .A3(new_n308_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n339_), .B1(new_n349_), .B2(new_n345_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n373_), .B1(new_n390_), .B2(new_n369_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n309_), .B1(new_n391_), .B2(new_n330_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n344_), .A2(new_n350_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n374_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n364_), .A2(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n308_), .B1(new_n392_), .B2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT92), .B1(new_n389_), .B2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n361_), .A2(new_n376_), .A3(new_n308_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT92), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n397_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n386_), .B(KEYINPUT96), .ZN(new_n403_));
  OAI211_X1 g202(.A(KEYINPUT27), .B(new_n388_), .C1(new_n402_), .C2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n377_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n392_), .A2(new_n308_), .A3(new_n395_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n386_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n388_), .A2(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(KEYINPUT97), .B(KEYINPUT27), .Z(new_n410_));
  AND3_X1   g209(.A1(new_n409_), .A2(KEYINPUT98), .A3(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(KEYINPUT98), .B1(new_n409_), .B2(new_n410_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n404_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT99), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  OAI211_X1 g214(.A(KEYINPUT99), .B(new_n404_), .C1(new_n411_), .C2(new_n412_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  OR2_X1    g216(.A1(G155gat), .A2(G162gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G155gat), .A2(G162gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT84), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT84), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n423_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(G141gat), .A2(G148gat), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT3), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT2), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n429_), .B1(G141gat), .B2(G148gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G141gat), .A2(G148gat), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n431_), .A2(KEYINPUT2), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n428_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT85), .B1(new_n425_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n431_), .A2(KEYINPUT2), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n429_), .A2(G141gat), .A3(G148gat), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n435_), .A2(new_n436_), .B1(new_n427_), .B2(new_n426_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n422_), .A2(new_n424_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT85), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n420_), .B1(new_n434_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT83), .ZN(new_n442_));
  OR3_X1    g241(.A1(new_n419_), .A2(new_n442_), .A3(KEYINPUT1), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n442_), .B1(new_n419_), .B2(KEYINPUT1), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n419_), .A2(KEYINPUT1), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n443_), .A2(new_n418_), .A3(new_n444_), .A4(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n426_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n446_), .A2(new_n447_), .A3(new_n431_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n441_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT29), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n364_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  XOR2_X1   g251(.A(G22gat), .B(G50gat), .Z(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  XOR2_X1   g254(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n450_), .A2(new_n451_), .A3(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G228gat), .A2(G233gat), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n460_), .B(G78gat), .Z(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(new_n203_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n457_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n463_));
  NOR3_X1   g262(.A1(new_n459_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n462_), .B1(new_n459_), .B2(new_n463_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n455_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n466_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n454_), .B1(new_n468_), .B2(new_n464_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(G127gat), .B(G134gat), .Z(new_n472_));
  XOR2_X1   g271(.A(G113gat), .B(G120gat), .Z(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G127gat), .B(G134gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G113gat), .B(G120gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n474_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT82), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n474_), .A2(KEYINPUT82), .A3(new_n477_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n482_), .B1(new_n441_), .B2(new_n449_), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n439_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n478_), .B(new_n448_), .C1(new_n486_), .C2(new_n420_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G225gat), .A2(G233gat), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n483_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n483_), .A2(KEYINPUT4), .A3(new_n487_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n488_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n491_), .B1(new_n483_), .B2(KEYINPUT4), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n489_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G1gat), .B(G29gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT90), .B(KEYINPUT0), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G57gat), .B(G85gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n493_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT94), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n489_), .B(new_n498_), .C1(new_n490_), .C2(new_n492_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n493_), .A2(KEYINPUT94), .A3(new_n499_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G227gat), .A2(G233gat), .ZN(new_n507_));
  INV_X1    g306(.A(G15gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT30), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n360_), .B(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(new_n482_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G71gat), .B(G99gat), .ZN(new_n513_));
  INV_X1    g312(.A(G43gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT31), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n512_), .B(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n506_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n417_), .A2(new_n471_), .A3(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n470_), .A2(new_n505_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n413_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT95), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n387_), .A2(KEYINPUT32), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n407_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(KEYINPUT93), .B1(new_n401_), .B2(new_n524_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT93), .ZN(new_n528_));
  AOI211_X1 g327(.A(new_n528_), .B(new_n523_), .C1(new_n397_), .C2(new_n400_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n526_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n522_), .B1(new_n530_), .B2(new_n505_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n307_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n399_), .B1(new_n532_), .B2(new_n398_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n400_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n524_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n528_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n401_), .A2(KEYINPUT93), .A3(new_n524_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n525_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n538_), .A2(KEYINPUT95), .A3(new_n504_), .A4(new_n503_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n502_), .A2(KEYINPUT91), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n540_), .A2(KEYINPUT33), .ZN(new_n541_));
  INV_X1    g340(.A(new_n409_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(KEYINPUT33), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n483_), .A2(new_n487_), .A3(new_n491_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n488_), .B1(new_n483_), .B2(KEYINPUT4), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n499_), .B(new_n544_), .C1(new_n490_), .C2(new_n545_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .A4(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n531_), .A2(new_n539_), .A3(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n521_), .B1(new_n548_), .B2(new_n471_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n517_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n519_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT70), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT68), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n295_), .B(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(new_n228_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n296_), .A2(new_n244_), .A3(new_n218_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n228_), .A2(KEYINPUT12), .A3(new_n299_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n557_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G230gat), .A2(G233gat), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n561_), .B(KEYINPUT64), .Z(new_n562_));
  OAI21_X1  g361(.A(new_n552_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n558_), .A2(new_n555_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(new_n562_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n558_), .A2(new_n559_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n562_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n566_), .A2(KEYINPUT70), .A3(new_n567_), .A4(new_n557_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n563_), .A2(new_n565_), .A3(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G120gat), .B(G148gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT5), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G176gat), .B(G204gat), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n571_), .B(new_n572_), .Z(new_n573_));
  NAND2_X1  g372(.A1(new_n569_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n573_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n563_), .A2(new_n565_), .A3(new_n568_), .A4(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT13), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n574_), .A2(KEYINPUT13), .A3(new_n576_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n286_), .A2(new_n239_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G229gat), .A2(G233gat), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n233_), .A2(new_n286_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n286_), .B(new_n239_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n583_), .ZN(new_n587_));
  AOI22_X1  g386(.A1(new_n584_), .A2(new_n585_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G113gat), .B(G141gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G169gat), .B(G197gat), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n589_), .B(new_n590_), .Z(new_n591_));
  NAND2_X1  g390(.A1(new_n588_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT80), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n588_), .A2(new_n591_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n581_), .A2(new_n597_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n551_), .A2(new_n598_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n305_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n600_), .A2(new_n281_), .A3(new_n506_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT38), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n598_), .A2(KEYINPUT100), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT100), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n605_), .B1(new_n581_), .B2(new_n597_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n302_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n551_), .A2(new_n270_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(G1gat), .B1(new_n609_), .B2(new_n505_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n601_), .A2(new_n602_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n603_), .A2(new_n610_), .A3(new_n611_), .ZN(G1324gat));
  INV_X1    g411(.A(new_n417_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n600_), .A2(new_n282_), .A3(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT101), .ZN(new_n615_));
  OAI21_X1  g414(.A(G8gat), .B1(new_n609_), .B2(new_n417_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT39), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT40), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n615_), .A2(KEYINPUT40), .A3(new_n617_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(G1325gat));
  OAI21_X1  g421(.A(G15gat), .B1(new_n609_), .B2(new_n517_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT41), .Z(new_n624_));
  NAND3_X1  g423(.A1(new_n600_), .A2(new_n508_), .A3(new_n550_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(G1326gat));
  OAI21_X1  g425(.A(G22gat), .B1(new_n609_), .B2(new_n471_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT42), .ZN(new_n628_));
  INV_X1    g427(.A(G22gat), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n600_), .A2(new_n629_), .A3(new_n470_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT102), .Z(G1327gat));
  AOI21_X1  g431(.A(new_n303_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT43), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n551_), .A2(new_n634_), .A3(new_n272_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n634_), .B1(new_n551_), .B2(new_n272_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n633_), .B(KEYINPUT44), .C1(new_n635_), .C2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT103), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n551_), .A2(new_n272_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(KEYINPUT43), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n551_), .A2(new_n634_), .A3(new_n272_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n643_), .A2(KEYINPUT103), .A3(KEYINPUT44), .A4(new_n633_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n639_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n633_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT44), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n645_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(G29gat), .B1(new_n650_), .B2(new_n505_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n270_), .A2(new_n303_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n599_), .A2(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n505_), .A2(G29gat), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT104), .Z(new_n655_));
  OAI21_X1  g454(.A(new_n651_), .B1(new_n653_), .B2(new_n655_), .ZN(G1328gat));
  INV_X1    g455(.A(KEYINPUT108), .ZN(new_n657_));
  INV_X1    g456(.A(G36gat), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n599_), .A2(new_n658_), .A3(new_n613_), .A4(new_n652_), .ZN(new_n659_));
  XOR2_X1   g458(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n580_), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT13), .B1(new_n574_), .B2(new_n576_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT100), .B1(new_n664_), .B2(new_n596_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n581_), .A2(new_n605_), .A3(new_n597_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n302_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n667_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n613_), .B1(new_n668_), .B2(KEYINPUT44), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n669_), .B1(new_n639_), .B2(new_n644_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n661_), .B1(new_n670_), .B2(new_n658_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT46), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n657_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n417_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n658_), .B1(new_n645_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n661_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n677_), .A2(KEYINPUT108), .A3(KEYINPUT46), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n673_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT106), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT46), .B1(new_n671_), .B2(new_n681_), .ZN(new_n682_));
  OAI211_X1 g481(.A(KEYINPUT106), .B(new_n661_), .C1(new_n670_), .C2(new_n658_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n680_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n681_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n685_));
  AND4_X1   g484(.A1(new_n680_), .A2(new_n685_), .A3(new_n683_), .A4(new_n672_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n679_), .B1(new_n684_), .B2(new_n686_), .ZN(G1329gat));
  INV_X1    g486(.A(KEYINPUT109), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n550_), .A2(G43gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n650_), .B2(new_n689_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n649_), .A2(KEYINPUT109), .A3(G43gat), .A4(new_n550_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n514_), .B1(new_n653_), .B2(new_n517_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n690_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT47), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT47), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n690_), .A2(new_n695_), .A3(new_n691_), .A4(new_n692_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(G1330gat));
  INV_X1    g496(.A(G50gat), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n471_), .A2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n599_), .A2(new_n470_), .A3(new_n652_), .ZN(new_n700_));
  AOI22_X1  g499(.A1(new_n649_), .A2(new_n699_), .B1(new_n698_), .B2(new_n700_), .ZN(G1331gat));
  NAND4_X1  g500(.A1(new_n608_), .A2(new_n303_), .A3(new_n597_), .A4(new_n581_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G57gat), .B1(new_n702_), .B2(new_n505_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n551_), .A2(new_n597_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n305_), .A2(new_n581_), .A3(new_n704_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n505_), .A2(G57gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n703_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT110), .ZN(G1332gat));
  OAI21_X1  g507(.A(G64gat), .B1(new_n702_), .B2(new_n417_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT48), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n417_), .A2(G64gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n710_), .B1(new_n705_), .B2(new_n711_), .ZN(G1333gat));
  OAI21_X1  g511(.A(G71gat), .B1(new_n702_), .B2(new_n517_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT49), .ZN(new_n714_));
  OR2_X1    g513(.A1(new_n517_), .A2(G71gat), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n714_), .B1(new_n705_), .B2(new_n715_), .ZN(G1334gat));
  OAI21_X1  g515(.A(G78gat), .B1(new_n702_), .B2(new_n471_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT50), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n471_), .A2(G78gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n705_), .B2(new_n719_), .ZN(G1335gat));
  AND2_X1   g519(.A1(new_n581_), .A2(new_n652_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n704_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n723_), .A2(new_n212_), .A3(new_n506_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n581_), .A2(new_n302_), .A3(new_n597_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(new_n506_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n724_), .B1(new_n728_), .B2(new_n212_), .ZN(G1336gat));
  OAI21_X1  g528(.A(new_n213_), .B1(new_n722_), .B2(new_n417_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT111), .Z(new_n731_));
  AND2_X1   g530(.A1(new_n613_), .A2(new_n208_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n726_), .B2(new_n732_), .ZN(G1337gat));
  NAND2_X1  g532(.A1(new_n726_), .A2(new_n550_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n550_), .A2(new_n202_), .ZN(new_n735_));
  AOI22_X1  g534(.A1(new_n734_), .A2(G99gat), .B1(new_n723_), .B2(new_n735_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n738_), .B(new_n739_), .Z(G1338gat));
  NAND3_X1  g539(.A1(new_n723_), .A2(new_n203_), .A3(new_n470_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n726_), .A2(new_n470_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(G106gat), .ZN(new_n743_));
  XOR2_X1   g542(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n744_));
  AND2_X1   g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n743_), .A2(new_n744_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n741_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g547(.A1(new_n664_), .A2(new_n303_), .A3(new_n597_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n272_), .A2(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT54), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n596_), .A2(new_n576_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT55), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n563_), .A2(new_n753_), .A3(new_n568_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT114), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT114), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n563_), .A2(new_n756_), .A3(new_n753_), .A4(new_n568_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n566_), .A2(KEYINPUT55), .A3(new_n567_), .A4(new_n557_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n560_), .A2(new_n562_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n755_), .A2(new_n757_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n573_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT56), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n762_), .A2(KEYINPUT56), .A3(new_n573_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n752_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n585_), .A2(new_n582_), .A3(new_n587_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n591_), .B1(new_n586_), .B2(new_n583_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n593_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n577_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n270_), .B1(new_n767_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT57), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n773_), .A2(KEYINPUT115), .A3(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT115), .ZN(new_n776_));
  INV_X1    g575(.A(new_n270_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n752_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n760_), .B1(new_n754_), .B2(KEYINPUT114), .ZN(new_n779_));
  AOI211_X1 g578(.A(new_n764_), .B(new_n575_), .C1(new_n779_), .C2(new_n757_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT56), .B1(new_n762_), .B2(new_n573_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n778_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n777_), .B1(new_n782_), .B2(new_n771_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n776_), .B1(new_n783_), .B2(KEYINPUT57), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(KEYINPUT57), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n770_), .A2(new_n576_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT116), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n770_), .A2(KEYINPUT116), .A3(new_n576_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n790_), .B1(new_n781_), .B2(new_n780_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT117), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT58), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n791_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n793_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n790_), .B(new_n795_), .C1(new_n781_), .C2(new_n780_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n794_), .A2(new_n272_), .A3(new_n796_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n775_), .A2(new_n784_), .A3(new_n785_), .A4(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n751_), .B1(new_n798_), .B2(new_n302_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n613_), .A2(new_n470_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n505_), .A2(new_n517_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(KEYINPUT59), .B1(new_n799_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n773_), .A2(new_n774_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n804_), .A2(new_n797_), .A3(new_n785_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n751_), .B1(new_n805_), .B2(new_n302_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n802_), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n807_), .A2(KEYINPUT118), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT59), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(KEYINPUT118), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n808_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(KEYINPUT119), .B1(new_n806_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n811_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n796_), .A2(new_n272_), .ZN(new_n815_));
  AOI22_X1  g614(.A1(new_n815_), .A2(new_n794_), .B1(KEYINPUT57), .B2(new_n783_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n303_), .B1(new_n816_), .B2(new_n804_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n813_), .B(new_n814_), .C1(new_n817_), .C2(new_n751_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n803_), .A2(new_n812_), .A3(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(G113gat), .B1(new_n819_), .B2(new_n597_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n799_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n807_), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n597_), .A2(G113gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n820_), .B1(new_n822_), .B2(new_n823_), .ZN(G1340gat));
  NAND4_X1  g623(.A1(new_n803_), .A2(new_n812_), .A3(new_n581_), .A4(new_n818_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(G120gat), .ZN(new_n826_));
  INV_X1    g625(.A(new_n822_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT60), .ZN(new_n828_));
  AOI21_X1  g627(.A(G120gat), .B1(new_n581_), .B2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n829_), .B1(new_n828_), .B2(G120gat), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n827_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n826_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT120), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n826_), .A2(KEYINPUT120), .A3(new_n831_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(G1341gat));
  OAI21_X1  g635(.A(G127gat), .B1(new_n819_), .B2(new_n302_), .ZN(new_n837_));
  OR2_X1    g636(.A1(new_n302_), .A2(G127gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n822_), .B2(new_n838_), .ZN(G1342gat));
  NAND4_X1  g638(.A1(new_n803_), .A2(new_n812_), .A3(new_n272_), .A4(new_n818_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(G134gat), .ZN(new_n841_));
  OR4_X1    g640(.A1(G134gat), .A2(new_n799_), .A3(new_n270_), .A4(new_n802_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT121), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n841_), .A2(KEYINPUT121), .A3(new_n842_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(G1343gat));
  NOR4_X1   g646(.A1(new_n613_), .A2(new_n505_), .A3(new_n471_), .A4(new_n550_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n821_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n596_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n581_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g653(.A1(new_n850_), .A2(new_n303_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT61), .B(G155gat), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1346gat));
  OR3_X1    g656(.A1(new_n849_), .A2(G162gat), .A3(new_n270_), .ZN(new_n858_));
  OAI21_X1  g657(.A(G162gat), .B1(new_n849_), .B2(new_n273_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(G1347gat));
  NAND2_X1  g659(.A1(new_n613_), .A2(new_n518_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n806_), .A2(new_n470_), .A3(new_n861_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT123), .ZN(new_n863_));
  XNOR2_X1  g662(.A(KEYINPUT22), .B(G169gat), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n863_), .A2(new_n596_), .A3(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n332_), .B1(new_n862_), .B2(new_n596_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n866_), .A2(KEYINPUT122), .A3(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n868_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n869_));
  AOI21_X1  g668(.A(KEYINPUT122), .B1(new_n866_), .B2(new_n867_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n865_), .B1(new_n869_), .B2(new_n870_), .ZN(G1348gat));
  NAND2_X1  g670(.A1(new_n581_), .A2(G176gat), .ZN(new_n872_));
  NOR4_X1   g671(.A1(new_n799_), .A2(new_n470_), .A3(new_n861_), .A4(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n863_), .A2(new_n581_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n873_), .B1(new_n874_), .B2(new_n333_), .ZN(G1349gat));
  NOR2_X1   g674(.A1(new_n302_), .A2(new_n349_), .ZN(new_n876_));
  NOR4_X1   g675(.A1(new_n799_), .A2(new_n302_), .A3(new_n470_), .A4(new_n861_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT124), .ZN(new_n878_));
  OR2_X1    g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(G183gat), .B1(new_n877_), .B2(new_n878_), .ZN(new_n880_));
  AOI22_X1  g679(.A1(new_n863_), .A2(new_n876_), .B1(new_n879_), .B2(new_n880_), .ZN(G1350gat));
  NAND2_X1  g680(.A1(new_n863_), .A2(new_n272_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(G190gat), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n863_), .A2(new_n777_), .A3(new_n345_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1351gat));
  NAND3_X1  g684(.A1(new_n470_), .A2(new_n505_), .A3(new_n517_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(KEYINPUT125), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n886_), .A2(KEYINPUT125), .ZN(new_n888_));
  AND3_X1   g687(.A1(new_n613_), .A2(new_n887_), .A3(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n821_), .A2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n597_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(new_n312_), .ZN(G1352gat));
  INV_X1    g691(.A(new_n890_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n581_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n311_), .A2(KEYINPUT126), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n894_), .B(new_n895_), .ZN(G1353gat));
  NAND2_X1  g695(.A1(new_n893_), .A2(new_n303_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n898_));
  AND2_X1   g697(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n897_), .A2(new_n898_), .A3(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n900_), .B1(new_n897_), .B2(new_n898_), .ZN(G1354gat));
  NOR3_X1   g700(.A1(new_n890_), .A2(new_n319_), .A3(new_n273_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n890_), .A2(new_n270_), .ZN(new_n903_));
  OR2_X1    g702(.A1(new_n903_), .A2(KEYINPUT127), .ZN(new_n904_));
  AOI21_X1  g703(.A(G218gat), .B1(new_n903_), .B2(KEYINPUT127), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n902_), .B1(new_n904_), .B2(new_n905_), .ZN(G1355gat));
endmodule


