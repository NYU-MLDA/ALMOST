//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 1 1 0 0 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n853_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n898_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  XOR2_X1   g002(.A(G211gat), .B(G218gat), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G197gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G204gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT89), .B(G204gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n207_), .B1(new_n208_), .B2(new_n206_), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n209_), .A2(KEYINPUT21), .ZN(new_n210_));
  INV_X1    g009(.A(G204gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G197gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT88), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n208_), .A2(new_n206_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  AND3_X1   g014(.A1(new_n215_), .A2(KEYINPUT90), .A3(KEYINPUT21), .ZN(new_n216_));
  AOI21_X1  g015(.A(KEYINPUT90), .B1(new_n215_), .B2(KEYINPUT21), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n205_), .B(new_n210_), .C1(new_n216_), .C2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n209_), .A2(KEYINPUT21), .A3(new_n204_), .ZN(new_n219_));
  XOR2_X1   g018(.A(KEYINPUT91), .B(KEYINPUT24), .Z(new_n220_));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT92), .ZN(new_n223_));
  INV_X1    g022(.A(G169gat), .ZN(new_n224_));
  INV_X1    g023(.A(G176gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT92), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n220_), .A2(new_n227_), .A3(new_n221_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n223_), .A2(new_n226_), .A3(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT25), .B(G183gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT26), .B(G190gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n220_), .A2(new_n226_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT23), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n233_), .A2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n229_), .A2(new_n232_), .A3(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT22), .B(G169gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(new_n225_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT80), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n221_), .B(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT93), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n235_), .B1(G183gat), .B2(G190gat), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT93), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n240_), .A2(new_n242_), .A3(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n244_), .A2(new_n245_), .A3(new_n247_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n218_), .A2(new_n219_), .A3(new_n238_), .A4(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(KEYINPUT97), .A3(KEYINPUT20), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n242_), .A2(KEYINPUT24), .A3(new_n226_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT81), .ZN(new_n252_));
  NAND2_X1  g051(.A1(KEYINPUT79), .A2(G190gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT78), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n253_), .A2(new_n254_), .A3(KEYINPUT26), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n253_), .B1(new_n254_), .B2(KEYINPUT26), .ZN(new_n256_));
  INV_X1    g055(.A(G190gat), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n254_), .B1(KEYINPUT26), .B2(new_n257_), .ZN(new_n258_));
  NOR3_X1   g057(.A1(new_n255_), .A2(new_n256_), .A3(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n236_), .B1(new_n259_), .B2(new_n230_), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n252_), .B(new_n260_), .C1(KEYINPUT24), .C2(new_n226_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n240_), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n262_), .A2(KEYINPUT82), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(KEYINPUT82), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n263_), .A2(new_n242_), .A3(new_n245_), .A4(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n261_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n218_), .A2(new_n219_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n250_), .A2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT97), .B1(new_n249_), .B2(KEYINPUT20), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n203_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT20), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n248_), .A2(KEYINPUT94), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT94), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n244_), .A2(new_n274_), .A3(new_n245_), .A4(new_n247_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(new_n238_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n272_), .B1(new_n277_), .B2(new_n267_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n261_), .A2(new_n265_), .A3(new_n218_), .A4(new_n219_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT98), .B1(new_n280_), .B2(new_n203_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT98), .ZN(new_n282_));
  INV_X1    g081(.A(new_n203_), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n278_), .A2(new_n282_), .A3(new_n283_), .A4(new_n279_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n271_), .A2(new_n281_), .A3(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G8gat), .B(G36gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G64gat), .B(G92gat), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n288_), .B(new_n289_), .Z(new_n290_));
  NAND2_X1  g089(.A1(new_n285_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT99), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n276_), .A2(new_n218_), .A3(new_n219_), .A4(new_n238_), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n294_), .A2(KEYINPUT95), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n272_), .B1(new_n294_), .B2(KEYINPUT95), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n295_), .A2(new_n296_), .A3(new_n283_), .A4(new_n268_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n290_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n280_), .A2(new_n203_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n297_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n300_), .A2(KEYINPUT27), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n285_), .A2(KEYINPUT99), .A3(new_n290_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n293_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G78gat), .B(G106gat), .ZN(new_n304_));
  INV_X1    g103(.A(G50gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306_));
  OR2_X1    g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307_));
  NOR2_X1   g106(.A1(G141gat), .A2(G148gat), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n308_), .B(KEYINPUT3), .Z(new_n309_));
  NAND2_X1  g108(.A1(G141gat), .A2(G148gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n310_), .B(KEYINPUT2), .Z(new_n311_));
  OAI211_X1 g110(.A(new_n306_), .B(new_n307_), .C1(new_n309_), .C2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n308_), .B(KEYINPUT86), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n306_), .A2(KEYINPUT1), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT87), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT87), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n306_), .A2(new_n316_), .A3(KEYINPUT1), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n317_), .A3(new_n307_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n306_), .A2(KEYINPUT1), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n313_), .B(new_n310_), .C1(new_n318_), .C2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n312_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT29), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n267_), .A2(new_n305_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n305_), .B1(new_n267_), .B2(new_n322_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n304_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n325_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n304_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n327_), .A2(new_n328_), .A3(new_n323_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n326_), .A2(new_n329_), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n321_), .A2(KEYINPUT29), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n331_), .A2(KEYINPUT28), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(KEYINPUT28), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G228gat), .A2(G233gat), .ZN(new_n334_));
  INV_X1    g133(.A(G22gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n332_), .A2(new_n333_), .A3(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n337_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n339_));
  OR2_X1    g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n330_), .A2(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n338_), .A2(new_n339_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(new_n326_), .A3(new_n329_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT84), .B(G99gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT31), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G15gat), .B(G43gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G227gat), .A2(G233gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G127gat), .B(G134gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(G113gat), .ZN(new_n352_));
  INV_X1    g151(.A(G120gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  OR2_X1    g153(.A1(new_n351_), .A2(G113gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n351_), .A2(G113gat), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n355_), .A2(G120gat), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n354_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT85), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n354_), .A2(KEYINPUT85), .A3(new_n357_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT83), .B(KEYINPUT30), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n360_), .A2(new_n361_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n362_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(G71gat), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n261_), .A2(new_n367_), .A3(new_n265_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n367_), .B1(new_n261_), .B2(new_n265_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n363_), .B(new_n366_), .C1(new_n369_), .C2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n370_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n366_), .A2(new_n363_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(new_n373_), .A3(new_n368_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n350_), .B1(new_n371_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n371_), .A2(new_n374_), .A3(new_n350_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n344_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n377_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n380_), .A2(new_n375_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(new_n341_), .A3(new_n343_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  AOI22_X1  g182(.A1(new_n360_), .A2(new_n361_), .B1(new_n320_), .B2(new_n312_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n358_), .A2(new_n321_), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT4), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n364_), .A2(new_n321_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT4), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n386_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G225gat), .A2(G233gat), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n384_), .A2(new_n385_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n391_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G1gat), .B(G29gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(G85gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT0), .ZN(new_n398_));
  INV_X1    g197(.A(G57gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n393_), .A2(new_n395_), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n400_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n391_), .B1(new_n386_), .B2(new_n389_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n395_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n402_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n401_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT100), .B(KEYINPUT27), .ZN(new_n408_));
  INV_X1    g207(.A(new_n300_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n298_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n408_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n303_), .A2(new_n383_), .A3(new_n407_), .A4(new_n411_), .ZN(new_n412_));
  NOR3_X1   g211(.A1(new_n384_), .A2(new_n391_), .A3(new_n385_), .ZN(new_n413_));
  AOI211_X1 g212(.A(new_n400_), .B(new_n413_), .C1(new_n390_), .C2(new_n391_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT33), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n401_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n410_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n393_), .A2(KEYINPUT33), .A3(new_n395_), .A4(new_n400_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n416_), .A2(new_n300_), .A3(new_n417_), .A4(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n298_), .A2(KEYINPUT32), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n285_), .A2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n297_), .A2(new_n299_), .A3(new_n420_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(new_n406_), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n419_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(new_n344_), .A3(new_n381_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n412_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT66), .ZN(new_n428_));
  INV_X1    g227(.A(G99gat), .ZN(new_n429_));
  INV_X1    g228(.A(G106gat), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT7), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G99gat), .A2(G106gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT6), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT6), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n435_), .A2(G99gat), .A3(G106gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT7), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n428_), .A2(new_n438_), .A3(new_n429_), .A4(new_n430_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n432_), .A2(new_n437_), .A3(new_n439_), .ZN(new_n440_));
  XOR2_X1   g239(.A(G85gat), .B(G92gat), .Z(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT8), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(KEYINPUT67), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n441_), .A2(KEYINPUT9), .ZN(new_n445_));
  XOR2_X1   g244(.A(KEYINPUT10), .B(G99gat), .Z(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n430_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(KEYINPUT65), .B(G85gat), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT9), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n448_), .A2(new_n449_), .A3(G92gat), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n445_), .A2(new_n447_), .A3(new_n437_), .A4(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT67), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n440_), .A2(new_n452_), .A3(new_n441_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT8), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n452_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n455_));
  OAI211_X1 g254(.A(new_n444_), .B(new_n451_), .C1(new_n454_), .C2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT68), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n442_), .A2(KEYINPUT67), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n459_), .A2(KEYINPUT8), .A3(new_n453_), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n460_), .A2(KEYINPUT68), .A3(new_n444_), .A4(new_n451_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G57gat), .B(G64gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT11), .ZN(new_n463_));
  XOR2_X1   g262(.A(G71gat), .B(G78gat), .Z(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  OR2_X1    g264(.A1(new_n462_), .A2(KEYINPUT11), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n458_), .A2(new_n461_), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT12), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n458_), .A2(new_n461_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n467_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G230gat), .A2(G233gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT64), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n467_), .B(KEYINPUT69), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n476_), .A2(KEYINPUT12), .A3(new_n456_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n470_), .A2(new_n473_), .A3(new_n475_), .A4(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n475_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n468_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n467_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n479_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n478_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G120gat), .B(G148gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT5), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(G176gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(G204gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n483_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n478_), .A2(new_n482_), .A3(new_n487_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT13), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n489_), .A2(KEYINPUT13), .A3(new_n490_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G113gat), .B(G141gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(new_n224_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(new_n206_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G15gat), .B(G22gat), .ZN(new_n500_));
  INV_X1    g299(.A(G1gat), .ZN(new_n501_));
  INV_X1    g300(.A(G8gat), .ZN(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT14), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n500_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G1gat), .B(G8gat), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n504_), .B(new_n505_), .Z(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  OR2_X1    g306(.A1(G29gat), .A2(G36gat), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT71), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G29gat), .A2(G36gat), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  AND2_X1   g310(.A1(G29gat), .A2(G36gat), .ZN(new_n512_));
  NOR2_X1   g311(.A1(G29gat), .A2(G36gat), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT71), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(G43gat), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n511_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n515_), .B1(new_n511_), .B2(new_n514_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n305_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n512_), .A2(new_n513_), .A3(KEYINPUT71), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n509_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n520_));
  OAI21_X1  g319(.A(G43gat), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n511_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n521_), .A2(G50gat), .A3(new_n522_), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n518_), .A2(KEYINPUT15), .A3(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(KEYINPUT15), .B1(new_n518_), .B2(new_n523_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n507_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT77), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G229gat), .A2(G233gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n518_), .A2(new_n523_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n507_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  OAI211_X1 g331(.A(KEYINPUT77), .B(new_n507_), .C1(new_n524_), .C2(new_n525_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n528_), .A2(new_n529_), .A3(new_n532_), .A4(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n529_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n506_), .B1(new_n523_), .B2(new_n518_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n535_), .B1(new_n531_), .B2(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n499_), .B1(new_n534_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n534_), .A2(new_n537_), .A3(new_n499_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n495_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n427_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G134gat), .B(G162gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G190gat), .B(G218gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n547_), .B(new_n548_), .Z(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n550_), .A2(KEYINPUT36), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n530_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n524_), .A2(new_n525_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n456_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n552_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G232gat), .A2(G233gat), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n557_), .B(KEYINPUT70), .Z(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT34), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT35), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(KEYINPUT72), .B1(new_n556_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n559_), .A2(new_n560_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n556_), .A2(new_n564_), .A3(new_n562_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT72), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n566_), .B(new_n561_), .C1(new_n552_), .C2(new_n555_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n563_), .A2(new_n565_), .A3(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n550_), .A2(KEYINPUT36), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n551_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n568_), .A2(new_n551_), .A3(new_n569_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n571_), .A2(KEYINPUT37), .A3(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT37), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n568_), .A2(new_n551_), .A3(new_n569_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n574_), .B1(new_n575_), .B2(new_n570_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n467_), .B(new_n506_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G231gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G127gat), .B(G155gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT16), .ZN(new_n581_));
  INV_X1    g380(.A(G183gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(G211gat), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT17), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n585_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n579_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT69), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n579_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT75), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n577_), .A2(new_n578_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n577_), .A2(new_n578_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n592_), .A2(KEYINPUT69), .A3(new_n593_), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n590_), .A2(new_n591_), .A3(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n591_), .B1(new_n590_), .B2(new_n594_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n586_), .B(KEYINPUT76), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n588_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n573_), .A2(new_n576_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n544_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n602_), .A2(new_n501_), .A3(new_n406_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT38), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT101), .ZN(new_n606_));
  INV_X1    g405(.A(new_n599_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n575_), .A2(new_n570_), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n608_), .A2(KEYINPUT102), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(KEYINPUT102), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n607_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n544_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(G1gat), .B1(new_n614_), .B2(new_n407_), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n606_), .B(new_n615_), .C1(KEYINPUT38), .C2(new_n604_), .ZN(G1324gat));
  INV_X1    g415(.A(new_n544_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n303_), .A2(new_n411_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n617_), .A2(KEYINPUT103), .A3(new_n618_), .A4(new_n611_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n611_), .A2(new_n427_), .A3(new_n543_), .A4(new_n618_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT103), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n619_), .A2(new_n622_), .A3(G8gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT39), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n602_), .A2(new_n502_), .A3(new_n618_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT40), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n624_), .A2(KEYINPUT40), .A3(new_n625_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1325gat));
  INV_X1    g429(.A(G15gat), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n631_), .B1(new_n613_), .B2(new_n378_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT41), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n602_), .A2(new_n631_), .A3(new_n378_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(G1326gat));
  INV_X1    g434(.A(new_n344_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n602_), .A2(new_n335_), .A3(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n613_), .A2(new_n636_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(G22gat), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n639_), .A2(KEYINPUT104), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(KEYINPUT104), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n640_), .A2(KEYINPUT42), .A3(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT42), .B1(new_n640_), .B2(new_n641_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n637_), .B1(new_n642_), .B2(new_n643_), .ZN(G1327gat));
  INV_X1    g443(.A(new_n608_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n544_), .A2(new_n645_), .A3(new_n599_), .ZN(new_n646_));
  AOI21_X1  g445(.A(G29gat), .B1(new_n646_), .B2(new_n406_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n573_), .A2(new_n576_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n427_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT43), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n427_), .A2(new_n651_), .A3(new_n648_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n653_), .A2(KEYINPUT44), .A3(new_n543_), .A4(new_n607_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n654_), .A2(G29gat), .A3(new_n406_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n427_), .A2(new_n651_), .A3(new_n648_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n651_), .B1(new_n427_), .B2(new_n648_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n543_), .B(new_n607_), .C1(new_n657_), .C2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n647_), .B1(new_n656_), .B2(new_n661_), .ZN(G1328gat));
  NAND3_X1  g461(.A1(new_n661_), .A2(new_n654_), .A3(new_n618_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(G36gat), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT106), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT46), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n665_), .A2(KEYINPUT46), .ZN(new_n667_));
  INV_X1    g466(.A(G36gat), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n617_), .A2(new_n668_), .A3(new_n608_), .A4(new_n607_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT105), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n618_), .A2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n303_), .A2(KEYINPUT105), .A3(new_n411_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(KEYINPUT45), .B1(new_n669_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT45), .ZN(new_n675_));
  INV_X1    g474(.A(new_n673_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n646_), .A2(new_n675_), .A3(new_n668_), .A4(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n674_), .A2(new_n677_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n664_), .A2(new_n666_), .A3(new_n667_), .A4(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n618_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n668_), .B1(new_n681_), .B2(new_n654_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n674_), .A2(new_n677_), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n665_), .B(KEYINPUT46), .C1(new_n682_), .C2(new_n683_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n679_), .A2(new_n684_), .ZN(G1329gat));
  NAND4_X1  g484(.A1(new_n661_), .A2(new_n654_), .A3(G43gat), .A4(new_n378_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n646_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n515_), .B1(new_n687_), .B2(new_n381_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g489(.A1(new_n661_), .A2(new_n654_), .A3(G50gat), .A4(new_n636_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n305_), .B1(new_n687_), .B2(new_n344_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1331gat));
  NAND3_X1  g492(.A1(new_n427_), .A2(new_n542_), .A3(new_n495_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n694_), .A2(new_n601_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G57gat), .B1(new_n695_), .B2(new_n406_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n694_), .A2(new_n612_), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n697_), .A2(KEYINPUT107), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(KEYINPUT107), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n407_), .A2(new_n399_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n696_), .B1(new_n700_), .B2(new_n701_), .ZN(G1332gat));
  INV_X1    g501(.A(G64gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n695_), .A2(new_n703_), .A3(new_n676_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n698_), .A2(new_n676_), .A3(new_n699_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT48), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n705_), .A2(new_n706_), .A3(G64gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n705_), .B2(G64gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n704_), .B1(new_n707_), .B2(new_n708_), .ZN(G1333gat));
  NAND2_X1  g508(.A1(new_n378_), .A2(new_n367_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT108), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n695_), .A2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n698_), .A2(new_n378_), .A3(new_n699_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT49), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n713_), .A2(new_n714_), .A3(G71gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n713_), .B2(G71gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(G1334gat));
  INV_X1    g516(.A(G78gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n695_), .A2(new_n718_), .A3(new_n636_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n698_), .A2(new_n636_), .A3(new_n699_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT50), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n720_), .A2(new_n721_), .A3(G78gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n720_), .B2(G78gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n719_), .B1(new_n722_), .B2(new_n723_), .ZN(G1335gat));
  NOR3_X1   g523(.A1(new_n694_), .A2(new_n645_), .A3(new_n599_), .ZN(new_n725_));
  AOI21_X1  g524(.A(G85gat), .B1(new_n725_), .B2(new_n406_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT109), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n727_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n650_), .A2(KEYINPUT109), .A3(new_n652_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n495_), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n730_), .A2(new_n541_), .A3(new_n599_), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n728_), .A2(new_n729_), .A3(new_n731_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n406_), .A2(new_n448_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n726_), .B1(new_n732_), .B2(new_n733_), .ZN(G1336gat));
  AOI21_X1  g533(.A(G92gat), .B1(new_n725_), .B2(new_n618_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n676_), .A2(G92gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n732_), .B2(new_n736_), .ZN(G1337gat));
  NAND4_X1  g536(.A1(new_n728_), .A2(new_n729_), .A3(new_n378_), .A4(new_n731_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n378_), .A2(new_n446_), .ZN(new_n739_));
  AOI22_X1  g538(.A1(new_n738_), .A2(G99gat), .B1(new_n725_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n741_), .A2(KEYINPUT51), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(KEYINPUT51), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n740_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n742_), .B1(new_n740_), .B2(new_n743_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1338gat));
  NAND3_X1  g545(.A1(new_n725_), .A2(new_n430_), .A3(new_n636_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n653_), .A2(new_n636_), .A3(new_n731_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT52), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n748_), .A2(new_n749_), .A3(G106gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n748_), .B2(G106gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n747_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT53), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT53), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n754_), .B(new_n747_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1339gat));
  XNOR2_X1  g555(.A(KEYINPUT111), .B(KEYINPUT112), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT54), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n600_), .A2(new_n542_), .A3(new_n730_), .A4(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n758_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n573_), .A2(new_n576_), .A3(new_n542_), .A4(new_n599_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(new_n495_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n759_), .A2(new_n762_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n528_), .A2(new_n535_), .A3(new_n532_), .A4(new_n533_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n529_), .B1(new_n531_), .B2(new_n536_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n764_), .A2(new_n498_), .A3(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n490_), .A2(new_n540_), .A3(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n470_), .A2(new_n473_), .A3(new_n477_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n479_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n769_), .A2(KEYINPUT55), .A3(new_n478_), .ZN(new_n770_));
  OR2_X1    g569(.A1(new_n478_), .A2(KEYINPUT55), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n770_), .A2(new_n488_), .A3(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT56), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n775_), .B1(new_n768_), .B2(new_n479_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n487_), .B1(new_n776_), .B2(new_n478_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n777_), .A2(KEYINPUT56), .A3(new_n771_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n767_), .B1(new_n774_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT114), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT58), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n767_), .ZN(new_n782_));
  AND4_X1   g581(.A1(KEYINPUT56), .A2(new_n770_), .A3(new_n488_), .A4(new_n771_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT56), .B1(new_n777_), .B2(new_n771_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n782_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT58), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n785_), .A2(KEYINPUT114), .A3(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n781_), .A2(new_n787_), .A3(new_n648_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT57), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n491_), .A2(new_n540_), .A3(new_n766_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n540_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n490_), .B1(new_n791_), .B2(new_n538_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n541_), .A2(KEYINPUT113), .A3(new_n490_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n774_), .A2(new_n778_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n790_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n789_), .B1(new_n799_), .B2(new_n608_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n796_), .B1(new_n774_), .B2(new_n778_), .ZN(new_n801_));
  OAI211_X1 g600(.A(KEYINPUT57), .B(new_n645_), .C1(new_n801_), .C2(new_n790_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n788_), .A2(new_n800_), .A3(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n763_), .B1(new_n803_), .B2(new_n607_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n379_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n680_), .A2(new_n805_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n804_), .A2(new_n407_), .A3(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(G113gat), .B1(new_n807_), .B2(new_n541_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT59), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n803_), .A2(new_n607_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n763_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n407_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n806_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n809_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NOR4_X1   g613(.A1(new_n804_), .A2(KEYINPUT59), .A3(new_n407_), .A4(new_n806_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n541_), .A2(G113gat), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(KEYINPUT115), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n808_), .B1(new_n816_), .B2(new_n818_), .ZN(G1340gat));
  OAI21_X1  g618(.A(new_n353_), .B1(new_n730_), .B2(KEYINPUT60), .ZN(new_n820_));
  OAI21_X1  g619(.A(KEYINPUT116), .B1(new_n353_), .B2(KEYINPUT60), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n807_), .B(new_n822_), .C1(new_n823_), .C2(new_n820_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n814_), .A2(new_n815_), .A3(new_n730_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n825_), .B2(new_n353_), .ZN(G1341gat));
  INV_X1    g625(.A(G127gat), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n607_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n814_), .A2(new_n815_), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(G127gat), .B1(new_n807_), .B2(new_n599_), .ZN(new_n831_));
  OAI21_X1  g630(.A(KEYINPUT117), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n812_), .A2(new_n813_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT59), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n807_), .A2(new_n809_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n834_), .A2(new_n835_), .A3(new_n828_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n837_));
  INV_X1    g636(.A(new_n831_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n836_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n832_), .A2(new_n839_), .ZN(G1342gat));
  INV_X1    g639(.A(G134gat), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n609_), .A2(new_n610_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n841_), .B1(new_n833_), .B2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT118), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n834_), .A2(G134gat), .A3(new_n835_), .A4(new_n648_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n847_), .B(new_n841_), .C1(new_n833_), .C2(new_n843_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n845_), .A2(new_n846_), .A3(new_n848_), .ZN(G1343gat));
  NOR4_X1   g648(.A1(new_n804_), .A2(new_n407_), .A3(new_n382_), .A4(new_n676_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n541_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n495_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g653(.A(KEYINPUT119), .B(KEYINPUT120), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  XOR2_X1   g655(.A(KEYINPUT61), .B(G155gat), .Z(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n850_), .A2(new_n599_), .A3(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n858_), .B1(new_n850_), .B2(new_n599_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n856_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n812_), .A2(new_n381_), .A3(new_n636_), .A4(new_n673_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n857_), .B1(new_n863_), .B2(new_n607_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n864_), .A2(new_n855_), .A3(new_n859_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n862_), .A2(new_n865_), .ZN(G1346gat));
  AOI21_X1  g665(.A(G162gat), .B1(new_n850_), .B2(new_n842_), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n648_), .A2(G162gat), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n850_), .B2(new_n868_), .ZN(G1347gat));
  NOR2_X1   g668(.A1(new_n804_), .A2(new_n636_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n671_), .A2(new_n407_), .A3(new_n378_), .A4(new_n672_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(KEYINPUT121), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n870_), .A2(new_n541_), .A3(new_n872_), .ZN(new_n873_));
  XOR2_X1   g672(.A(KEYINPUT122), .B(KEYINPUT62), .Z(new_n874_));
  AND3_X1   g673(.A1(new_n873_), .A2(G169gat), .A3(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n873_), .B2(G169gat), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n870_), .A2(new_n872_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n541_), .A2(new_n239_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(KEYINPUT123), .ZN(new_n879_));
  OAI22_X1  g678(.A1(new_n875_), .A2(new_n876_), .B1(new_n877_), .B2(new_n879_), .ZN(G1348gat));
  NAND2_X1  g679(.A1(new_n810_), .A2(new_n811_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n881_), .A2(KEYINPUT125), .A3(new_n344_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT125), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n804_), .B2(new_n636_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n730_), .A2(new_n225_), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n882_), .A2(new_n884_), .A3(new_n872_), .A4(new_n885_), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n886_), .A2(KEYINPUT126), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(KEYINPUT126), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n870_), .A2(new_n495_), .A3(new_n872_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n225_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT124), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT124), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n889_), .A2(new_n892_), .A3(new_n225_), .ZN(new_n893_));
  AOI22_X1  g692(.A1(new_n887_), .A2(new_n888_), .B1(new_n891_), .B2(new_n893_), .ZN(G1349gat));
  NOR3_X1   g693(.A1(new_n877_), .A2(new_n230_), .A3(new_n607_), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n882_), .A2(new_n884_), .A3(new_n599_), .A4(new_n872_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n895_), .B1(new_n582_), .B2(new_n896_), .ZN(G1350gat));
  AND2_X1   g696(.A1(new_n573_), .A2(new_n576_), .ZN(new_n898_));
  OAI21_X1  g697(.A(G190gat), .B1(new_n877_), .B2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n842_), .A2(new_n231_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n877_), .B2(new_n900_), .ZN(G1351gat));
  NOR2_X1   g700(.A1(new_n804_), .A2(new_n382_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n673_), .A2(new_n406_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n542_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(new_n206_), .ZN(G1352gat));
  INV_X1    g705(.A(new_n904_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(new_n495_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(G204gat), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n909_), .B1(new_n908_), .B2(new_n208_), .ZN(G1353gat));
  AOI21_X1  g709(.A(new_n607_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n911_));
  XOR2_X1   g710(.A(new_n911_), .B(KEYINPUT127), .Z(new_n912_));
  NAND2_X1  g711(.A1(new_n907_), .A2(new_n912_), .ZN(new_n913_));
  OR2_X1    g712(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n913_), .B(new_n914_), .ZN(G1354gat));
  AND3_X1   g714(.A1(new_n907_), .A2(G218gat), .A3(new_n648_), .ZN(new_n916_));
  AOI21_X1  g715(.A(G218gat), .B1(new_n907_), .B2(new_n842_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1355gat));
endmodule


