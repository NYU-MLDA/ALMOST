//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 0 1 0 0 0 0 1 0 1 0 0 1 0 1 0 1 0 0 0 1 0 1 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n926_, new_n927_, new_n928_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_;
  INV_X1    g000(.A(KEYINPUT29), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT82), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT82), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n209_), .B1(G155gat), .B2(G162gat), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT1), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n211_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT83), .ZN(new_n216_));
  OAI22_X1  g015(.A1(new_n215_), .A2(new_n216_), .B1(KEYINPUT1), .B2(new_n213_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n208_), .A2(new_n210_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n218_), .B1(KEYINPUT1), .B2(new_n213_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n219_), .A2(KEYINPUT83), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n206_), .B1(new_n217_), .B2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n205_), .B(KEYINPUT3), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n203_), .B(KEYINPUT2), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n218_), .A2(new_n214_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n202_), .B1(new_n221_), .B2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G211gat), .B(G218gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT84), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G197gat), .B(G204gat), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n229_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n232_), .A2(KEYINPUT21), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(KEYINPUT21), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n229_), .A2(new_n231_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  OAI211_X1 g035(.A(G228gat), .B(G233gat), .C1(new_n227_), .C2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n236_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G228gat), .A2(G233gat), .ZN(new_n239_));
  AOI22_X1  g038(.A1(new_n219_), .A2(KEYINPUT83), .B1(new_n212_), .B2(new_n214_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n240_), .B1(KEYINPUT83), .B2(new_n219_), .ZN(new_n241_));
  AOI22_X1  g040(.A1(new_n241_), .A2(new_n206_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n238_), .B(new_n239_), .C1(new_n242_), .C2(new_n202_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G78gat), .B(G106gat), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n237_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n245_), .B1(new_n237_), .B2(new_n243_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT28), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n242_), .A2(new_n249_), .A3(new_n202_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n221_), .A2(new_n226_), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT28), .B1(new_n251_), .B2(KEYINPUT29), .ZN(new_n252_));
  XOR2_X1   g051(.A(G22gat), .B(G50gat), .Z(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n250_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n254_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT85), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n246_), .B(new_n248_), .C1(new_n257_), .C2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n250_), .A2(new_n252_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(new_n253_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n250_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n246_), .A2(new_n258_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n246_), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n263_), .B(new_n264_), .C1(new_n265_), .C2(new_n247_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n259_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(G127gat), .B(G134gat), .Z(new_n269_));
  XNOR2_X1  g068(.A(G113gat), .B(G120gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  XOR2_X1   g070(.A(new_n271_), .B(KEYINPUT31), .Z(new_n272_));
  NAND2_X1  g071(.A1(G227gat), .A2(G233gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(G15gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(G71gat), .B(G99gat), .Z(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT80), .B(G43gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G183gat), .A2(G190gat), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT23), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT76), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n279_), .B(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n281_), .B1(new_n283_), .B2(new_n280_), .ZN(new_n284_));
  OR3_X1    g083(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT77), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n284_), .A2(KEYINPUT77), .A3(new_n285_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT25), .B(G183gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT26), .B(G190gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT75), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n288_), .A2(new_n289_), .A3(new_n292_), .A4(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT22), .B(G169gat), .ZN(new_n299_));
  INV_X1    g098(.A(G176gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n294_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT78), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n283_), .A2(KEYINPUT23), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n304_), .B1(KEYINPUT23), .B2(new_n279_), .ZN(new_n305_));
  OR2_X1    g104(.A1(G183gat), .A2(G190gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n303_), .A2(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(KEYINPUT79), .B(KEYINPUT30), .Z(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n298_), .A2(new_n308_), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n310_), .B1(new_n298_), .B2(new_n308_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n278_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n313_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n278_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n315_), .A2(new_n311_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n314_), .A2(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n272_), .B1(new_n318_), .B2(KEYINPUT81), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT81), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n314_), .A2(new_n317_), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n314_), .A2(new_n317_), .A3(new_n320_), .A4(new_n272_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n268_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT92), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n271_), .B(KEYINPUT91), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n242_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(KEYINPUT92), .B1(new_n251_), .B2(new_n271_), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n327_), .A2(new_n221_), .A3(new_n226_), .ZN(new_n330_));
  OAI211_X1 g129(.A(new_n328_), .B(KEYINPUT4), .C1(new_n329_), .C2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G225gat), .A2(G233gat), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT4), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n251_), .A2(new_n334_), .A3(new_n271_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n331_), .A2(new_n333_), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT93), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT93), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n331_), .A2(new_n338_), .A3(new_n333_), .A4(new_n335_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n329_), .A2(new_n330_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n328_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(new_n332_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G1gat), .B(G29gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT0), .ZN(new_n346_));
  INV_X1    g145(.A(G57gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(G85gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n340_), .A2(new_n344_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT33), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n340_), .A2(KEYINPUT33), .A3(new_n344_), .A4(new_n351_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n331_), .A2(new_n335_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n332_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n333_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n351_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n298_), .A2(new_n236_), .A3(new_n308_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n284_), .A2(new_n306_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT88), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n294_), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n364_), .A2(KEYINPUT87), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(KEYINPUT87), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(new_n366_), .A3(new_n301_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n296_), .A2(new_n293_), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n369_), .A2(new_n285_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n305_), .A2(new_n292_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT86), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n305_), .A2(KEYINPUT86), .A3(new_n292_), .A4(new_n370_), .ZN(new_n374_));
  AOI22_X1  g173(.A1(new_n363_), .A2(new_n368_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  OAI211_X1 g174(.A(KEYINPUT20), .B(new_n360_), .C1(new_n375_), .C2(new_n236_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G226gat), .A2(G233gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT19), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n375_), .A2(new_n236_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n298_), .A2(new_n308_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n238_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n378_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n380_), .A2(new_n382_), .A3(KEYINPUT20), .A4(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n379_), .A2(new_n384_), .ZN(new_n385_));
  XOR2_X1   g184(.A(G64gat), .B(G92gat), .Z(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT90), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G8gat), .B(G36gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n385_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n391_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n379_), .A2(new_n393_), .A3(new_n384_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n359_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n354_), .A2(new_n355_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT32), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n391_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT94), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(new_n379_), .A3(new_n384_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT95), .B(KEYINPUT20), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n361_), .B(KEYINPUT88), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n403_), .A2(new_n367_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n236_), .A2(new_n371_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n402_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n382_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n378_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n408_), .B1(new_n378_), .B2(new_n376_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(new_n399_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n401_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n340_), .A2(new_n344_), .A3(new_n351_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n351_), .B1(new_n340_), .B2(new_n344_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n412_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n325_), .B1(new_n397_), .B2(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n413_), .A2(new_n414_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n267_), .A2(new_n324_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n259_), .A2(new_n322_), .A3(new_n266_), .A4(new_n323_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n409_), .A2(new_n391_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT96), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n394_), .A2(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n379_), .A2(new_n384_), .A3(KEYINPUT96), .A4(new_n393_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n421_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT27), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT27), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n392_), .A2(new_n427_), .A3(new_n394_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n417_), .A2(new_n420_), .A3(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n416_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT67), .ZN(new_n432_));
  NOR2_X1   g231(.A1(G99gat), .A2(G106gat), .ZN(new_n433_));
  NOR2_X1   g232(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G99gat), .A2(G106gat), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT6), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n439_));
  OAI22_X1  g238(.A1(KEYINPUT65), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n435_), .A2(new_n438_), .A3(new_n439_), .A4(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(G92gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n349_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G85gat), .A2(G92gat), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n441_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT8), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G57gat), .B(G64gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G71gat), .B(G78gat), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(new_n450_), .A3(KEYINPUT11), .ZN(new_n451_));
  XOR2_X1   g250(.A(G71gat), .B(G78gat), .Z(new_n452_));
  INV_X1    g251(.A(G64gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(G57gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n347_), .A2(G64gat), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(new_n455_), .A3(KEYINPUT11), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n452_), .A2(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n449_), .A2(KEYINPUT11), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n451_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(G85gat), .B1(KEYINPUT64), .B2(G92gat), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT64), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n460_), .B1(new_n461_), .B2(new_n442_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT9), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  OR2_X1    g263(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n465_));
  INV_X1    g264(.A(G106gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n438_), .A2(new_n439_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n443_), .A2(new_n461_), .A3(KEYINPUT9), .A4(new_n444_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n464_), .A2(new_n468_), .A3(new_n469_), .A4(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n441_), .A2(KEYINPUT8), .A3(new_n445_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n448_), .A2(new_n459_), .A3(new_n471_), .A4(new_n472_), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n473_), .A2(KEYINPUT66), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n448_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n459_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n473_), .A2(KEYINPUT66), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n474_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(G230gat), .ZN(new_n480_));
  INV_X1    g279(.A(G233gat), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n479_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n482_), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n473_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT12), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n475_), .A2(new_n486_), .A3(new_n476_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n486_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n485_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G120gat), .B(G148gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT5), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G176gat), .B(G204gat), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n491_), .B(new_n492_), .Z(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n483_), .A2(new_n489_), .A3(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n494_), .B1(new_n483_), .B2(new_n489_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n432_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n483_), .A2(new_n489_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(new_n493_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(KEYINPUT67), .A3(new_n495_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT13), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n498_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n502_), .B1(new_n498_), .B2(new_n501_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G113gat), .B(G141gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G169gat), .B(G197gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G229gat), .A2(G233gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G29gat), .B(G36gat), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT69), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  XOR2_X1   g313(.A(G43gat), .B(G50gat), .Z(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G15gat), .B(G22gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT72), .B(G1gat), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n518_), .A2(G8gat), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT14), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n517_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(G1gat), .B(G8gat), .Z(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n522_), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n517_), .B(new_n524_), .C1(new_n519_), .C2(new_n520_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n516_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT73), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n516_), .A2(new_n526_), .A3(KEYINPUT73), .ZN(new_n530_));
  INV_X1    g329(.A(new_n526_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n515_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n514_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n512_), .B(KEYINPUT69), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n515_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT15), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT15), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n533_), .A2(new_n535_), .A3(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n531_), .A2(new_n537_), .A3(new_n539_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n529_), .A2(new_n530_), .B1(new_n540_), .B2(KEYINPUT74), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT74), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n531_), .A2(new_n537_), .A3(new_n542_), .A4(new_n539_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n511_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n516_), .A2(new_n526_), .ZN(new_n545_));
  AOI211_X1 g344(.A(new_n510_), .B(new_n545_), .C1(new_n529_), .C2(new_n530_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n509_), .B1(new_n544_), .B2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n529_), .A2(new_n530_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n540_), .A2(KEYINPUT74), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n548_), .A2(new_n549_), .A3(new_n543_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n510_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n546_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(new_n552_), .A3(new_n508_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n547_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n505_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n537_), .A2(new_n475_), .A3(new_n539_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n536_), .A2(new_n475_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G232gat), .A2(G233gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT34), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT35), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n558_), .A2(new_n559_), .A3(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n562_), .A2(new_n563_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n566_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n558_), .A2(new_n568_), .A3(new_n559_), .A4(new_n564_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G190gat), .B(G218gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G134gat), .B(G162gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n572_), .A2(KEYINPUT36), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n567_), .A2(new_n569_), .A3(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n572_), .B(KEYINPUT36), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n575_), .B1(new_n567_), .B2(new_n569_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n574_), .B1(KEYINPUT71), .B2(new_n576_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n576_), .A2(KEYINPUT71), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n579_), .A2(KEYINPUT97), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(KEYINPUT97), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(G127gat), .B(G155gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT16), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G183gat), .B(G211gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT17), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G231gat), .A2(G233gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n459_), .B(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(new_n526_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n587_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT17), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n590_), .B1(new_n592_), .B2(new_n586_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n582_), .A2(new_n594_), .ZN(new_n595_));
  NOR3_X1   g394(.A1(new_n431_), .A2(new_n557_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n417_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(G1gat), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n496_), .A2(new_n497_), .A3(new_n432_), .ZN(new_n600_));
  AOI21_X1  g399(.A(KEYINPUT67), .B1(new_n500_), .B2(new_n495_), .ZN(new_n601_));
  OAI21_X1  g400(.A(KEYINPUT13), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n498_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT68), .ZN(new_n605_));
  OAI21_X1  g404(.A(KEYINPUT37), .B1(new_n574_), .B2(new_n576_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT70), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT37), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n577_), .A2(new_n609_), .A3(new_n578_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n606_), .A2(new_n607_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n608_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(new_n594_), .ZN(new_n613_));
  NOR4_X1   g412(.A1(new_n431_), .A2(new_n555_), .A3(new_n605_), .A4(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n518_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n614_), .A2(new_n597_), .A3(new_n615_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n616_), .A2(KEYINPUT38), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(KEYINPUT38), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n599_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT98), .ZN(G1324gat));
  INV_X1    g419(.A(G8gat), .ZN(new_n621_));
  INV_X1    g420(.A(new_n429_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n614_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT39), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n596_), .A2(new_n622_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n624_), .B1(new_n625_), .B2(G8gat), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n626_), .A2(KEYINPUT99), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n625_), .A2(new_n624_), .A3(G8gat), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n628_), .B1(new_n626_), .B2(KEYINPUT99), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n623_), .B1(new_n627_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT40), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  OAI211_X1 g431(.A(KEYINPUT40), .B(new_n623_), .C1(new_n627_), .C2(new_n629_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(G1325gat));
  INV_X1    g433(.A(new_n324_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n596_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(G15gat), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n637_), .A2(KEYINPUT41), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(KEYINPUT41), .ZN(new_n639_));
  INV_X1    g438(.A(G15gat), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n614_), .A2(new_n640_), .A3(new_n635_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n638_), .A2(new_n639_), .A3(new_n641_), .ZN(G1326gat));
  INV_X1    g441(.A(G22gat), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n643_), .B1(new_n596_), .B2(new_n267_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT42), .Z(new_n645_));
  NAND3_X1  g444(.A1(new_n614_), .A2(new_n643_), .A3(new_n267_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(G1327gat));
  INV_X1    g446(.A(new_n325_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n396_), .A2(new_n355_), .ZN(new_n649_));
  AOI22_X1  g448(.A1(new_n337_), .A2(new_n339_), .B1(new_n332_), .B2(new_n343_), .ZN(new_n650_));
  AOI21_X1  g449(.A(KEYINPUT33), .B1(new_n650_), .B2(new_n351_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n649_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n340_), .A2(new_n344_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(new_n350_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n411_), .B1(new_n654_), .B2(new_n352_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n648_), .B1(new_n652_), .B2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n417_), .A2(new_n420_), .A3(new_n429_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n659_));
  INV_X1    g458(.A(new_n579_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n594_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT101), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n658_), .A2(new_n659_), .A3(new_n556_), .A4(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n556_), .ZN(new_n665_));
  OAI21_X1  g464(.A(KEYINPUT102), .B1(new_n431_), .B2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(G29gat), .B1(new_n668_), .B2(new_n597_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n612_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n670_), .B1(new_n416_), .B2(new_n430_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT43), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT43), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n673_), .B(new_n670_), .C1(new_n416_), .C2(new_n430_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n556_), .A2(new_n661_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT100), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n675_), .A2(KEYINPUT44), .A3(new_n678_), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n679_), .A2(G29gat), .A3(new_n597_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n675_), .A2(new_n678_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n669_), .B1(new_n680_), .B2(new_n683_), .ZN(G1328gat));
  NOR2_X1   g483(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n429_), .A2(G36gat), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n664_), .A2(new_n666_), .A3(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT45), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT45), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n664_), .A2(new_n666_), .A3(new_n689_), .A4(new_n686_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n685_), .B1(new_n688_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT103), .ZN(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT104), .B1(new_n692_), .B2(KEYINPUT46), .ZN(new_n693_));
  AOI21_X1  g492(.A(KEYINPUT44), .B1(new_n675_), .B2(new_n678_), .ZN(new_n694_));
  AOI211_X1 g493(.A(new_n682_), .B(new_n677_), .C1(new_n672_), .C2(new_n674_), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n694_), .A2(new_n695_), .A3(new_n429_), .ZN(new_n696_));
  INV_X1    g495(.A(G36gat), .ZN(new_n697_));
  OAI211_X1 g496(.A(new_n691_), .B(new_n693_), .C1(new_n696_), .C2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n683_), .A2(new_n622_), .A3(new_n679_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(G36gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n693_), .B1(new_n701_), .B2(new_n691_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n699_), .A2(new_n702_), .ZN(G1329gat));
  NAND2_X1  g502(.A1(new_n683_), .A2(new_n679_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n635_), .A2(G43gat), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n667_), .A2(new_n324_), .ZN(new_n706_));
  OAI22_X1  g505(.A1(new_n704_), .A2(new_n705_), .B1(G43gat), .B2(new_n706_), .ZN(new_n707_));
  XOR2_X1   g506(.A(KEYINPUT105), .B(KEYINPUT47), .Z(new_n708_));
  XNOR2_X1  g507(.A(new_n707_), .B(new_n708_), .ZN(G1330gat));
  OR3_X1    g508(.A1(new_n667_), .A2(G50gat), .A3(new_n268_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n683_), .A2(new_n267_), .A3(new_n679_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n711_), .A2(KEYINPUT106), .ZN(new_n712_));
  OAI21_X1  g511(.A(G50gat), .B1(new_n711_), .B2(KEYINPUT106), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n710_), .B1(new_n712_), .B2(new_n713_), .ZN(G1331gat));
  INV_X1    g513(.A(new_n605_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n431_), .A2(new_n554_), .A3(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n716_), .A2(new_n594_), .A3(new_n582_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G57gat), .B1(new_n717_), .B2(new_n417_), .ZN(new_n718_));
  NOR4_X1   g517(.A1(new_n431_), .A2(new_n554_), .A3(new_n604_), .A4(new_n613_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n719_), .A2(new_n347_), .A3(new_n597_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1332gat));
  OAI21_X1  g520(.A(G64gat), .B1(new_n717_), .B2(new_n429_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT48), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n719_), .A2(new_n453_), .A3(new_n622_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1333gat));
  OAI21_X1  g524(.A(G71gat), .B1(new_n717_), .B2(new_n324_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT49), .ZN(new_n727_));
  INV_X1    g526(.A(G71gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n719_), .A2(new_n728_), .A3(new_n635_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1334gat));
  OAI21_X1  g529(.A(G78gat), .B1(new_n717_), .B2(new_n268_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT50), .ZN(new_n732_));
  INV_X1    g531(.A(G78gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n719_), .A2(new_n733_), .A3(new_n267_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(G1335gat));
  AND2_X1   g534(.A1(new_n716_), .A2(new_n663_), .ZN(new_n736_));
  AOI21_X1  g535(.A(G85gat), .B1(new_n736_), .B2(new_n597_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT107), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n737_), .A2(KEYINPUT107), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n505_), .A2(new_n661_), .A3(new_n555_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n672_), .B2(new_n674_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n743_), .A2(new_n349_), .A3(new_n417_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n739_), .A2(new_n740_), .A3(new_n744_), .ZN(G1336gat));
  OAI21_X1  g544(.A(G92gat), .B1(new_n743_), .B2(new_n429_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n736_), .A2(new_n442_), .A3(new_n622_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1337gat));
  AND3_X1   g547(.A1(new_n635_), .A2(new_n465_), .A3(new_n467_), .ZN(new_n749_));
  AOI21_X1  g548(.A(KEYINPUT109), .B1(new_n736_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(G99gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n742_), .B2(new_n635_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n752_), .A2(KEYINPUT108), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n752_), .A2(KEYINPUT108), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n750_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT51), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n757_), .B(new_n750_), .C1(new_n753_), .C2(new_n754_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1338gat));
  NAND3_X1  g558(.A1(new_n736_), .A2(new_n466_), .A3(new_n267_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n742_), .A2(new_n267_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n762_), .B2(G106gat), .ZN(new_n763_));
  AOI211_X1 g562(.A(KEYINPUT52), .B(new_n466_), .C1(new_n742_), .C2(new_n267_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n760_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g565(.A(KEYINPUT115), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n545_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n767_), .B(new_n508_), .C1(new_n768_), .C2(new_n511_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n541_), .A2(new_n511_), .A3(new_n543_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n530_), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT73), .B1(new_n516_), .B2(new_n526_), .ZN(new_n773_));
  OAI22_X1  g572(.A1(new_n772_), .A2(new_n773_), .B1(new_n526_), .B2(new_n516_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n510_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n767_), .B1(new_n775_), .B2(new_n508_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n546_), .B1(new_n510_), .B2(new_n550_), .ZN(new_n777_));
  OAI22_X1  g576(.A1(new_n771_), .A2(new_n776_), .B1(new_n777_), .B2(new_n508_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n778_), .A2(new_n496_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT112), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n473_), .A2(new_n484_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n477_), .A2(KEYINPUT12), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n475_), .A2(new_n486_), .A3(new_n476_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n781_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n780_), .B1(new_n784_), .B2(KEYINPUT55), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n489_), .A2(KEYINPUT112), .A3(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT113), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(new_n489_), .B2(new_n786_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n782_), .A2(new_n783_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n791_), .A2(KEYINPUT113), .A3(KEYINPUT55), .A4(new_n485_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT66), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n473_), .B(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n484_), .B1(new_n791_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n788_), .A2(new_n793_), .A3(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(KEYINPUT56), .A3(new_n493_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT56), .B1(new_n798_), .B2(new_n493_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n799_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n796_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n494_), .B1(new_n803_), .B2(new_n793_), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n804_), .A2(KEYINPUT116), .A3(KEYINPUT56), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n779_), .B1(new_n802_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT58), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  OAI211_X1 g607(.A(KEYINPUT58), .B(new_n779_), .C1(new_n802_), .C2(new_n805_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(new_n670_), .A3(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT57), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n778_), .B1(new_n498_), .B2(new_n501_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n804_), .B2(KEYINPUT56), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n489_), .A2(KEYINPUT112), .A3(new_n786_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT112), .B1(new_n489_), .B2(new_n786_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n797_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n790_), .A2(new_n792_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n493_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT56), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(KEYINPUT114), .A3(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n814_), .A2(new_n821_), .A3(new_n799_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n554_), .A2(new_n495_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n812_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n811_), .B1(new_n825_), .B2(new_n660_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n810_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  AOI211_X1 g627(.A(new_n820_), .B(new_n494_), .C1(new_n803_), .C2(new_n793_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n819_), .A2(new_n820_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n813_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n823_), .B1(new_n831_), .B2(new_n821_), .ZN(new_n832_));
  OAI211_X1 g631(.A(KEYINPUT57), .B(new_n579_), .C1(new_n832_), .C2(new_n812_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n828_), .A2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n827_), .B1(new_n810_), .B2(new_n826_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n661_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT110), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n547_), .A2(new_n594_), .A3(new_n553_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n837_), .B(new_n838_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n612_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n837_), .B1(new_n604_), .B2(new_n838_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT54), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT111), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  OR3_X1    g643(.A1(new_n840_), .A2(new_n841_), .A3(KEYINPUT54), .ZN(new_n845_));
  OAI211_X1 g644(.A(KEYINPUT111), .B(KEYINPUT54), .C1(new_n840_), .C2(new_n841_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n844_), .A2(new_n845_), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n836_), .A2(new_n847_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n622_), .A2(new_n417_), .A3(new_n419_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n850_), .A2(KEYINPUT59), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n554_), .A2(KEYINPUT119), .A3(G113gat), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(KEYINPUT119), .B2(G113gat), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n810_), .A2(new_n833_), .A3(new_n826_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n661_), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n856_), .A2(KEYINPUT117), .A3(new_n847_), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT117), .B1(new_n856_), .B2(new_n847_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n857_), .A2(new_n858_), .A3(new_n850_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n852_), .B(new_n854_), .C1(new_n859_), .C2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n858_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n856_), .A2(new_n847_), .A3(KEYINPUT117), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n862_), .A2(new_n554_), .A3(new_n863_), .A4(new_n849_), .ZN(new_n864_));
  INV_X1    g663(.A(G113gat), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n861_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n861_), .A2(KEYINPUT120), .A3(new_n866_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1340gat));
  INV_X1    g670(.A(KEYINPUT60), .ZN(new_n872_));
  INV_X1    g671(.A(G120gat), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n505_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n874_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n859_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n876_), .B(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n852_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n879_));
  OAI21_X1  g678(.A(G120gat), .B1(new_n879_), .B2(new_n715_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n880_), .ZN(G1341gat));
  OAI21_X1  g680(.A(G127gat), .B1(new_n879_), .B2(new_n661_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n859_), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n661_), .A2(G127gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n882_), .B1(new_n883_), .B2(new_n884_), .ZN(G1342gat));
  OAI21_X1  g684(.A(G134gat), .B1(new_n879_), .B2(new_n612_), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n582_), .A2(G134gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n883_), .B2(new_n887_), .ZN(G1343gat));
  NOR3_X1   g687(.A1(new_n857_), .A2(new_n858_), .A3(new_n418_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n622_), .A2(new_n417_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n889_), .A2(new_n554_), .A3(new_n890_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g691(.A1(new_n889_), .A2(new_n605_), .A3(new_n890_), .ZN(new_n893_));
  XOR2_X1   g692(.A(KEYINPUT122), .B(G148gat), .Z(new_n894_));
  XOR2_X1   g693(.A(new_n893_), .B(new_n894_), .Z(G1345gat));
  NAND3_X1  g694(.A1(new_n889_), .A2(new_n594_), .A3(new_n890_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(KEYINPUT61), .B(G155gat), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n896_), .B(new_n897_), .ZN(G1346gat));
  NAND2_X1  g697(.A1(new_n889_), .A2(new_n890_), .ZN(new_n899_));
  OAI21_X1  g698(.A(G162gat), .B1(new_n899_), .B2(new_n612_), .ZN(new_n900_));
  OR2_X1    g699(.A1(new_n582_), .A2(G162gat), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n899_), .B2(new_n901_), .ZN(G1347gat));
  INV_X1    g701(.A(G169gat), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n597_), .A2(new_n429_), .A3(new_n324_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n268_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n905_), .B1(new_n836_), .B2(new_n847_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n903_), .B1(new_n906_), .B2(new_n554_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n908_));
  OAI21_X1  g707(.A(KEYINPUT123), .B1(new_n907_), .B2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n910_));
  AOI211_X1 g709(.A(new_n555_), .B(new_n905_), .C1(new_n836_), .C2(new_n847_), .ZN(new_n911_));
  OAI211_X1 g710(.A(new_n910_), .B(KEYINPUT62), .C1(new_n911_), .C2(new_n903_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n907_), .A2(new_n908_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n909_), .A2(new_n912_), .A3(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n911_), .A2(new_n299_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1348gat));
  AOI21_X1  g715(.A(G176gat), .B1(new_n906_), .B2(new_n505_), .ZN(new_n917_));
  NOR3_X1   g716(.A1(new_n857_), .A2(new_n858_), .A3(new_n267_), .ZN(new_n918_));
  AND3_X1   g717(.A1(new_n904_), .A2(G176gat), .A3(new_n605_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n917_), .B1(new_n918_), .B2(new_n919_), .ZN(G1349gat));
  INV_X1    g719(.A(new_n906_), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n921_), .A2(new_n290_), .A3(new_n661_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n918_), .A2(new_n594_), .A3(new_n904_), .ZN(new_n923_));
  INV_X1    g722(.A(G183gat), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n922_), .B1(new_n923_), .B2(new_n924_), .ZN(G1350gat));
  OAI21_X1  g724(.A(G190gat), .B1(new_n921_), .B2(new_n612_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n580_), .A2(new_n291_), .A3(new_n581_), .ZN(new_n927_));
  XOR2_X1   g726(.A(new_n927_), .B(KEYINPUT124), .Z(new_n928_));
  OAI21_X1  g727(.A(new_n926_), .B1(new_n921_), .B2(new_n928_), .ZN(G1351gat));
  NOR2_X1   g728(.A1(new_n597_), .A2(new_n429_), .ZN(new_n930_));
  NAND4_X1  g729(.A1(new_n889_), .A2(G197gat), .A3(new_n554_), .A4(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n418_), .ZN(new_n934_));
  NAND4_X1  g733(.A1(new_n862_), .A2(new_n934_), .A3(new_n863_), .A4(new_n930_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n935_), .A2(new_n555_), .ZN(new_n936_));
  OAI21_X1  g735(.A(KEYINPUT125), .B1(new_n936_), .B2(G197gat), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n933_), .B1(new_n937_), .B2(new_n931_), .ZN(G1352gat));
  NOR2_X1   g737(.A1(new_n935_), .A2(new_n715_), .ZN(new_n939_));
  XOR2_X1   g738(.A(new_n939_), .B(G204gat), .Z(G1353gat));
  AOI21_X1  g739(.A(new_n661_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n889_), .A2(new_n930_), .A3(new_n941_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n943_));
  XOR2_X1   g742(.A(new_n942_), .B(new_n943_), .Z(G1354gat));
  XOR2_X1   g743(.A(KEYINPUT127), .B(G218gat), .Z(new_n945_));
  NAND2_X1  g744(.A1(new_n670_), .A2(new_n945_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n935_), .A2(new_n946_), .ZN(new_n947_));
  NOR3_X1   g746(.A1(new_n935_), .A2(KEYINPUT126), .A3(new_n582_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n948_), .A2(new_n945_), .ZN(new_n949_));
  OAI21_X1  g748(.A(KEYINPUT126), .B1(new_n935_), .B2(new_n582_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n947_), .B1(new_n949_), .B2(new_n950_), .ZN(G1355gat));
endmodule


