//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 1 0 0 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n588_, new_n589_, new_n590_, new_n592_, new_n593_, new_n594_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n629_, new_n630_, new_n631_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n648_,
    new_n649_, new_n650_, new_n652_, new_n653_, new_n654_, new_n656_,
    new_n657_, new_n658_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n797_, new_n799_,
    new_n800_, new_n802_, new_n803_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n827_,
    new_n828_, new_n830_, new_n831_, new_n832_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n856_,
    new_n857_, new_n858_;
  INV_X1    g000(.A(KEYINPUT102), .ZN(new_n202_));
  XOR2_X1   g001(.A(G155gat), .B(G162gat), .Z(new_n203_));
  NAND2_X1  g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT2), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n204_), .B1(new_n205_), .B2(KEYINPUT88), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(KEYINPUT88), .ZN(new_n207_));
  MUX2_X1   g006(.A(new_n204_), .B(new_n206_), .S(new_n207_), .Z(new_n208_));
  OR2_X1    g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT3), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n203_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT1), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n203_), .A2(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n213_), .A2(new_n204_), .A3(new_n209_), .A4(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n211_), .A2(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n216_), .A2(KEYINPUT29), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G78gat), .B(G106gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  AND2_X1   g018(.A1(G228gat), .A2(G233gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G204gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(G197gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT90), .B(G197gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n223_), .B1(new_n224_), .B2(new_n222_), .ZN(new_n225_));
  XOR2_X1   g024(.A(G211gat), .B(G218gat), .Z(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(KEYINPUT21), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n225_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT91), .B(KEYINPUT21), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT92), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n229_), .A2(KEYINPUT92), .A3(new_n230_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n226_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G197gat), .A2(G204gat), .ZN(new_n236_));
  OAI211_X1 g035(.A(KEYINPUT21), .B(new_n236_), .C1(new_n224_), .C2(G204gat), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n228_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n239_), .A2(KEYINPUT93), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT93), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n216_), .A2(KEYINPUT29), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n221_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  AND3_X1   g044(.A1(new_n239_), .A2(new_n221_), .A3(new_n244_), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT89), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NOR3_X1   g047(.A1(new_n245_), .A2(KEYINPUT89), .A3(new_n246_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n219_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n249_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n219_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n251_), .A2(new_n252_), .A3(new_n247_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n250_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G22gat), .B(G50gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT28), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n254_), .A2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G8gat), .B(G36gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(G92gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT18), .B(G64gat), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n260_), .B(new_n261_), .Z(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G226gat), .A2(G233gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT19), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT26), .B(G190gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT94), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT25), .B(G183gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  OR2_X1    g069(.A1(G169gat), .A2(G176gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G169gat), .A2(G176gat), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(KEYINPUT24), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n274_), .A2(KEYINPUT95), .ZN(new_n275_));
  INV_X1    g074(.A(G183gat), .ZN(new_n276_));
  INV_X1    g075(.A(G190gat), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT23), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT23), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n279_), .A2(G183gat), .A3(G190gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  OR2_X1    g080(.A1(new_n271_), .A2(KEYINPUT24), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n274_), .A2(KEYINPUT95), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n275_), .A2(new_n281_), .A3(new_n282_), .A4(new_n283_), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n280_), .A2(KEYINPUT83), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n280_), .A2(KEYINPUT83), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n285_), .A2(new_n278_), .A3(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n287_), .B1(G183gat), .B2(G190gat), .ZN(new_n288_));
  INV_X1    g087(.A(new_n272_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT22), .B(G169gat), .ZN(new_n290_));
  INV_X1    g089(.A(G176gat), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n289_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n288_), .A2(new_n292_), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n284_), .B(new_n293_), .C1(new_n240_), .C2(new_n242_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT20), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT26), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(G190gat), .ZN(new_n297_));
  XOR2_X1   g096(.A(KEYINPUT81), .B(G190gat), .Z(new_n298_));
  OAI211_X1 g097(.A(new_n269_), .B(new_n297_), .C1(new_n298_), .C2(new_n296_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n273_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT82), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(new_n287_), .A3(new_n282_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n281_), .B1(new_n298_), .B2(G183gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n292_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n295_), .B1(new_n305_), .B2(new_n239_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n266_), .B1(new_n294_), .B2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n238_), .A2(new_n302_), .A3(new_n304_), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n293_), .B(KEYINPUT96), .Z(new_n309_));
  AND2_X1   g108(.A1(new_n284_), .A2(new_n309_), .ZN(new_n310_));
  OAI211_X1 g109(.A(KEYINPUT20), .B(new_n308_), .C1(new_n310_), .C2(new_n238_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n311_), .A2(new_n265_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n263_), .B1(new_n307_), .B2(new_n312_), .ZN(new_n313_));
  AOI211_X1 g112(.A(new_n295_), .B(new_n265_), .C1(new_n305_), .C2(new_n239_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n310_), .A2(new_n238_), .ZN(new_n315_));
  AOI22_X1  g114(.A1(new_n311_), .A2(new_n265_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n262_), .ZN(new_n317_));
  AND3_X1   g116(.A1(new_n313_), .A2(KEYINPUT27), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT27), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n311_), .A2(new_n265_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n314_), .A2(new_n315_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT97), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n322_), .A2(new_n323_), .A3(new_n263_), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT97), .B1(new_n316_), .B2(new_n262_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(new_n325_), .A3(new_n317_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n318_), .B1(new_n319_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n216_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G127gat), .B(G134gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G113gat), .B(G120gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n330_), .ZN(new_n332_));
  MUX2_X1   g131(.A(new_n331_), .B(new_n332_), .S(KEYINPUT85), .Z(new_n333_));
  NOR2_X1   g132(.A1(new_n328_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n334_), .A2(KEYINPUT4), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n328_), .A2(new_n331_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n336_), .B1(new_n333_), .B2(new_n328_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n335_), .B1(KEYINPUT4), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G225gat), .A2(G233gat), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n337_), .B1(G225gat), .B2(G233gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G1gat), .B(G29gat), .ZN(new_n342_));
  INV_X1    g141(.A(G85gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(KEYINPUT0), .B(G57gat), .Z(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  OR3_X1    g145(.A1(new_n340_), .A2(new_n341_), .A3(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n346_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n250_), .A2(new_n253_), .A3(new_n256_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n258_), .A2(new_n327_), .A3(new_n350_), .A4(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT101), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n262_), .A2(KEYINPUT32), .ZN(new_n354_));
  OR3_X1    g153(.A1(new_n322_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n354_), .B1(new_n307_), .B2(new_n312_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n353_), .B1(new_n322_), .B2(new_n354_), .ZN(new_n357_));
  AND4_X1   g156(.A1(new_n349_), .A2(new_n355_), .A3(new_n356_), .A4(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n346_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT100), .ZN(new_n360_));
  INV_X1    g159(.A(new_n338_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n360_), .B1(new_n339_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n326_), .A2(KEYINPUT98), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT98), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n324_), .A2(new_n325_), .A3(new_n364_), .A4(new_n317_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n362_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(KEYINPUT99), .A2(KEYINPUT33), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n347_), .B(new_n367_), .Z(new_n368_));
  AOI21_X1  g167(.A(new_n358_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n258_), .A2(new_n351_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n202_), .B(new_n352_), .C1(new_n369_), .C2(new_n371_), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n352_), .A2(new_n202_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n305_), .B(KEYINPUT84), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(G43gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G71gat), .B(G99gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT30), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G227gat), .A2(G233gat), .ZN(new_n378_));
  INV_X1    g177(.A(G15gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n377_), .B(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n375_), .B(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT87), .ZN(new_n383_));
  XOR2_X1   g182(.A(KEYINPUT86), .B(KEYINPUT31), .Z(new_n384_));
  XNOR2_X1  g183(.A(new_n333_), .B(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT87), .ZN(new_n387_));
  OR3_X1    g186(.A1(new_n382_), .A2(new_n387_), .A3(new_n385_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n372_), .A2(new_n373_), .A3(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n389_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n327_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n371_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n391_), .A2(new_n393_), .A3(new_n350_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n390_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G15gat), .B(G22gat), .ZN(new_n396_));
  INV_X1    g195(.A(G1gat), .ZN(new_n397_));
  INV_X1    g196(.A(G8gat), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT14), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n396_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G1gat), .B(G8gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  XOR2_X1   g201(.A(G43gat), .B(G50gat), .Z(new_n403_));
  XNOR2_X1  g202(.A(G29gat), .B(G36gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n402_), .A2(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(new_n406_), .B(KEYINPUT78), .Z(new_n407_));
  NAND2_X1  g206(.A1(new_n402_), .A2(new_n405_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT79), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G229gat), .A2(G233gat), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  XOR2_X1   g211(.A(new_n405_), .B(KEYINPUT15), .Z(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n402_), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n407_), .A2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n412_), .B1(new_n411_), .B2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G113gat), .B(G141gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G169gat), .B(G197gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n416_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT80), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n416_), .A2(new_n420_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n395_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT103), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  XOR2_X1   g226(.A(G57gat), .B(G64gat), .Z(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n429_), .A2(KEYINPUT11), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n429_), .A2(KEYINPUT11), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G71gat), .B(G78gat), .ZN(new_n432_));
  OR3_X1    g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n429_), .A2(new_n432_), .A3(KEYINPUT11), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT69), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G99gat), .A2(G106gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT6), .ZN(new_n439_));
  INV_X1    g238(.A(G99gat), .ZN(new_n440_));
  INV_X1    g239(.A(G106gat), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT65), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n440_), .B(new_n441_), .C1(new_n442_), .C2(KEYINPUT7), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT7), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n444_), .B(KEYINPUT65), .C1(G99gat), .C2(G106gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n439_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT8), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G85gat), .B(G92gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n447_), .A2(new_n448_), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT67), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n446_), .A2(KEYINPUT66), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT66), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n443_), .A2(new_n445_), .A3(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n453_), .A2(new_n439_), .A3(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n450_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n452_), .B1(new_n457_), .B2(KEYINPUT8), .ZN(new_n458_));
  AOI211_X1 g257(.A(KEYINPUT67), .B(new_n448_), .C1(new_n456_), .C2(new_n450_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n451_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT68), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT68), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n462_), .B(new_n451_), .C1(new_n458_), .C2(new_n459_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n449_), .A2(KEYINPUT9), .ZN(new_n465_));
  INV_X1    g264(.A(G92gat), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n343_), .A2(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n465_), .B1(KEYINPUT9), .B2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT64), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT10), .B(G99gat), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n441_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n469_), .A2(new_n472_), .A3(new_n439_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n437_), .B1(new_n464_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n473_), .ZN(new_n475_));
  AOI211_X1 g274(.A(KEYINPUT69), .B(new_n475_), .C1(new_n461_), .C2(new_n463_), .ZN(new_n476_));
  OAI211_X1 g275(.A(KEYINPUT12), .B(new_n436_), .C1(new_n474_), .C2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n460_), .A2(new_n473_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n436_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n480_), .A2(KEYINPUT12), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT70), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n460_), .A2(new_n435_), .A3(new_n473_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(G230gat), .ZN(new_n485_));
  INV_X1    g284(.A(G233gat), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n482_), .B1(new_n484_), .B2(new_n487_), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n483_), .B(KEYINPUT70), .C1(new_n485_), .C2(new_n486_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n477_), .A2(new_n481_), .A3(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n487_), .B1(new_n480_), .B2(new_n484_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G176gat), .B(G204gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G120gat), .B(G148gat), .ZN(new_n496_));
  XOR2_X1   g295(.A(new_n495_), .B(new_n496_), .Z(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n491_), .A2(new_n492_), .A3(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT72), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n491_), .A2(new_n492_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n500_), .B1(new_n501_), .B2(new_n498_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT13), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n478_), .A2(new_n405_), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n443_), .A2(new_n445_), .A3(new_n454_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n454_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n449_), .B1(new_n507_), .B2(new_n439_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT67), .B1(new_n508_), .B2(new_n448_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n457_), .A2(new_n452_), .A3(KEYINPUT8), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n462_), .B1(new_n511_), .B2(new_n451_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n463_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n473_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT69), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n464_), .A2(new_n437_), .A3(new_n473_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n504_), .B1(new_n517_), .B2(new_n413_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G232gat), .A2(G233gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT34), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT35), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(KEYINPUT73), .B1(new_n517_), .B2(new_n413_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n521_), .A2(new_n522_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n518_), .B(new_n523_), .C1(new_n524_), .C2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G134gat), .B(G162gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(G218gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT74), .B(G190gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n531_), .A2(KEYINPUT36), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n413_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n533_), .B1(new_n405_), .B2(new_n478_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT73), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n534_), .A2(new_n536_), .A3(new_n525_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n527_), .A2(new_n532_), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT75), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n527_), .A2(KEYINPUT75), .A3(new_n537_), .A4(new_n532_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n532_), .B1(new_n527_), .B2(new_n537_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n531_), .A2(KEYINPUT36), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(KEYINPUT76), .A2(KEYINPUT37), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(KEYINPUT76), .A2(KEYINPUT37), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n546_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n540_), .A2(new_n541_), .B1(new_n544_), .B2(new_n543_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n551_), .A2(KEYINPUT76), .A3(KEYINPUT37), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  XOR2_X1   g352(.A(new_n435_), .B(new_n402_), .Z(new_n554_));
  NAND2_X1  g353(.A1(G231gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G183gat), .B(G211gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G127gat), .B(G155gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n559_), .B(new_n560_), .Z(new_n561_));
  XOR2_X1   g360(.A(new_n561_), .B(KEYINPUT17), .Z(new_n562_));
  OR2_X1    g361(.A1(new_n556_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n561_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n556_), .A2(KEYINPUT17), .A3(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n553_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n395_), .A2(KEYINPUT103), .A3(new_n424_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n427_), .A2(new_n503_), .A3(new_n567_), .A4(new_n568_), .ZN(new_n569_));
  NOR3_X1   g368(.A1(new_n569_), .A2(G1gat), .A3(new_n350_), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n570_), .A2(KEYINPUT38), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n551_), .B1(new_n390_), .B2(new_n394_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n566_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n503_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n424_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  AND3_X1   g375(.A1(new_n572_), .A2(new_n573_), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(G1gat), .B1(new_n578_), .B2(new_n350_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n570_), .A2(KEYINPUT38), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n571_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n581_), .B(KEYINPUT104), .Z(G1324gat));
  AOI21_X1  g381(.A(new_n398_), .B1(new_n577_), .B2(new_n392_), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n583_), .B(KEYINPUT39), .Z(new_n584_));
  NAND2_X1  g383(.A1(new_n392_), .A2(new_n398_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n584_), .B1(new_n569_), .B2(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n586_), .B(KEYINPUT40), .Z(G1325gat));
  AOI21_X1  g386(.A(new_n379_), .B1(new_n577_), .B2(new_n391_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT41), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n391_), .A2(new_n379_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n589_), .B1(new_n569_), .B2(new_n590_), .ZN(G1326gat));
  OAI21_X1  g390(.A(G22gat), .B1(new_n578_), .B2(new_n370_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT42), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n370_), .A2(G22gat), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n593_), .B1(new_n569_), .B2(new_n594_), .ZN(G1327gat));
  NOR2_X1   g394(.A1(new_n546_), .A2(new_n573_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n427_), .A2(new_n503_), .A3(new_n568_), .A4(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(G29gat), .B1(new_n598_), .B2(new_n349_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n395_), .A2(new_n553_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT43), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT43), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n395_), .A2(new_n602_), .A3(new_n553_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n604_), .A2(new_n566_), .A3(new_n576_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT44), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  AND3_X1   g406(.A1(new_n607_), .A2(G29gat), .A3(new_n349_), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n605_), .A2(new_n606_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n599_), .B1(new_n608_), .B2(new_n609_), .ZN(G1328gat));
  NAND3_X1  g409(.A1(new_n609_), .A2(new_n392_), .A3(new_n607_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(G36gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n327_), .B(KEYINPUT105), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n597_), .A2(G36gat), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT106), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NOR4_X1   g416(.A1(new_n597_), .A2(KEYINPUT106), .A3(G36gat), .A4(new_n614_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n617_), .A2(KEYINPUT45), .A3(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT45), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n615_), .A2(new_n616_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n621_), .B1(new_n622_), .B2(new_n618_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n612_), .A2(new_n620_), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT46), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n612_), .A2(new_n620_), .A3(new_n623_), .A4(KEYINPUT46), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(G1329gat));
  NAND4_X1  g427(.A1(new_n609_), .A2(G43gat), .A3(new_n391_), .A4(new_n607_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n597_), .A2(new_n389_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n629_), .B1(G43gat), .B2(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g431(.A1(new_n597_), .A2(G50gat), .A3(new_n370_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n609_), .A2(new_n371_), .A3(new_n607_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT107), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n634_), .A2(new_n635_), .A3(G50gat), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n635_), .B1(new_n634_), .B2(G50gat), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n633_), .B1(new_n636_), .B2(new_n637_), .ZN(G1331gat));
  NOR2_X1   g437(.A1(new_n503_), .A2(new_n424_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n572_), .A2(new_n573_), .A3(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G57gat), .B1(new_n640_), .B2(new_n350_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n639_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n642_), .B1(new_n390_), .B2(new_n394_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(new_n567_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n350_), .A2(G57gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n641_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n646_), .B(KEYINPUT108), .Z(G1332gat));
  OAI21_X1  g446(.A(G64gat), .B1(new_n640_), .B2(new_n614_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT48), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n614_), .A2(G64gat), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n649_), .B1(new_n644_), .B2(new_n650_), .ZN(G1333gat));
  OAI21_X1  g450(.A(G71gat), .B1(new_n640_), .B2(new_n389_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT49), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n389_), .A2(G71gat), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n653_), .B1(new_n644_), .B2(new_n654_), .ZN(G1334gat));
  OAI21_X1  g454(.A(G78gat), .B1(new_n640_), .B2(new_n370_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT50), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n370_), .A2(G78gat), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n657_), .B1(new_n644_), .B2(new_n658_), .ZN(G1335gat));
  INV_X1    g458(.A(new_n553_), .ZN(new_n660_));
  AOI211_X1 g459(.A(KEYINPUT43), .B(new_n660_), .C1(new_n390_), .C2(new_n394_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n602_), .B1(new_n395_), .B2(new_n553_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n566_), .B(new_n639_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n663_), .A2(new_n343_), .A3(new_n350_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n643_), .A2(new_n596_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(G85gat), .B1(new_n666_), .B2(new_n349_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n664_), .A2(new_n667_), .ZN(G1336gat));
  NOR3_X1   g467(.A1(new_n663_), .A2(new_n466_), .A3(new_n614_), .ZN(new_n669_));
  AOI21_X1  g468(.A(G92gat), .B1(new_n666_), .B2(new_n392_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1337gat));
  OAI21_X1  g470(.A(G99gat), .B1(new_n663_), .B2(new_n389_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n666_), .A2(new_n391_), .A3(new_n471_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT51), .ZN(G1338gat));
  NOR3_X1   g474(.A1(new_n665_), .A2(G106gat), .A3(new_n370_), .ZN(new_n676_));
  OAI21_X1  g475(.A(KEYINPUT109), .B1(new_n663_), .B2(new_n370_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n642_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT109), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n678_), .A2(new_n679_), .A3(new_n566_), .A4(new_n371_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n677_), .A2(new_n680_), .A3(G106gat), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT52), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT52), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n677_), .A2(new_n680_), .A3(new_n683_), .A4(G106gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n676_), .B1(new_n682_), .B2(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n685_), .B(new_n687_), .ZN(G1339gat));
  NAND2_X1  g487(.A1(new_n391_), .A2(new_n393_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n549_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n551_), .A2(new_n547_), .A3(new_n690_), .ZN(new_n691_));
  AND4_X1   g490(.A1(KEYINPUT76), .A2(new_n542_), .A3(KEYINPUT37), .A4(new_n545_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n411_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n420_), .B1(new_n415_), .B2(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n694_), .B1(new_n693_), .B2(new_n410_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT114), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n696_), .A2(new_n421_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n500_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT56), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n477_), .A2(new_n483_), .A3(new_n481_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n487_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n477_), .A2(KEYINPUT55), .A3(new_n481_), .A4(new_n490_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT55), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n491_), .A2(KEYINPUT112), .A3(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(KEYINPUT112), .B1(new_n491_), .B2(new_n704_), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n703_), .A2(new_n705_), .A3(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n699_), .B1(new_n707_), .B2(new_n498_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n477_), .A2(new_n481_), .A3(new_n490_), .ZN(new_n709_));
  AOI22_X1  g508(.A1(new_n709_), .A2(KEYINPUT55), .B1(new_n700_), .B2(new_n487_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT112), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n711_), .B1(new_n709_), .B2(KEYINPUT55), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n491_), .A2(KEYINPUT112), .A3(new_n704_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n710_), .A2(new_n712_), .A3(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n714_), .A2(KEYINPUT56), .A3(new_n497_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n698_), .B1(new_n708_), .B2(new_n715_), .ZN(new_n716_));
  OAI22_X1  g515(.A1(new_n691_), .A2(new_n692_), .B1(new_n716_), .B2(KEYINPUT58), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT116), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(KEYINPUT58), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT58), .ZN(new_n720_));
  INV_X1    g519(.A(new_n715_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT56), .B1(new_n714_), .B2(new_n497_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n720_), .B1(new_n723_), .B2(new_n698_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT116), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n724_), .A2(new_n553_), .A3(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n718_), .A2(new_n719_), .A3(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n708_), .A2(KEYINPUT113), .A3(new_n715_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT113), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n714_), .A2(new_n729_), .A3(KEYINPUT56), .A4(new_n497_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n730_), .A2(new_n500_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n728_), .A2(new_n731_), .A3(new_n424_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n502_), .A2(new_n697_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n551_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(KEYINPUT115), .B1(new_n734_), .B2(KEYINPUT57), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(KEYINPUT57), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT115), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT57), .ZN(new_n738_));
  INV_X1    g537(.A(new_n733_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n714_), .A2(new_n497_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n729_), .B1(new_n740_), .B2(new_n699_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n575_), .B1(new_n741_), .B2(new_n715_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n739_), .B1(new_n742_), .B2(new_n731_), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n737_), .B(new_n738_), .C1(new_n743_), .C2(new_n551_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n727_), .A2(new_n735_), .A3(new_n736_), .A4(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n566_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT54), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n567_), .A2(new_n747_), .A3(new_n575_), .A4(new_n503_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT111), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NOR3_X1   g549(.A1(new_n553_), .A2(new_n566_), .A3(new_n424_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(new_n503_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT54), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n751_), .A2(KEYINPUT111), .A3(new_n747_), .A4(new_n503_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n750_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n755_));
  AOI211_X1 g554(.A(new_n350_), .B(new_n689_), .C1(new_n746_), .C2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(G113gat), .B1(new_n756_), .B2(new_n424_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n746_), .A2(new_n755_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n689_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n758_), .A2(new_n349_), .A3(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n738_), .B1(new_n743_), .B2(new_n551_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n727_), .A2(new_n736_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n566_), .ZN(new_n763_));
  AOI211_X1 g562(.A(KEYINPUT59), .B(new_n689_), .C1(new_n763_), .C2(new_n755_), .ZN(new_n764_));
  AOI22_X1  g563(.A1(KEYINPUT59), .A2(new_n760_), .B1(new_n764_), .B2(new_n349_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n765_), .B1(KEYINPUT117), .B2(G113gat), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(G113gat), .B1(new_n575_), .B2(KEYINPUT117), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n757_), .B1(new_n767_), .B2(new_n768_), .ZN(G1340gat));
  INV_X1    g568(.A(G120gat), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n770_), .B1(new_n503_), .B2(KEYINPUT60), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n756_), .B(new_n771_), .C1(KEYINPUT60), .C2(new_n770_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT118), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n765_), .A2(new_n574_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n773_), .B1(new_n775_), .B2(new_n770_), .ZN(G1341gat));
  INV_X1    g575(.A(G127gat), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n777_), .B1(new_n765_), .B2(new_n573_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n760_), .A2(G127gat), .A3(new_n566_), .ZN(new_n779_));
  OAI21_X1  g578(.A(KEYINPUT119), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n763_), .A2(new_n755_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT59), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n781_), .A2(new_n782_), .A3(new_n349_), .A4(new_n759_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n756_), .B2(new_n782_), .ZN(new_n784_));
  OAI21_X1  g583(.A(G127gat), .B1(new_n784_), .B2(new_n566_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT119), .ZN(new_n786_));
  INV_X1    g585(.A(new_n779_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n785_), .A2(new_n786_), .A3(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n780_), .A2(new_n788_), .ZN(G1342gat));
  AOI21_X1  g588(.A(G134gat), .B1(new_n756_), .B2(new_n551_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n553_), .A2(G134gat), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n765_), .B2(new_n791_), .ZN(G1343gat));
  NOR2_X1   g591(.A1(new_n391_), .A2(new_n370_), .ZN(new_n793_));
  AND4_X1   g592(.A1(new_n349_), .A2(new_n758_), .A3(new_n614_), .A4(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n424_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n574_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g597(.A1(new_n794_), .A2(new_n573_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(KEYINPUT61), .B(G155gat), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n799_), .B(new_n800_), .ZN(G1346gat));
  AOI21_X1  g600(.A(G162gat), .B1(new_n794_), .B2(new_n551_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n553_), .A2(G162gat), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n794_), .B2(new_n803_), .ZN(G1347gat));
  INV_X1    g603(.A(KEYINPUT120), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n614_), .A2(new_n349_), .A3(new_n389_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n806_), .A2(new_n370_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n781_), .A2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n805_), .B1(new_n808_), .B2(new_n575_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n781_), .A2(KEYINPUT120), .A3(new_n424_), .A4(new_n807_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(G169gat), .A3(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT121), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT121), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n809_), .A2(new_n813_), .A3(G169gat), .A4(new_n810_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n812_), .A2(KEYINPUT62), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n808_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n816_), .A2(new_n290_), .A3(new_n424_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT62), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n811_), .A2(KEYINPUT121), .A3(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n815_), .A2(new_n817_), .A3(new_n819_), .ZN(G1348gat));
  AOI21_X1  g619(.A(G176gat), .B1(new_n816_), .B2(new_n574_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n371_), .B1(new_n746_), .B2(new_n755_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(KEYINPUT122), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n823_), .A2(new_n806_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n503_), .A2(new_n291_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n821_), .B1(new_n824_), .B2(new_n825_), .ZN(G1349gat));
  NOR3_X1   g625(.A1(new_n808_), .A2(new_n566_), .A3(new_n269_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n823_), .A2(new_n573_), .A3(new_n806_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n827_), .B1(new_n828_), .B2(new_n276_), .ZN(G1350gat));
  OAI21_X1  g628(.A(G190gat), .B1(new_n808_), .B2(new_n660_), .ZN(new_n830_));
  XOR2_X1   g629(.A(new_n830_), .B(KEYINPUT123), .Z(new_n831_));
  NAND3_X1  g630(.A1(new_n816_), .A2(new_n268_), .A3(new_n551_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(G1351gat));
  NAND2_X1  g632(.A1(new_n793_), .A2(new_n350_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n834_), .A2(KEYINPUT124), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n835_), .A2(new_n614_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(KEYINPUT124), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n758_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT125), .ZN(new_n839_));
  AOI22_X1  g638(.A1(new_n746_), .A2(new_n755_), .B1(KEYINPUT124), .B2(new_n834_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT125), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n841_), .A3(new_n836_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n839_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n424_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n574_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n222_), .A2(KEYINPUT126), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(G1353gat));
  NOR2_X1   g647(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(KEYINPUT127), .ZN(new_n850_));
  NAND2_X1  g649(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n851_));
  AND4_X1   g650(.A1(new_n573_), .A2(new_n843_), .A3(new_n850_), .A4(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n566_), .B1(new_n839_), .B2(new_n842_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n850_), .B1(new_n853_), .B2(new_n851_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n852_), .A2(new_n854_), .ZN(G1354gat));
  NAND3_X1  g654(.A1(new_n843_), .A2(G218gat), .A3(new_n553_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n546_), .B1(new_n839_), .B2(new_n842_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(G218gat), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(G1355gat));
endmodule


