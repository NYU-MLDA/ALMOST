//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 1 1 0 0 0 0 0 1 0 1 0 1 0 0 1 0 1 1 1 1 1 1 0 0 0 0 0 1 1 1 1 0 1 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n927_, new_n929_, new_n930_,
    new_n931_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_,
    new_n959_, new_n960_;
  XOR2_X1   g000(.A(G29gat), .B(G36gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G29gat), .B(G36gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G43gat), .B(G50gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT78), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G15gat), .B(G22gat), .ZN(new_n211_));
  INV_X1    g010(.A(G1gat), .ZN(new_n212_));
  INV_X1    g011(.A(G8gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT14), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G1gat), .B(G8gat), .ZN(new_n216_));
  XOR2_X1   g015(.A(new_n215_), .B(new_n216_), .Z(new_n217_));
  NAND2_X1  g016(.A1(new_n210_), .A2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n208_), .B(KEYINPUT15), .ZN(new_n219_));
  INV_X1    g018(.A(new_n217_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n218_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G229gat), .A2(G233gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n224_), .A2(KEYINPUT79), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(KEYINPUT79), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n210_), .B(new_n217_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n223_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n225_), .A2(new_n226_), .A3(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT80), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G113gat), .B(G141gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G169gat), .B(G197gat), .ZN(new_n234_));
  XOR2_X1   g033(.A(new_n233_), .B(new_n234_), .Z(new_n235_));
  XNOR2_X1  g034(.A(new_n232_), .B(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G78gat), .B(G106gat), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n240_));
  INV_X1    g039(.A(G141gat), .ZN(new_n241_));
  INV_X1    g040(.A(G148gat), .ZN(new_n242_));
  AND4_X1   g041(.A1(KEYINPUT90), .A2(new_n240_), .A3(new_n241_), .A4(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(G141gat), .A2(G148gat), .ZN(new_n244_));
  AOI21_X1  g043(.A(KEYINPUT90), .B1(new_n244_), .B2(new_n240_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G141gat), .A2(G148gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT2), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT2), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(G141gat), .A3(G148gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n241_), .A2(new_n242_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT3), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT91), .B1(new_n246_), .B2(new_n254_), .ZN(new_n255_));
  AOI22_X1  g054(.A1(new_n248_), .A2(new_n250_), .B1(new_n252_), .B2(KEYINPUT3), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT91), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n256_), .B(new_n257_), .C1(new_n245_), .C2(new_n243_), .ZN(new_n258_));
  AND2_X1   g057(.A1(G155gat), .A2(G162gat), .ZN(new_n259_));
  NOR2_X1   g058(.A1(G155gat), .A2(G162gat), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n255_), .A2(new_n258_), .A3(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n244_), .B(KEYINPUT89), .ZN(new_n263_));
  AOI22_X1  g062(.A1(new_n259_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n264_));
  INV_X1    g063(.A(new_n261_), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n263_), .B(new_n264_), .C1(KEYINPUT1), .C2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n262_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT92), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT92), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n262_), .A2(new_n269_), .A3(new_n266_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n268_), .A2(KEYINPUT29), .A3(new_n270_), .ZN(new_n271_));
  XOR2_X1   g070(.A(G197gat), .B(G204gat), .Z(new_n272_));
  NOR2_X1   g071(.A1(new_n272_), .A2(KEYINPUT21), .ZN(new_n273_));
  XOR2_X1   g072(.A(G211gat), .B(G218gat), .Z(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(G197gat), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n276_), .A2(KEYINPUT94), .A3(G204gat), .ZN(new_n277_));
  OAI211_X1 g076(.A(KEYINPUT21), .B(new_n277_), .C1(new_n272_), .C2(KEYINPUT94), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n275_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n272_), .A2(new_n274_), .A3(KEYINPUT21), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G228gat), .A2(G233gat), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n271_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT95), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT95), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n271_), .A2(new_n286_), .A3(new_n283_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n267_), .A2(KEYINPUT29), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n282_), .B1(new_n289_), .B2(new_n281_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n239_), .B1(new_n288_), .B2(new_n291_), .ZN(new_n292_));
  AOI211_X1 g091(.A(new_n238_), .B(new_n290_), .C1(new_n285_), .C2(new_n287_), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT97), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n268_), .A2(new_n270_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT29), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT93), .B(KEYINPUT28), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(G22gat), .B(G50gat), .Z(new_n301_));
  INV_X1    g100(.A(new_n270_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n269_), .B1(new_n262_), .B2(new_n266_), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n296_), .B(new_n298_), .C1(new_n302_), .C2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n300_), .A2(new_n301_), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n301_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n304_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n298_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n306_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n305_), .A2(new_n309_), .ZN(new_n310_));
  AND3_X1   g109(.A1(new_n271_), .A2(new_n286_), .A3(new_n283_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n286_), .B1(new_n271_), .B2(new_n283_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n291_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n238_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n310_), .B1(new_n314_), .B2(KEYINPUT96), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n288_), .A2(new_n291_), .A3(new_n239_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT97), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n314_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n294_), .A2(new_n315_), .A3(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n315_), .B1(new_n294_), .B2(new_n318_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G127gat), .B(G134gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G113gat), .B(G120gat), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n324_), .A2(KEYINPUT87), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n322_), .B(new_n323_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n325_), .B1(new_n326_), .B2(KEYINPUT87), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n268_), .A2(new_n327_), .A3(new_n270_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n262_), .A2(new_n326_), .A3(new_n266_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G225gat), .A2(G233gat), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n328_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  AND3_X1   g130(.A1(new_n328_), .A2(KEYINPUT4), .A3(new_n329_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT4), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n268_), .A2(new_n333_), .A3(new_n327_), .A4(new_n270_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n330_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n331_), .B1(new_n332_), .B2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G1gat), .B(G29gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(G85gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT0), .B(G57gat), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n339_), .B(new_n340_), .Z(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n337_), .A2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n328_), .A2(KEYINPUT4), .A3(new_n329_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n344_), .A2(new_n335_), .A3(new_n334_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n345_), .A2(new_n331_), .A3(new_n341_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n343_), .A2(new_n346_), .ZN(new_n347_));
  XOR2_X1   g146(.A(G8gat), .B(G36gat), .Z(new_n348_));
  XNOR2_X1  g147(.A(G64gat), .B(G92gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT32), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT104), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G183gat), .A2(G190gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT23), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT23), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n358_), .A2(G183gat), .A3(G190gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(G190gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT81), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT81), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(G190gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n360_), .B1(new_n365_), .B2(G183gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G169gat), .A2(G176gat), .ZN(new_n367_));
  INV_X1    g166(.A(G176gat), .ZN(new_n368_));
  INV_X1    g167(.A(G169gat), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT22), .B1(new_n369_), .B2(KEYINPUT84), .ZN(new_n370_));
  OR2_X1    g169(.A1(new_n369_), .A2(KEYINPUT22), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n368_), .B(new_n370_), .C1(new_n371_), .C2(KEYINPUT84), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n366_), .A2(new_n367_), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT82), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT25), .B(G183gat), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT26), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n376_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n374_), .B(new_n375_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT24), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n380_), .A2(new_n369_), .A3(new_n368_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n367_), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n381_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT83), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n356_), .A2(new_n386_), .A3(KEYINPUT23), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n386_), .B1(new_n356_), .B2(KEYINPUT23), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n359_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n379_), .A2(new_n385_), .A3(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n378_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT81), .B(G190gat), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n392_), .B1(new_n393_), .B2(new_n376_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n374_), .B1(new_n394_), .B2(new_n375_), .ZN(new_n395_));
  OAI211_X1 g194(.A(KEYINPUT85), .B(new_n373_), .C1(new_n391_), .C2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n378_), .B1(new_n365_), .B2(KEYINPUT26), .ZN(new_n398_));
  INV_X1    g197(.A(new_n375_), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT82), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n357_), .A2(KEYINPUT83), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n387_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n384_), .B1(new_n402_), .B2(new_n359_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n400_), .A2(new_n379_), .A3(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(KEYINPUT85), .B1(new_n404_), .B2(new_n373_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n281_), .B1(new_n397_), .B2(new_n405_), .ZN(new_n406_));
  OR2_X1    g205(.A1(G183gat), .A2(G190gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n390_), .A2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT22), .B(G169gat), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n382_), .B1(new_n409_), .B2(new_n368_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT26), .B(G190gat), .ZN(new_n412_));
  AOI22_X1  g211(.A1(new_n375_), .A2(new_n412_), .B1(new_n359_), .B2(new_n357_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n385_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n411_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT103), .ZN(new_n416_));
  INV_X1    g215(.A(new_n281_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT103), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n411_), .A2(new_n418_), .A3(new_n414_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n416_), .A2(new_n417_), .A3(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n406_), .A2(KEYINPUT20), .A3(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G226gat), .A2(G233gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT19), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n421_), .A2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n373_), .B1(new_n391_), .B2(new_n395_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT85), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(new_n396_), .A3(new_n417_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n423_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT20), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n430_), .B1(new_n281_), .B2(new_n415_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n428_), .A2(new_n429_), .A3(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n355_), .B1(new_n424_), .B2(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT104), .B1(new_n421_), .B2(new_n423_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n354_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n428_), .A2(new_n431_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n423_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT98), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n436_), .A2(KEYINPUT98), .A3(new_n423_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n415_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n423_), .B1(new_n417_), .B2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n406_), .A2(KEYINPUT20), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT99), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n427_), .A2(new_n396_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n430_), .B1(new_n447_), .B2(new_n281_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n448_), .A2(KEYINPUT99), .A3(new_n443_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n446_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n441_), .A2(new_n450_), .A3(new_n353_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n347_), .A2(new_n435_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT105), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n334_), .A2(new_n330_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n341_), .B1(new_n455_), .B2(new_n344_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n328_), .A2(new_n329_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT102), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT102), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n328_), .A2(new_n459_), .A3(new_n329_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(new_n335_), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n456_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT101), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT33), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n345_), .A2(new_n331_), .A3(new_n341_), .A4(new_n465_), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n462_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n441_), .A2(new_n352_), .A3(new_n450_), .ZN(new_n468_));
  AOI21_X1  g267(.A(KEYINPUT99), .B1(new_n448_), .B2(new_n443_), .ZN(new_n469_));
  AND4_X1   g268(.A1(KEYINPUT99), .A2(new_n406_), .A3(KEYINPUT20), .A4(new_n443_), .ZN(new_n470_));
  AOI21_X1  g269(.A(KEYINPUT98), .B1(new_n436_), .B2(new_n423_), .ZN(new_n471_));
  AOI211_X1 g270(.A(new_n438_), .B(new_n429_), .C1(new_n428_), .C2(new_n431_), .ZN(new_n472_));
  OAI22_X1  g271(.A1(new_n469_), .A2(new_n470_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n352_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n346_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n467_), .A2(new_n468_), .A3(new_n475_), .A4(new_n476_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n347_), .A2(new_n435_), .A3(KEYINPUT105), .A4(new_n451_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n454_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n321_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n475_), .A2(new_n468_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT27), .ZN(new_n482_));
  AOI22_X1  g281(.A1(new_n439_), .A2(new_n440_), .B1(new_n446_), .B2(new_n449_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n482_), .B1(new_n483_), .B2(new_n352_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n474_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n485_));
  AOI22_X1  g284(.A1(new_n481_), .A2(new_n482_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n347_), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n486_), .B(new_n487_), .C1(new_n319_), .C2(new_n320_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G15gat), .B(G43gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT86), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT30), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n447_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(G99gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n427_), .A2(KEYINPUT30), .A3(new_n396_), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n493_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n494_), .B1(new_n493_), .B2(new_n495_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n491_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n493_), .A2(new_n495_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(G99gat), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n493_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(new_n490_), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G227gat), .A2(G233gat), .ZN(new_n503_));
  INV_X1    g302(.A(G71gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n498_), .A2(new_n502_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT88), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n505_), .B1(new_n498_), .B2(new_n502_), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT31), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n498_), .A2(new_n502_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n505_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT31), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n513_), .A2(new_n507_), .A3(new_n514_), .A4(new_n506_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n510_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n327_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n510_), .A2(new_n327_), .A3(new_n515_), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n480_), .A2(new_n488_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n510_), .A2(new_n327_), .A3(new_n515_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n327_), .B1(new_n510_), .B2(new_n515_), .ZN(new_n522_));
  NOR3_X1   g321(.A1(new_n521_), .A2(new_n522_), .A3(new_n347_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n294_), .A2(new_n318_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n315_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n294_), .A2(new_n315_), .A3(new_n318_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n473_), .A2(new_n474_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n352_), .B1(new_n441_), .B2(new_n450_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n482_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n485_), .A2(KEYINPUT27), .A3(new_n468_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n528_), .A2(new_n533_), .ZN(new_n534_));
  AOI22_X1  g333(.A1(new_n520_), .A2(KEYINPUT106), .B1(new_n523_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT106), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n533_), .B1(new_n527_), .B2(new_n526_), .ZN(new_n537_));
  AOI22_X1  g336(.A1(new_n537_), .A2(new_n487_), .B1(new_n321_), .B2(new_n479_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n521_), .A2(new_n522_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n536_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n237_), .B1(new_n535_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G232gat), .A2(G233gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT34), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT35), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT71), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G85gat), .A2(G92gat), .ZN(new_n547_));
  INV_X1    g346(.A(G85gat), .ZN(new_n548_));
  INV_X1    g347(.A(G92gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(G99gat), .A2(G106gat), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT7), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G99gat), .A2(G106gat), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT6), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n547_), .B(new_n550_), .C1(new_n553_), .C2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT8), .ZN(new_n558_));
  INV_X1    g357(.A(new_n556_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT9), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT65), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n547_), .A2(new_n561_), .A3(new_n560_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n561_), .B1(new_n547_), .B2(new_n560_), .ZN(new_n563_));
  OAI221_X1 g362(.A(new_n550_), .B1(new_n560_), .B2(new_n547_), .C1(new_n562_), .C2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(KEYINPUT10), .B(G99gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT64), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n559_), .B(new_n564_), .C1(new_n566_), .C2(G106gat), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n558_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(new_n208_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n543_), .A2(KEYINPUT35), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT72), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n572_), .A2(KEYINPUT73), .ZN(new_n573_));
  INV_X1    g372(.A(new_n568_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(new_n219_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n575_), .B1(new_n572_), .B2(KEYINPUT73), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n546_), .B1(new_n573_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT74), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G190gat), .B(G218gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT75), .ZN(new_n581_));
  XOR2_X1   g380(.A(G134gat), .B(G162gat), .Z(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n584_), .A2(KEYINPUT36), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n575_), .A2(new_n545_), .A3(new_n569_), .A4(new_n571_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n579_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT77), .B(KEYINPUT37), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n579_), .A2(new_n586_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n583_), .B(KEYINPUT36), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n587_), .B(new_n588_), .C1(new_n589_), .C2(new_n591_), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n579_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n590_), .B(KEYINPUT76), .Z(new_n594_));
  AOI21_X1  g393(.A(new_n594_), .B1(new_n579_), .B2(new_n586_), .ZN(new_n595_));
  OAI21_X1  g394(.A(KEYINPUT37), .B1(new_n593_), .B2(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n592_), .A2(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(KEYINPUT66), .B(G71gat), .Z(new_n598_));
  INV_X1    g397(.A(G78gat), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT66), .B(G71gat), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(G78gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G57gat), .B(G64gat), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n600_), .B(new_n602_), .C1(KEYINPUT11), .C2(new_n603_), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n604_), .A2(KEYINPUT67), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(KEYINPUT67), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n603_), .A2(KEYINPUT11), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n605_), .A2(new_n606_), .A3(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n608_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(new_n574_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(new_n574_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT12), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n613_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G230gat), .A2(G233gat), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n611_), .A2(KEYINPUT68), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n611_), .A2(KEYINPUT68), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n618_), .A2(KEYINPUT12), .A3(new_n574_), .A4(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n616_), .A2(new_n617_), .A3(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n611_), .A2(new_n568_), .ZN(new_n622_));
  OAI211_X1 g421(.A(G230gat), .B(G233gat), .C1(new_n614_), .C2(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(KEYINPUT69), .B(KEYINPUT5), .Z(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT70), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G120gat), .B(G148gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G176gat), .B(G204gat), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n627_), .B(new_n628_), .Z(new_n629_));
  AND3_X1   g428(.A1(new_n621_), .A2(new_n623_), .A3(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n621_), .B2(new_n623_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n632_), .A2(KEYINPUT13), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(KEYINPUT13), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT17), .ZN(new_n636_));
  XOR2_X1   g435(.A(G127gat), .B(G155gat), .Z(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT16), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G183gat), .B(G211gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n618_), .A2(new_n619_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(G231gat), .A2(G233gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n217_), .B(new_n642_), .ZN(new_n643_));
  AOI211_X1 g442(.A(new_n636_), .B(new_n640_), .C1(new_n641_), .C2(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n644_), .B1(new_n641_), .B2(new_n643_), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n611_), .A2(new_n643_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n611_), .A2(new_n643_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n640_), .B(KEYINPUT17), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n646_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n645_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n597_), .A2(new_n635_), .A3(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n541_), .A2(new_n652_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n653_), .A2(G1gat), .A3(new_n487_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT107), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n655_), .A2(KEYINPUT38), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(KEYINPUT38), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n539_), .A2(new_n487_), .A3(new_n534_), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n454_), .A2(new_n478_), .A3(new_n477_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n488_), .B1(new_n659_), .B2(new_n528_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n518_), .A2(new_n519_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n660_), .A2(KEYINPUT106), .A3(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n540_), .A2(new_n658_), .A3(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n587_), .B1(new_n589_), .B2(new_n591_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT108), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n663_), .A2(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n667_), .A2(KEYINPUT109), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT109), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n669_), .B1(new_n663_), .B2(new_n666_), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n635_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(new_n236_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n673_), .A2(new_n651_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n671_), .A2(new_n347_), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(G1gat), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n656_), .A2(new_n657_), .A3(new_n676_), .ZN(G1324gat));
  NAND4_X1  g476(.A1(new_n541_), .A2(new_n213_), .A3(new_n533_), .A4(new_n652_), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n533_), .B(new_n674_), .C1(new_n668_), .C2(new_n670_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT39), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n679_), .A2(new_n680_), .A3(G8gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n679_), .B2(G8gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n678_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT40), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  OAI211_X1 g484(.A(KEYINPUT40), .B(new_n678_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1325gat));
  OAI211_X1 g486(.A(new_n539_), .B(new_n674_), .C1(new_n668_), .C2(new_n670_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT110), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n688_), .A2(new_n689_), .A3(G15gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n688_), .B2(G15gat), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n692_));
  OR3_X1    g491(.A1(new_n690_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n694_));
  OR3_X1    g493(.A1(new_n653_), .A2(G15gat), .A3(new_n661_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n693_), .A2(new_n694_), .A3(new_n695_), .ZN(G1326gat));
  OR3_X1    g495(.A1(new_n653_), .A2(G22gat), .A3(new_n321_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n671_), .A2(new_n528_), .A3(new_n674_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT42), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n698_), .A2(new_n699_), .A3(G22gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n698_), .B2(G22gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n697_), .B1(new_n700_), .B2(new_n701_), .ZN(G1327gat));
  NOR3_X1   g501(.A1(new_n635_), .A2(new_n664_), .A3(new_n650_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n541_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(G29gat), .B1(new_n705_), .B2(new_n347_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n673_), .A2(new_n650_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n592_), .A2(new_n596_), .ZN(new_n708_));
  AOI211_X1 g507(.A(KEYINPUT43), .B(new_n708_), .C1(new_n535_), .C2(new_n540_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n710_), .B1(new_n663_), .B2(new_n597_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n709_), .B2(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(KEYINPUT44), .B1(new_n712_), .B2(KEYINPUT111), .ZN(new_n713_));
  INV_X1    g512(.A(new_n707_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n662_), .A2(new_n658_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n520_), .A2(KEYINPUT106), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n597_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT43), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n663_), .A2(new_n710_), .A3(new_n597_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n714_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT111), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  AOI22_X1  g521(.A1(new_n713_), .A2(new_n722_), .B1(KEYINPUT44), .B2(new_n720_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n347_), .A2(G29gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n706_), .B1(new_n723_), .B2(new_n724_), .ZN(G1328gat));
  NOR2_X1   g524(.A1(new_n486_), .A2(G36gat), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  OR3_X1    g526(.A1(new_n704_), .A2(KEYINPUT45), .A3(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(KEYINPUT45), .B1(new_n704_), .B2(new_n727_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  OAI211_X1 g529(.A(KEYINPUT44), .B(new_n707_), .C1(new_n709_), .C2(new_n711_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(new_n533_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n713_), .B2(new_n722_), .ZN(new_n733_));
  INV_X1    g532(.A(G36gat), .ZN(new_n734_));
  OAI211_X1 g533(.A(KEYINPUT46), .B(new_n730_), .C1(new_n733_), .C2(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n486_), .B1(new_n720_), .B2(KEYINPUT44), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n737_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n738_));
  AOI211_X1 g537(.A(KEYINPUT111), .B(new_n714_), .C1(new_n718_), .C2(new_n719_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n736_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  AOI22_X1  g539(.A1(new_n740_), .A2(G36gat), .B1(new_n729_), .B2(new_n728_), .ZN(new_n741_));
  XOR2_X1   g540(.A(KEYINPUT112), .B(KEYINPUT46), .Z(new_n742_));
  OAI21_X1  g541(.A(new_n735_), .B1(new_n741_), .B2(new_n742_), .ZN(G1329gat));
  INV_X1    g542(.A(G43gat), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n661_), .A2(new_n744_), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n731_), .B(new_n745_), .C1(new_n738_), .C2(new_n739_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n744_), .B1(new_n704_), .B2(new_n661_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT47), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT47), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n746_), .A2(new_n750_), .A3(new_n747_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(G1330gat));
  AOI21_X1  g551(.A(G50gat), .B1(new_n705_), .B2(new_n528_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n528_), .A2(G50gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n723_), .B2(new_n754_), .ZN(G1331gat));
  NOR3_X1   g554(.A1(new_n672_), .A2(new_n236_), .A3(new_n651_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n671_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n347_), .A2(G57gat), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n759_), .A2(KEYINPUT113), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n757_), .A2(new_n761_), .A3(new_n758_), .ZN(new_n762_));
  AOI211_X1 g561(.A(new_n236_), .B(new_n672_), .C1(new_n535_), .C2(new_n540_), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n763_), .A2(new_n650_), .A3(new_n708_), .ZN(new_n764_));
  AOI21_X1  g563(.A(G57gat), .B1(new_n764_), .B2(new_n347_), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n760_), .A2(new_n762_), .A3(new_n765_), .ZN(G1332gat));
  INV_X1    g565(.A(G64gat), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n764_), .A2(new_n767_), .A3(new_n533_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n671_), .A2(new_n533_), .A3(new_n756_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(G64gat), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n770_), .A2(KEYINPUT48), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n770_), .A2(KEYINPUT48), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(G1333gat));
  NAND3_X1  g572(.A1(new_n764_), .A2(new_n504_), .A3(new_n539_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n671_), .A2(new_n539_), .A3(new_n756_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(G71gat), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n776_), .A2(KEYINPUT49), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(KEYINPUT49), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n774_), .B1(new_n777_), .B2(new_n778_), .ZN(G1334gat));
  NAND3_X1  g578(.A1(new_n764_), .A2(new_n599_), .A3(new_n528_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n528_), .B(new_n756_), .C1(new_n668_), .C2(new_n670_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n781_), .A2(new_n782_), .A3(G78gat), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n781_), .B2(G78gat), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n780_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT114), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n787_), .B(new_n780_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(G1335gat));
  NAND3_X1  g588(.A1(new_n635_), .A2(new_n237_), .A3(new_n651_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(G85gat), .B1(new_n792_), .B2(new_n487_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n664_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n763_), .A2(new_n651_), .A3(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n795_), .A2(new_n548_), .A3(new_n347_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n793_), .A2(new_n796_), .ZN(G1336gat));
  OAI21_X1  g596(.A(G92gat), .B1(new_n792_), .B2(new_n486_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n795_), .A2(new_n549_), .A3(new_n533_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(G1337gat));
  NOR2_X1   g599(.A1(new_n661_), .A2(new_n566_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n795_), .A2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n494_), .B1(new_n791_), .B2(new_n539_), .ZN(new_n803_));
  OAI22_X1  g602(.A1(new_n802_), .A2(new_n803_), .B1(KEYINPUT115), .B2(KEYINPUT51), .ZN(new_n804_));
  NAND2_X1  g603(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n804_), .B(new_n805_), .ZN(G1338gat));
  INV_X1    g605(.A(G106gat), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n795_), .A2(new_n807_), .A3(new_n528_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n790_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n528_), .B(new_n809_), .C1(new_n709_), .C2(new_n711_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n811_));
  AND4_X1   g610(.A1(KEYINPUT116), .A2(new_n810_), .A3(new_n811_), .A4(G106gat), .ZN(new_n812_));
  OAI21_X1  g611(.A(G106gat), .B1(new_n811_), .B2(KEYINPUT116), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  AOI22_X1  g613(.A1(new_n810_), .A2(new_n814_), .B1(KEYINPUT116), .B2(new_n811_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n808_), .B1(new_n812_), .B2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT53), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n818_), .B(new_n808_), .C1(new_n812_), .C2(new_n815_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(G1339gat));
  NAND4_X1  g619(.A1(new_n708_), .A2(new_n672_), .A3(new_n237_), .A4(new_n650_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n821_), .B(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n235_), .B1(new_n227_), .B2(new_n223_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT119), .ZN(new_n826_));
  AOI22_X1  g625(.A1(new_n825_), .A2(new_n826_), .B1(new_n228_), .B2(new_n222_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n826_), .B2(new_n825_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n225_), .A2(new_n226_), .A3(new_n229_), .A4(new_n235_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT120), .B1(new_n632_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n830_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT120), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n832_), .B(new_n833_), .C1(new_n630_), .C2(new_n631_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n831_), .A2(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT55), .B1(new_n617_), .B2(KEYINPUT117), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n836_), .B1(KEYINPUT55), .B2(new_n617_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n616_), .A2(new_n620_), .A3(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n836_), .B1(new_n616_), .B2(new_n620_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT118), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n616_), .A2(new_n620_), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n843_), .B(new_n839_), .C1(new_n844_), .C2(new_n836_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n629_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n842_), .A2(new_n845_), .A3(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT56), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n842_), .A2(new_n845_), .A3(KEYINPUT56), .A4(new_n846_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n630_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n835_), .B1(new_n851_), .B2(new_n236_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n824_), .B1(new_n852_), .B2(new_n794_), .ZN(new_n853_));
  AOI211_X1 g652(.A(new_n630_), .B(new_n237_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n854_));
  OAI211_X1 g653(.A(KEYINPUT57), .B(new_n664_), .C1(new_n854_), .C2(new_n835_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n853_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT58), .B1(new_n851_), .B2(new_n832_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n708_), .ZN(new_n859_));
  AOI211_X1 g658(.A(new_n630_), .B(new_n830_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n597_), .B(KEYINPUT121), .C1(new_n860_), .C2(KEYINPUT58), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(KEYINPUT58), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n859_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n856_), .A2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n823_), .B1(new_n864_), .B2(new_n651_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n539_), .A2(new_n347_), .A3(new_n534_), .ZN(new_n866_));
  XOR2_X1   g665(.A(new_n866_), .B(KEYINPUT122), .Z(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n865_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(G113gat), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n869_), .A2(new_n870_), .A3(new_n236_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(KEYINPUT59), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(new_n865_), .B2(new_n868_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n237_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n871_), .B1(new_n875_), .B2(new_n870_), .ZN(G1340gat));
  XNOR2_X1  g675(.A(KEYINPUT123), .B(G120gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(new_n672_), .B2(KEYINPUT60), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n869_), .B(new_n878_), .C1(KEYINPUT60), .C2(new_n877_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n672_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(new_n877_), .ZN(G1341gat));
  INV_X1    g680(.A(new_n823_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n853_), .A2(new_n855_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n861_), .A2(new_n862_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n883_), .B1(new_n884_), .B2(new_n859_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n882_), .B1(new_n885_), .B2(new_n650_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n886_), .A2(new_n650_), .A3(new_n867_), .ZN(new_n887_));
  INV_X1    g686(.A(G127gat), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT124), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n887_), .A2(KEYINPUT124), .A3(new_n888_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n872_), .A2(new_n874_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n650_), .A2(G127gat), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n891_), .A2(new_n892_), .B1(new_n893_), .B2(new_n895_), .ZN(G1342gat));
  INV_X1    g695(.A(G134gat), .ZN(new_n897_));
  INV_X1    g696(.A(new_n666_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n869_), .A2(new_n897_), .A3(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n708_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(new_n897_), .ZN(G1343gat));
  NAND3_X1  g700(.A1(new_n661_), .A2(new_n347_), .A3(new_n537_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n865_), .A2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n236_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n635_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g706(.A1(new_n903_), .A2(new_n650_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT61), .B(G155gat), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(G1346gat));
  INV_X1    g709(.A(G162gat), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n903_), .A2(new_n911_), .A3(new_n898_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n903_), .A2(new_n597_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n912_), .B1(new_n914_), .B2(new_n911_), .ZN(G1347gat));
  NOR4_X1   g714(.A1(new_n661_), .A2(new_n347_), .A3(new_n528_), .A4(new_n486_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n886_), .A2(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(G169gat), .B1(new_n917_), .B2(new_n237_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n886_), .A2(new_n916_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n921_), .A2(new_n409_), .A3(new_n236_), .ZN(new_n922_));
  OAI211_X1 g721(.A(KEYINPUT62), .B(G169gat), .C1(new_n917_), .C2(new_n237_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n920_), .A2(new_n922_), .A3(new_n923_), .ZN(G1348gat));
  NAND3_X1  g723(.A1(new_n886_), .A2(new_n635_), .A3(new_n916_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g725(.A1(new_n886_), .A2(new_n650_), .A3(new_n916_), .ZN(new_n927_));
  MUX2_X1   g726(.A(new_n375_), .B(G183gat), .S(new_n927_), .Z(G1350gat));
  NAND3_X1  g727(.A1(new_n921_), .A2(new_n412_), .A3(new_n898_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n921_), .A2(new_n597_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n930_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n929_), .B1(new_n931_), .B2(new_n361_), .ZN(G1351gat));
  INV_X1    g731(.A(KEYINPUT125), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n528_), .A2(new_n487_), .A3(new_n533_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n539_), .A2(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n935_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n933_), .B1(new_n865_), .B2(new_n936_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n650_), .B1(new_n856_), .B2(new_n863_), .ZN(new_n938_));
  OAI211_X1 g737(.A(KEYINPUT125), .B(new_n935_), .C1(new_n938_), .C2(new_n823_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n937_), .A2(new_n939_), .ZN(new_n940_));
  AOI21_X1  g739(.A(G197gat), .B1(new_n940_), .B2(new_n236_), .ZN(new_n941_));
  AOI211_X1 g740(.A(new_n276_), .B(new_n237_), .C1(new_n937_), .C2(new_n939_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n941_), .A2(new_n942_), .ZN(G1352gat));
  AOI21_X1  g742(.A(KEYINPUT125), .B1(new_n886_), .B2(new_n935_), .ZN(new_n944_));
  INV_X1    g743(.A(new_n939_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n635_), .B1(new_n944_), .B2(new_n945_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(KEYINPUT126), .B(G204gat), .ZN(new_n947_));
  INV_X1    g746(.A(new_n947_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n946_), .A2(new_n948_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n940_), .A2(new_n635_), .A3(new_n947_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n949_), .A2(new_n950_), .ZN(G1353gat));
  OR2_X1    g750(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n952_), .B1(new_n940_), .B2(new_n650_), .ZN(new_n953_));
  XNOR2_X1  g752(.A(KEYINPUT63), .B(G211gat), .ZN(new_n954_));
  AOI211_X1 g753(.A(new_n651_), .B(new_n954_), .C1(new_n937_), .C2(new_n939_), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n953_), .A2(new_n955_), .ZN(G1354gat));
  NAND2_X1  g755(.A1(new_n940_), .A2(new_n898_), .ZN(new_n957_));
  INV_X1    g756(.A(G218gat), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n597_), .A2(G218gat), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n959_), .B(KEYINPUT127), .ZN(new_n960_));
  AOI22_X1  g759(.A1(new_n957_), .A2(new_n958_), .B1(new_n940_), .B2(new_n960_), .ZN(G1355gat));
endmodule


