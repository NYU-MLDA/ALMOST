//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 1 1 0 1 0 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n842_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n885_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT20), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G197gat), .A2(G204gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT91), .B(G197gat), .ZN(new_n206_));
  INV_X1    g005(.A(G204gat), .ZN(new_n207_));
  OAI211_X1 g006(.A(KEYINPUT92), .B(new_n205_), .C1(new_n206_), .C2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT21), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n208_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT91), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n213_), .A2(G197gat), .ZN(new_n214_));
  INV_X1    g013(.A(G197gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n215_), .A2(KEYINPUT91), .ZN(new_n216_));
  OAI21_X1  g015(.A(G204gat), .B1(new_n214_), .B2(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(KEYINPUT92), .B1(new_n217_), .B2(new_n205_), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT93), .B1(new_n212_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT92), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n215_), .A2(KEYINPUT91), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n213_), .A2(G197gat), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n207_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n220_), .B1(new_n223_), .B2(new_n204_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT93), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n224_), .A2(new_n225_), .A3(new_n208_), .A4(new_n211_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n219_), .A2(new_n226_), .ZN(new_n227_));
  XOR2_X1   g026(.A(G211gat), .B(G218gat), .Z(new_n228_));
  NAND3_X1  g027(.A1(new_n221_), .A2(new_n222_), .A3(new_n207_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n210_), .B1(G197gat), .B2(G204gat), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n228_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n210_), .B1(new_n223_), .B2(new_n204_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n227_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT82), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT22), .B(G169gat), .ZN(new_n237_));
  INV_X1    g036(.A(G176gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT23), .ZN(new_n241_));
  OR2_X1    g040(.A1(G183gat), .A2(G190gat), .ZN(new_n242_));
  AOI22_X1  g041(.A1(new_n236_), .A2(new_n239_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n237_), .A2(KEYINPUT82), .A3(new_n238_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G169gat), .A2(G176gat), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  OR2_X1    g045(.A1(G169gat), .A2(G176gat), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n247_), .A2(KEYINPUT24), .A3(new_n245_), .ZN(new_n248_));
  OR3_X1    g047(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n241_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(G183gat), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT81), .B1(new_n251_), .B2(KEYINPUT25), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT26), .B(G190gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT25), .B(G183gat), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n252_), .B(new_n253_), .C1(new_n254_), .C2(KEYINPUT81), .ZN(new_n255_));
  AOI22_X1  g054(.A1(new_n243_), .A2(new_n246_), .B1(new_n250_), .B2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n203_), .B1(new_n235_), .B2(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n233_), .B1(new_n219_), .B2(new_n226_), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n248_), .A2(new_n249_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n254_), .A2(new_n253_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n261_), .A2(new_n241_), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n239_), .A2(new_n245_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n241_), .A2(new_n242_), .ZN(new_n264_));
  AOI22_X1  g063(.A1(new_n260_), .A2(new_n262_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n259_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n258_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G226gat), .A2(G233gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n202_), .B1(new_n267_), .B2(new_n271_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n258_), .A2(KEYINPUT98), .A3(new_n270_), .A4(new_n266_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n265_), .B1(new_n227_), .B2(new_n234_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n203_), .B1(new_n259_), .B2(new_n256_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT96), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n275_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(G218gat), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n279_), .A2(G211gat), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(G211gat), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT21), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n221_), .A2(new_n222_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n204_), .B1(new_n283_), .B2(G204gat), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n282_), .B1(new_n284_), .B2(KEYINPUT92), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n225_), .B1(new_n285_), .B2(new_n224_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n226_), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n256_), .B(new_n234_), .C1(new_n286_), .C2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT20), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT96), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n278_), .A2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(KEYINPUT97), .B1(new_n291_), .B2(new_n271_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT97), .ZN(new_n293_));
  AOI211_X1 g092(.A(new_n293_), .B(new_n270_), .C1(new_n278_), .C2(new_n290_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n274_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G8gat), .B(G36gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT18), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G64gat), .B(G92gat), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n297_), .B(new_n298_), .Z(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n295_), .A2(new_n300_), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n299_), .B(new_n274_), .C1(new_n292_), .C2(new_n294_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT27), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n267_), .A2(new_n271_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT102), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n278_), .A2(new_n270_), .A3(new_n290_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT102), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n267_), .A2(new_n309_), .A3(new_n271_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n307_), .A2(new_n308_), .A3(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n304_), .B1(new_n311_), .B2(new_n300_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(new_n302_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n305_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(G233gat), .ZN(new_n316_));
  OR2_X1    g115(.A1(KEYINPUT90), .A2(G228gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(KEYINPUT90), .A2(G228gat), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n316_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n259_), .A2(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(G155gat), .B(G162gat), .Z(new_n321_));
  NAND2_X1  g120(.A1(G141gat), .A2(G148gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT2), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n325_));
  NOR3_X1   g124(.A1(KEYINPUT86), .A2(G141gat), .A3(G148gat), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT3), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n324_), .B(new_n325_), .C1(new_n326_), .C2(new_n327_), .ZN(new_n328_));
  OR2_X1    g127(.A1(G141gat), .A2(G148gat), .ZN(new_n329_));
  NOR3_X1   g128(.A1(new_n329_), .A2(KEYINPUT86), .A3(KEYINPUT3), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n321_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT87), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  OAI211_X1 g132(.A(KEYINPUT87), .B(new_n321_), .C1(new_n328_), .C2(new_n330_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT1), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n321_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n336_), .A2(new_n329_), .A3(new_n322_), .A4(new_n337_), .ZN(new_n338_));
  AND3_X1   g137(.A1(new_n333_), .A2(new_n334_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT29), .ZN(new_n340_));
  NOR3_X1   g139(.A1(new_n339_), .A2(KEYINPUT89), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT89), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n333_), .A2(new_n334_), .A3(new_n338_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n342_), .B1(new_n343_), .B2(KEYINPUT29), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n320_), .B1(new_n341_), .B2(new_n344_), .ZN(new_n345_));
  XOR2_X1   g144(.A(G78gat), .B(G106gat), .Z(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n339_), .A2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n319_), .B1(new_n349_), .B2(new_n259_), .ZN(new_n350_));
  AND3_X1   g149(.A1(new_n345_), .A2(new_n347_), .A3(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n347_), .B1(new_n345_), .B2(new_n350_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n339_), .A2(new_n340_), .ZN(new_n354_));
  XOR2_X1   g153(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n355_));
  OR2_X1    g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(G22gat), .B(G50gat), .Z(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n354_), .A2(new_n355_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n356_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n358_), .B1(new_n356_), .B2(new_n359_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  OR2_X1    g161(.A1(new_n353_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n353_), .A2(new_n362_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G127gat), .B(G134gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT84), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT84), .ZN(new_n368_));
  INV_X1    g167(.A(G127gat), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n369_), .A2(G134gat), .ZN(new_n370_));
  INV_X1    g169(.A(G134gat), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n371_), .A2(G127gat), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n368_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G113gat), .B(G120gat), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n367_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n374_), .B1(new_n367_), .B2(new_n373_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n343_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n377_), .A2(new_n334_), .A3(new_n338_), .A4(new_n333_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G225gat), .A2(G233gat), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n383_), .B(KEYINPUT100), .Z(new_n384_));
  NOR3_X1   g183(.A1(new_n380_), .A2(new_n382_), .A3(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n379_), .A2(KEYINPUT4), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n379_), .A2(KEYINPUT4), .A3(new_n381_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT99), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT99), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n379_), .A2(new_n389_), .A3(new_n381_), .A4(KEYINPUT4), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n386_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n385_), .B1(new_n391_), .B2(new_n384_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G1gat), .B(G29gat), .ZN(new_n393_));
  INV_X1    g192(.A(G85gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT0), .B(G57gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n392_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n391_), .A2(new_n384_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n385_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n399_), .A2(new_n397_), .A3(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n398_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n377_), .B(KEYINPUT31), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G227gat), .A2(G233gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(G71gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(G99gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n256_), .B(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G15gat), .B(G43gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT83), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT30), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n408_), .B(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT85), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n404_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  OR3_X1    g213(.A1(new_n414_), .A2(new_n413_), .A3(new_n412_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n414_), .B1(new_n413_), .B2(new_n412_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n315_), .A2(new_n365_), .A3(new_n403_), .A4(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT27), .B1(new_n301_), .B2(new_n302_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n313_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n363_), .A2(new_n364_), .A3(new_n401_), .A4(new_n398_), .ZN(new_n422_));
  NOR3_X1   g221(.A1(new_n420_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT101), .ZN(new_n424_));
  INV_X1    g223(.A(new_n384_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n391_), .A2(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n380_), .A2(new_n382_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n397_), .B1(new_n427_), .B2(new_n384_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT33), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n392_), .A2(new_n430_), .A3(new_n397_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n430_), .B1(new_n392_), .B2(new_n397_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n429_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n424_), .B1(new_n303_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n401_), .A2(KEYINPUT33), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n392_), .A2(new_n430_), .A3(new_n397_), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n435_), .A2(new_n436_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n437_), .A2(KEYINPUT101), .A3(new_n302_), .A4(new_n301_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n299_), .A2(KEYINPUT32), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n311_), .A2(new_n439_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n402_), .B(new_n440_), .C1(new_n295_), .C2(new_n439_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n434_), .A2(new_n438_), .A3(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n423_), .B1(new_n442_), .B2(new_n365_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n419_), .B1(new_n443_), .B2(new_n418_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G1gat), .B(G8gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT76), .ZN(new_n447_));
  INV_X1    g246(.A(G15gat), .ZN(new_n448_));
  INV_X1    g247(.A(G22gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G15gat), .A2(G22gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G1gat), .A2(G8gat), .ZN(new_n452_));
  AOI22_X1  g251(.A1(new_n450_), .A2(new_n451_), .B1(KEYINPUT14), .B2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n447_), .B(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G29gat), .B(G36gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G43gat), .B(G50gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n454_), .A2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT80), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n454_), .A2(new_n457_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G229gat), .A2(G233gat), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n454_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n457_), .B(KEYINPUT15), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n459_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n464_), .B1(new_n463_), .B2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G113gat), .B(G141gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G169gat), .B(G197gat), .ZN(new_n470_));
  XOR2_X1   g269(.A(new_n469_), .B(new_n470_), .Z(new_n471_));
  XNOR2_X1  g270(.A(new_n468_), .B(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n445_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G120gat), .B(G148gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT5), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G176gat), .B(G204gat), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n476_), .B(new_n477_), .Z(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT64), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n480_), .A2(KEYINPUT9), .ZN(new_n481_));
  INV_X1    g280(.A(G92gat), .ZN(new_n482_));
  NOR3_X1   g281(.A1(new_n481_), .A2(new_n394_), .A3(new_n482_), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n480_), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n484_));
  XOR2_X1   g283(.A(KEYINPUT10), .B(G99gat), .Z(new_n485_));
  INV_X1    g284(.A(G106gat), .ZN(new_n486_));
  AOI22_X1  g285(.A1(new_n483_), .A2(new_n484_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G99gat), .A2(G106gat), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n487_), .B(new_n491_), .C1(new_n484_), .C2(new_n483_), .ZN(new_n492_));
  XOR2_X1   g291(.A(G85gat), .B(G92gat), .Z(new_n493_));
  NOR2_X1   g292(.A1(G99gat), .A2(G106gat), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT7), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n493_), .B1(new_n496_), .B2(new_n490_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT8), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n492_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n493_), .A2(KEYINPUT8), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT65), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n496_), .A2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n490_), .B1(new_n496_), .B2(new_n502_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n501_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n500_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT68), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G57gat), .B(G64gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT11), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT66), .ZN(new_n510_));
  XOR2_X1   g309(.A(G71gat), .B(G78gat), .Z(new_n511_));
  OAI21_X1  g310(.A(new_n511_), .B1(KEYINPUT11), .B2(new_n508_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n510_), .B(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n507_), .A2(KEYINPUT12), .A3(new_n514_), .ZN(new_n515_));
  AND2_X1   g314(.A1(G230gat), .A2(G233gat), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n516_), .B1(new_n506_), .B2(new_n513_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n506_), .A2(new_n513_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT70), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NOR3_X1   g322(.A1(new_n518_), .A2(KEYINPUT70), .A3(new_n520_), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n515_), .B(new_n517_), .C1(new_n523_), .C2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n506_), .A2(new_n513_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT67), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n516_), .B1(new_n528_), .B2(new_n518_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n479_), .B1(new_n525_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n525_), .A2(new_n529_), .A3(new_n479_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT72), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n532_), .A2(KEYINPUT71), .A3(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n533_), .B1(new_n532_), .B2(KEYINPUT71), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n531_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n532_), .A2(KEYINPUT71), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT72), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n532_), .A2(KEYINPUT71), .A3(new_n533_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n538_), .A2(new_n530_), .A3(new_n539_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n536_), .A2(new_n540_), .A3(KEYINPUT13), .ZN(new_n541_));
  AOI21_X1  g340(.A(KEYINPUT13), .B1(new_n536_), .B2(new_n540_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n543_), .A2(KEYINPUT73), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(KEYINPUT73), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n507_), .A2(new_n466_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G232gat), .A2(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n550_), .A2(KEYINPUT35), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n551_), .B1(new_n506_), .B2(new_n457_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n547_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n550_), .A2(KEYINPUT35), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(G190gat), .B(G218gat), .Z(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT75), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G134gat), .B(G162gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT36), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n555_), .A2(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n559_), .A2(KEYINPUT36), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n555_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT37), .ZN(new_n565_));
  XOR2_X1   g364(.A(G127gat), .B(G155gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(G183gat), .B(G211gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n570_), .A2(KEYINPUT17), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n571_), .A2(KEYINPUT78), .ZN(new_n572_));
  AND2_X1   g371(.A1(G231gat), .A2(G233gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n574_), .A2(new_n454_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n454_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(new_n514_), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n570_), .A2(KEYINPUT17), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n575_), .A2(new_n513_), .A3(new_n576_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n578_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT79), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT79), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n578_), .A2(new_n583_), .A3(new_n579_), .A4(new_n580_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n565_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n474_), .A2(new_n546_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT103), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n589_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n403_), .A2(G1gat), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n590_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT38), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n472_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT104), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n585_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n564_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n596_), .A2(new_n597_), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n598_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(new_n402_), .A3(new_n444_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(G1gat), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n593_), .A2(new_n594_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n595_), .A2(new_n605_), .A3(new_n606_), .ZN(G1324gat));
  NOR2_X1   g406(.A1(new_n315_), .A2(G8gat), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n590_), .A2(new_n591_), .A3(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n603_), .A2(new_n314_), .A3(new_n444_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n610_), .A2(new_n611_), .A3(G8gat), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n611_), .B1(new_n610_), .B2(G8gat), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n609_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT40), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n609_), .B(KEYINPUT40), .C1(new_n612_), .C2(new_n613_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1325gat));
  NAND2_X1  g417(.A1(new_n590_), .A2(new_n591_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n418_), .A2(new_n448_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n603_), .A2(new_n418_), .A3(new_n444_), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n621_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n622_));
  AOI21_X1  g421(.A(KEYINPUT41), .B1(new_n621_), .B2(G15gat), .ZN(new_n623_));
  OAI22_X1  g422(.A1(new_n619_), .A2(new_n620_), .B1(new_n622_), .B2(new_n623_), .ZN(G1326gat));
  INV_X1    g423(.A(new_n365_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(new_n449_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n603_), .A2(new_n625_), .A3(new_n444_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT42), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n627_), .A2(new_n628_), .A3(G22gat), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n628_), .B1(new_n627_), .B2(G22gat), .ZN(new_n630_));
  OAI22_X1  g429(.A1(new_n619_), .A2(new_n626_), .B1(new_n629_), .B2(new_n630_), .ZN(G1327gat));
  INV_X1    g430(.A(KEYINPUT43), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n564_), .B(KEYINPUT37), .Z(new_n633_));
  NAND2_X1  g432(.A1(new_n442_), .A2(new_n365_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n423_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n418_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  NOR4_X1   g435(.A1(new_n314_), .A2(new_n625_), .A3(new_n402_), .A4(new_n417_), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n632_), .B(new_n633_), .C1(new_n636_), .C2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT105), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT105), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n444_), .A2(new_n640_), .A3(new_n632_), .A4(new_n633_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n444_), .A2(new_n633_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT43), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n639_), .A2(new_n641_), .A3(new_n643_), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n598_), .A2(new_n599_), .A3(new_n602_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT44), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n644_), .A2(KEYINPUT44), .A3(new_n645_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(G29gat), .B1(new_n650_), .B2(new_n403_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n543_), .A2(new_n585_), .A3(new_n564_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n474_), .A2(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n403_), .A2(G29gat), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT106), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n651_), .A2(new_n656_), .ZN(G1328gat));
  INV_X1    g456(.A(KEYINPUT107), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n315_), .A2(G36gat), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n474_), .A2(new_n658_), .A3(new_n652_), .A4(new_n659_), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n652_), .A2(new_n472_), .A3(new_n444_), .A4(new_n659_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT107), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT45), .ZN(new_n664_));
  AND3_X1   g463(.A1(new_n644_), .A2(KEYINPUT44), .A3(new_n645_), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT44), .B1(new_n644_), .B2(new_n645_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n665_), .A2(new_n666_), .A3(new_n315_), .ZN(new_n667_));
  INV_X1    g466(.A(G36gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n664_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT46), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  OAI211_X1 g470(.A(KEYINPUT46), .B(new_n664_), .C1(new_n667_), .C2(new_n668_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1329gat));
  AND2_X1   g472(.A1(new_n653_), .A2(new_n418_), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n674_), .A2(G43gat), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n418_), .A2(G43gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n650_), .B2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT47), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT47), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n675_), .B(new_n679_), .C1(new_n650_), .C2(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(G1330gat));
  INV_X1    g480(.A(G50gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n653_), .A2(new_n682_), .A3(new_n625_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n650_), .A2(new_n365_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n684_), .A2(KEYINPUT108), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n648_), .A2(KEYINPUT108), .A3(new_n625_), .A4(new_n649_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(G50gat), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n683_), .B1(new_n685_), .B2(new_n687_), .ZN(G1331gat));
  INV_X1    g487(.A(new_n546_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n445_), .A2(new_n472_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n689_), .A2(new_n690_), .A3(new_n601_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(KEYINPUT111), .B(G57gat), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n691_), .A2(new_n403_), .A3(new_n692_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT112), .Z(new_n694_));
  AND3_X1   g493(.A1(new_n444_), .A2(KEYINPUT109), .A3(new_n473_), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT109), .B1(new_n444_), .B2(new_n473_), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n697_), .A2(new_n543_), .A3(new_n587_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT110), .Z(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(new_n402_), .ZN(new_n700_));
  INV_X1    g499(.A(G57gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n694_), .B1(new_n700_), .B2(new_n701_), .ZN(G1332gat));
  OAI21_X1  g501(.A(G64gat), .B1(new_n691_), .B2(new_n315_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT48), .ZN(new_n704_));
  INV_X1    g503(.A(new_n699_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n315_), .A2(G64gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n704_), .B1(new_n705_), .B2(new_n706_), .ZN(G1333gat));
  OAI21_X1  g506(.A(G71gat), .B1(new_n691_), .B2(new_n417_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT49), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n417_), .A2(G71gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(new_n705_), .B2(new_n710_), .ZN(G1334gat));
  OAI21_X1  g510(.A(G78gat), .B1(new_n691_), .B2(new_n365_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT50), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n365_), .A2(G78gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n713_), .B1(new_n705_), .B2(new_n714_), .ZN(G1335gat));
  NOR2_X1   g514(.A1(new_n585_), .A2(new_n564_), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n544_), .A2(new_n545_), .A3(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n697_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n719_), .A2(new_n394_), .A3(new_n402_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n543_), .A2(new_n473_), .A3(new_n599_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT113), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n644_), .A2(KEYINPUT114), .A3(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT114), .B1(new_n644_), .B2(new_n722_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n723_), .A2(new_n724_), .A3(new_n403_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n720_), .B1(new_n725_), .B2(new_n394_), .ZN(G1336gat));
  INV_X1    g525(.A(KEYINPUT116), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n717_), .B(new_n314_), .C1(new_n695_), .C2(new_n696_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n482_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT115), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n314_), .A2(G92gat), .ZN(new_n731_));
  NOR3_X1   g530(.A1(new_n723_), .A2(new_n724_), .A3(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n727_), .B1(new_n730_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT115), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n729_), .B(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n732_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(new_n736_), .A3(KEYINPUT116), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n733_), .A2(new_n737_), .ZN(G1337gat));
  AND2_X1   g537(.A1(new_n418_), .A2(new_n485_), .ZN(new_n739_));
  AOI22_X1  g538(.A1(new_n719_), .A2(new_n739_), .B1(KEYINPUT117), .B2(KEYINPUT51), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n644_), .A2(new_n418_), .A3(new_n722_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(G99gat), .ZN(new_n742_));
  OR2_X1    g541(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n740_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n740_), .B2(new_n742_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1338gat));
  NAND3_X1  g545(.A1(new_n644_), .A2(new_n722_), .A3(new_n625_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n747_), .A2(new_n748_), .A3(G106gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n747_), .B2(G106gat), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n625_), .A2(new_n486_), .ZN(new_n751_));
  OAI22_X1  g550(.A1(new_n749_), .A2(new_n750_), .B1(new_n718_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT53), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT53), .ZN(new_n754_));
  OAI221_X1 g553(.A(new_n754_), .B1(new_n718_), .B2(new_n751_), .C1(new_n749_), .C2(new_n750_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1339gat));
  NOR4_X1   g555(.A1(new_n314_), .A2(new_n625_), .A3(new_n403_), .A4(new_n417_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n515_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n516_), .B1(new_n759_), .B2(new_n528_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n521_), .B(new_n522_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n761_), .A2(KEYINPUT55), .A3(new_n515_), .A4(new_n517_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT55), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n525_), .A2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n760_), .A2(new_n762_), .A3(new_n764_), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n765_), .A2(KEYINPUT56), .A3(new_n478_), .ZN(new_n766_));
  AOI21_X1  g565(.A(KEYINPUT56), .B1(new_n765_), .B2(new_n478_), .ZN(new_n767_));
  OR2_X1    g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT118), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n468_), .A2(new_n471_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n467_), .A2(new_n463_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n471_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n772_), .B1(new_n461_), .B2(new_n463_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n769_), .B1(new_n770_), .B2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n468_), .A2(new_n471_), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n776_), .B(KEYINPUT118), .C1(new_n771_), .C2(new_n773_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n768_), .A2(KEYINPUT58), .A3(new_n532_), .A4(new_n778_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n778_), .B(new_n532_), .C1(new_n766_), .C2(new_n767_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT58), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n633_), .A2(new_n779_), .A3(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT57), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n472_), .B(new_n532_), .C1(new_n766_), .C2(new_n767_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n536_), .A2(new_n540_), .A3(new_n778_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n784_), .B1(new_n787_), .B2(new_n564_), .ZN(new_n788_));
  AOI211_X1 g587(.A(KEYINPUT57), .B(new_n600_), .C1(new_n785_), .C2(new_n786_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n783_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT119), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT119), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n783_), .B(new_n792_), .C1(new_n788_), .C2(new_n789_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n791_), .A2(new_n599_), .A3(new_n793_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n586_), .A2(new_n543_), .A3(new_n472_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n795_), .B(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n758_), .B1(new_n794_), .B2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(G113gat), .B1(new_n798_), .B2(new_n472_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n794_), .A2(new_n797_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n757_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT59), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT59), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n803_), .B1(new_n757_), .B2(KEYINPUT120), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(KEYINPUT120), .B2(new_n757_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n795_), .B(KEYINPUT54), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n790_), .A2(new_n599_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n805_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n802_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(G113gat), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n472_), .B2(KEYINPUT121), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(KEYINPUT121), .B2(new_n811_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n799_), .B1(new_n810_), .B2(new_n813_), .ZN(G1340gat));
  NOR3_X1   g613(.A1(new_n541_), .A2(new_n542_), .A3(KEYINPUT60), .ZN(new_n815_));
  INV_X1    g614(.A(G120gat), .ZN(new_n816_));
  MUX2_X1   g615(.A(KEYINPUT60), .B(new_n815_), .S(new_n816_), .Z(new_n817_));
  NAND2_X1  g616(.A1(new_n798_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT122), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n818_), .B(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n802_), .A2(new_n689_), .A3(new_n808_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n820_), .B1(new_n822_), .B2(new_n816_), .ZN(G1341gat));
  OAI21_X1  g622(.A(new_n369_), .B1(new_n801_), .B2(new_n599_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n599_), .A2(new_n369_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n808_), .B(new_n825_), .C1(new_n798_), .C2(new_n803_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT123), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n824_), .A2(KEYINPUT123), .A3(new_n826_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(G1342gat));
  OAI21_X1  g630(.A(G134gat), .B1(new_n809_), .B2(new_n565_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n798_), .A2(new_n371_), .A3(new_n600_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(G1343gat));
  NOR2_X1   g633(.A1(new_n418_), .A2(new_n365_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n314_), .A2(new_n403_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  AOI211_X1 g637(.A(new_n836_), .B(new_n838_), .C1(new_n794_), .C2(new_n797_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n472_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n689_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g642(.A(KEYINPUT61), .B(G155gat), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT124), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n846_), .B1(new_n839_), .B2(new_n585_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n800_), .A2(new_n585_), .A3(new_n835_), .A4(new_n837_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n848_), .A2(KEYINPUT124), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n845_), .B1(new_n847_), .B2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n839_), .A2(new_n846_), .A3(new_n585_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n848_), .A2(KEYINPUT124), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n852_), .A3(new_n844_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n850_), .A2(new_n853_), .ZN(G1346gat));
  AOI21_X1  g653(.A(G162gat), .B1(new_n839_), .B2(new_n600_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n633_), .A2(G162gat), .ZN(new_n856_));
  XOR2_X1   g655(.A(new_n856_), .B(KEYINPUT125), .Z(new_n857_));
  AOI21_X1  g656(.A(new_n855_), .B1(new_n839_), .B2(new_n857_), .ZN(G1347gat));
  NOR2_X1   g657(.A1(new_n806_), .A2(new_n807_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n315_), .A2(new_n402_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n418_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n365_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n859_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n472_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(G169gat), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n864_), .A2(new_n472_), .A3(new_n237_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n865_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n868_), .A2(new_n869_), .A3(new_n870_), .ZN(G1348gat));
  AOI21_X1  g670(.A(G176gat), .B1(new_n864_), .B2(new_n543_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n800_), .A2(new_n365_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(KEYINPUT126), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT126), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n800_), .A2(new_n875_), .A3(new_n365_), .ZN(new_n876_));
  AND3_X1   g675(.A1(new_n874_), .A2(new_n862_), .A3(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n546_), .A2(new_n238_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n872_), .B1(new_n877_), .B2(new_n878_), .ZN(G1349gat));
  INV_X1    g678(.A(new_n864_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n880_), .A2(new_n254_), .A3(new_n599_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n874_), .A2(new_n585_), .A3(new_n862_), .A4(new_n876_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n881_), .B1(new_n882_), .B2(new_n251_), .ZN(G1350gat));
  OAI21_X1  g682(.A(G190gat), .B1(new_n880_), .B2(new_n565_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n864_), .A2(new_n253_), .A3(new_n600_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1351gat));
  NAND3_X1  g685(.A1(new_n800_), .A2(new_n835_), .A3(new_n860_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(KEYINPUT127), .A2(G197gat), .ZN(new_n889_));
  OR2_X1    g688(.A1(KEYINPUT127), .A2(G197gat), .ZN(new_n890_));
  AOI22_X1  g689(.A1(new_n888_), .A2(new_n472_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n887_), .A2(new_n473_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(new_n890_), .ZN(G1352gat));
  NOR2_X1   g692(.A1(new_n887_), .A2(new_n546_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(new_n207_), .ZN(G1353gat));
  NOR2_X1   g694(.A1(new_n887_), .A2(new_n599_), .ZN(new_n896_));
  OR2_X1    g695(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  XOR2_X1   g697(.A(KEYINPUT63), .B(G211gat), .Z(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n896_), .B2(new_n899_), .ZN(G1354gat));
  OAI21_X1  g699(.A(G218gat), .B1(new_n887_), .B2(new_n565_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n600_), .A2(new_n279_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n887_), .B2(new_n902_), .ZN(G1355gat));
endmodule


