//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n590_, new_n591_, new_n592_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n790_, new_n791_, new_n793_, new_n794_,
    new_n795_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n819_, new_n820_, new_n821_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_;
  INV_X1    g000(.A(G141gat), .ZN(new_n202_));
  INV_X1    g001(.A(G148gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT84), .ZN(new_n204_));
  OAI211_X1 g003(.A(new_n202_), .B(new_n203_), .C1(new_n204_), .C2(KEYINPUT3), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n206_));
  OAI211_X1 g005(.A(new_n206_), .B(KEYINPUT84), .C1(G141gat), .C2(G148gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT85), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT2), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n209_), .A2(new_n210_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n204_), .A2(KEYINPUT3), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n208_), .A2(new_n212_), .A3(new_n214_), .A4(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G155gat), .B(G162gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT86), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n217_), .A2(KEYINPUT1), .ZN(new_n221_));
  AND2_X1   g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222_));
  AOI22_X1  g021(.A1(new_n222_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n202_), .A2(new_n203_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n221_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT86), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n216_), .A2(new_n226_), .A3(new_n218_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n220_), .A2(new_n225_), .A3(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n228_), .A2(KEYINPUT29), .ZN(new_n229_));
  XOR2_X1   g028(.A(new_n229_), .B(KEYINPUT89), .Z(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT88), .B(G204gat), .ZN(new_n231_));
  INV_X1    g030(.A(G197gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(G204gat), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n233_), .B(KEYINPUT21), .C1(new_n232_), .C2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G211gat), .B(G218gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n231_), .A2(G197gat), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n237_), .B1(G197gat), .B2(new_n234_), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n235_), .B(new_n236_), .C1(new_n238_), .C2(KEYINPUT21), .ZN(new_n239_));
  INV_X1    g038(.A(new_n236_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(KEYINPUT21), .A3(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n243_), .B1(KEYINPUT29), .B2(new_n228_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n230_), .B(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G22gat), .B(G50gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G78gat), .B(G106gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G228gat), .A2(G233gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n248_), .B(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n245_), .B(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G226gat), .A2(G233gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT19), .ZN(new_n256_));
  INV_X1    g055(.A(G183gat), .ZN(new_n257_));
  INV_X1    g056(.A(G190gat), .ZN(new_n258_));
  OR3_X1    g057(.A1(new_n257_), .A2(new_n258_), .A3(KEYINPUT23), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT23), .B1(new_n257_), .B2(new_n258_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT79), .ZN(new_n262_));
  INV_X1    g061(.A(G169gat), .ZN(new_n263_));
  INV_X1    g062(.A(G176gat), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n262_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT79), .B1(G169gat), .B2(G176gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT24), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n261_), .A2(new_n269_), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n270_), .A2(KEYINPUT91), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT25), .B(G183gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(G190gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT24), .B1(new_n263_), .B2(new_n264_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n276_), .A2(KEYINPUT90), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(KEYINPUT90), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n277_), .A2(new_n265_), .A3(new_n266_), .A4(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n270_), .A2(KEYINPUT91), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n271_), .A2(new_n274_), .A3(new_n279_), .A4(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n263_), .A2(new_n264_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT22), .B(G169gat), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n282_), .B1(new_n283_), .B2(new_n264_), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n260_), .B(KEYINPUT81), .Z(new_n285_));
  INV_X1    g084(.A(new_n259_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n284_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n281_), .A2(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT20), .B1(new_n290_), .B2(new_n242_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n287_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n267_), .A2(new_n275_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT80), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n292_), .A2(new_n294_), .A3(new_n269_), .A4(new_n274_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n261_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n284_), .B1(new_n296_), .B2(new_n288_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n243_), .B1(new_n295_), .B2(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n256_), .B1(new_n291_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n290_), .A2(new_n242_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n295_), .A2(new_n243_), .A3(new_n297_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n300_), .A2(new_n301_), .A3(KEYINPUT20), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n299_), .B1(new_n302_), .B2(new_n256_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G64gat), .B(G92gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G8gat), .B(G36gat), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n306_), .B(new_n307_), .Z(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n303_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n256_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n311_), .B1(new_n291_), .B2(new_n298_), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n300_), .A2(new_n301_), .A3(KEYINPUT20), .A4(new_n256_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(new_n308_), .ZN(new_n315_));
  AND3_X1   g114(.A1(new_n310_), .A2(KEYINPUT27), .A3(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(KEYINPUT98), .B(KEYINPUT27), .Z(new_n317_));
  NAND3_X1  g116(.A1(new_n312_), .A2(new_n313_), .A3(new_n309_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n317_), .B1(new_n315_), .B2(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT100), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NOR3_X1   g121(.A1(new_n316_), .A2(KEYINPUT100), .A3(new_n319_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n254_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(G113gat), .B(G120gat), .Z(new_n325_));
  XNOR2_X1  g124(.A(G127gat), .B(G134gat), .ZN(new_n326_));
  OR2_X1    g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n326_), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n327_), .A2(new_n328_), .A3(KEYINPUT83), .ZN(new_n329_));
  AOI21_X1  g128(.A(KEYINPUT83), .B1(new_n327_), .B2(new_n328_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT4), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n228_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT95), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT93), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n216_), .A2(new_n226_), .A3(new_n218_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n226_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n221_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n340_));
  NOR3_X1   g139(.A1(new_n338_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G113gat), .B(G120gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n326_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT83), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n337_), .B1(new_n341_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n341_), .A2(new_n343_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n228_), .A2(new_n331_), .A3(KEYINPUT93), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n345_), .A2(KEYINPUT4), .A3(new_n346_), .A4(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT94), .ZN(new_n349_));
  AND2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n348_), .A2(new_n349_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n336_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G225gat), .A2(G233gat), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n228_), .A2(KEYINPUT93), .A3(new_n331_), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT93), .B1(new_n228_), .B2(new_n331_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(new_n346_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n353_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G1gat), .B(G29gat), .ZN(new_n361_));
  INV_X1    g160(.A(G85gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT0), .B(G57gat), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n363_), .B(new_n364_), .Z(new_n365_));
  NAND4_X1  g164(.A1(new_n355_), .A2(KEYINPUT97), .A3(new_n360_), .A4(new_n365_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n358_), .A2(KEYINPUT94), .A3(KEYINPUT4), .A4(new_n346_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n348_), .A2(new_n349_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n335_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n360_), .B(new_n365_), .C1(new_n369_), .C2(new_n353_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT97), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n360_), .B1(new_n369_), .B2(new_n353_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n365_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n366_), .A2(new_n372_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G227gat), .A2(G233gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n344_), .B(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT82), .B(KEYINPUT30), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n295_), .A2(new_n297_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G15gat), .B(G43gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT31), .ZN(new_n384_));
  XOR2_X1   g183(.A(G71gat), .B(G99gat), .Z(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n382_), .B(new_n386_), .ZN(new_n387_));
  OR2_X1    g186(.A1(new_n381_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n381_), .A2(new_n387_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n377_), .A2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n324_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n308_), .A2(KEYINPUT32), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n394_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n395_), .B1(new_n303_), .B2(new_n394_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n253_), .B1(new_n376_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT33), .ZN(new_n398_));
  INV_X1    g197(.A(new_n360_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n399_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n398_), .B1(new_n400_), .B2(new_n365_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n315_), .A2(new_n318_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n359_), .A2(new_n353_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n403_), .B1(new_n369_), .B2(new_n353_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n402_), .B1(new_n404_), .B2(new_n365_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n373_), .A2(KEYINPUT33), .A3(new_n374_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n401_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT96), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT96), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n401_), .A2(new_n405_), .A3(new_n409_), .A4(new_n406_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n397_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n320_), .A2(new_n375_), .A3(new_n372_), .A4(new_n366_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n390_), .B1(new_n412_), .B2(new_n253_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT99), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT99), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n411_), .A2(new_n416_), .A3(new_n413_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n392_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G99gat), .A2(G106gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT6), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT66), .ZN(new_n421_));
  XOR2_X1   g220(.A(G85gat), .B(G92gat), .Z(new_n422_));
  AOI21_X1  g221(.A(new_n421_), .B1(KEYINPUT9), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(G92gat), .ZN(new_n424_));
  OR3_X1    g223(.A1(new_n362_), .A2(new_n424_), .A3(KEYINPUT9), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT10), .B(G99gat), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n426_), .A2(G106gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT65), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n423_), .A2(new_n425_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(G99gat), .ZN(new_n430_));
  INV_X1    g229(.A(G106gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT7), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n422_), .B1(new_n421_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT8), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n420_), .ZN(new_n437_));
  OAI211_X1 g236(.A(KEYINPUT8), .B(new_n422_), .C1(new_n433_), .C2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n429_), .A2(new_n436_), .A3(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G57gat), .B(G64gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT11), .ZN(new_n441_));
  XOR2_X1   g240(.A(new_n441_), .B(KEYINPUT67), .Z(new_n442_));
  NAND2_X1  g241(.A1(G71gat), .A2(G78gat), .ZN(new_n443_));
  INV_X1    g242(.A(G71gat), .ZN(new_n444_));
  INV_X1    g243(.A(G78gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n443_), .B(new_n446_), .C1(new_n440_), .C2(KEYINPUT11), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n442_), .B(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n439_), .A2(new_n449_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n448_), .A2(new_n429_), .A3(new_n436_), .A4(new_n438_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G230gat), .A2(G233gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT64), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT68), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n450_), .A2(KEYINPUT12), .A3(new_n451_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT12), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n439_), .A2(new_n458_), .A3(new_n449_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n454_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n456_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  AOI211_X1 g261(.A(KEYINPUT68), .B(new_n454_), .C1(new_n457_), .C2(new_n459_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n455_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G120gat), .B(G148gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(G204gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT5), .B(G176gat), .ZN(new_n467_));
  XOR2_X1   g266(.A(new_n466_), .B(new_n467_), .Z(new_n468_));
  NAND2_X1  g267(.A1(new_n464_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n468_), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n455_), .B(new_n470_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT13), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n469_), .A2(KEYINPUT13), .A3(new_n471_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n418_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G15gat), .B(G22gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G1gat), .A2(G8gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT14), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G1gat), .B(G8gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G231gat), .A2(G233gat), .ZN(new_n484_));
  XOR2_X1   g283(.A(new_n484_), .B(KEYINPUT73), .Z(new_n485_));
  XNOR2_X1  g284(.A(new_n483_), .B(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n448_), .B(new_n486_), .Z(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT74), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G127gat), .B(G155gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(G211gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(KEYINPUT16), .B(G183gat), .Z(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT17), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(new_n488_), .B(new_n494_), .Z(new_n495_));
  INV_X1    g294(.A(new_n487_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n496_), .A2(new_n493_), .A3(new_n492_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n498_), .B(KEYINPUT75), .Z(new_n499_));
  INV_X1    g298(.A(KEYINPUT37), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G29gat), .B(G36gat), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G43gat), .B(G50gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n503_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n501_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT15), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n439_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G232gat), .A2(G233gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT35), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n510_), .B(new_n515_), .C1(new_n439_), .C2(new_n507_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n513_), .A2(new_n514_), .ZN(new_n517_));
  XOR2_X1   g316(.A(new_n516_), .B(new_n517_), .Z(new_n518_));
  XNOR2_X1  g317(.A(G190gat), .B(G218gat), .ZN(new_n519_));
  INV_X1    g318(.A(G162gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT70), .B(G134gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n518_), .B1(KEYINPUT36), .B2(new_n524_), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n524_), .A2(KEYINPUT36), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT72), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n500_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  XOR2_X1   g328(.A(new_n526_), .B(KEYINPUT71), .Z(new_n530_));
  NAND2_X1  g329(.A1(new_n518_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n527_), .A2(new_n531_), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n529_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n529_), .A2(new_n532_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n499_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n509_), .A2(new_n483_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT77), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n483_), .A2(new_n507_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G229gat), .A2(G233gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n483_), .B(new_n507_), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n543_), .B(KEYINPUT76), .Z(new_n544_));
  NAND3_X1  g343(.A1(new_n544_), .A2(G229gat), .A3(G233gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G113gat), .B(G141gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G169gat), .B(G197gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n546_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n549_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n542_), .A2(new_n545_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT78), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n477_), .A2(new_n535_), .A3(new_n555_), .ZN(new_n556_));
  NOR3_X1   g355(.A1(new_n556_), .A2(G1gat), .A3(new_n377_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n557_), .A2(KEYINPUT38), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n558_), .B(KEYINPUT104), .Z(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(KEYINPUT38), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT101), .ZN(new_n561_));
  INV_X1    g360(.A(new_n553_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n476_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT102), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n564_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(new_n498_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT103), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n532_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n418_), .A2(new_n571_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n566_), .A2(KEYINPUT103), .A3(new_n498_), .A4(new_n567_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n570_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(G1gat), .B1(new_n574_), .B2(new_n377_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n559_), .A2(new_n561_), .A3(new_n575_), .ZN(G1324gat));
  OR2_X1    g375(.A1(new_n322_), .A2(new_n323_), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n556_), .A2(G8gat), .A3(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(G8gat), .B1(new_n574_), .B2(new_n577_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n579_), .A2(KEYINPUT39), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(KEYINPUT39), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n578_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n582_), .B(new_n583_), .Z(G1325gat));
  INV_X1    g383(.A(new_n390_), .ZN(new_n585_));
  OAI21_X1  g384(.A(G15gat), .B1(new_n574_), .B2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT41), .ZN(new_n587_));
  NOR3_X1   g386(.A1(new_n556_), .A2(G15gat), .A3(new_n585_), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n587_), .A2(new_n588_), .ZN(G1326gat));
  OAI21_X1  g388(.A(G22gat), .B1(new_n574_), .B2(new_n254_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT42), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n254_), .A2(G22gat), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n591_), .B1(new_n556_), .B2(new_n592_), .ZN(G1327gat));
  INV_X1    g392(.A(KEYINPUT109), .ZN(new_n594_));
  XOR2_X1   g393(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n595_));
  NAND2_X1  g394(.A1(new_n533_), .A2(new_n534_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n595_), .B1(new_n418_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT107), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  OR3_X1    g398(.A1(new_n418_), .A2(KEYINPUT43), .A3(new_n596_), .ZN(new_n600_));
  OAI211_X1 g399(.A(KEYINPUT107), .B(new_n595_), .C1(new_n418_), .C2(new_n596_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n599_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT108), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT44), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n499_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n566_), .A2(new_n567_), .ZN(new_n608_));
  AOI211_X1 g407(.A(new_n607_), .B(new_n608_), .C1(new_n603_), .C2(new_n604_), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n602_), .A2(new_n606_), .A3(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n606_), .B1(new_n602_), .B2(new_n609_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n376_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(G29gat), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n477_), .A2(new_n499_), .A3(new_n555_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n614_), .A2(new_n532_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NOR3_X1   g415(.A1(new_n616_), .A2(G29gat), .A3(new_n377_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n594_), .B1(new_n613_), .B2(new_n618_), .ZN(new_n619_));
  AOI211_X1 g418(.A(KEYINPUT109), .B(new_n617_), .C1(new_n612_), .C2(G29gat), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(G1328gat));
  INV_X1    g420(.A(KEYINPUT46), .ZN(new_n622_));
  INV_X1    g421(.A(G36gat), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n602_), .A2(new_n609_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(new_n605_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n602_), .A2(new_n606_), .A3(new_n609_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n577_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n623_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n615_), .A2(new_n623_), .A3(new_n628_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT45), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n622_), .B1(new_n629_), .B2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n630_), .B(KEYINPUT45), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n577_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n634_), .B(KEYINPUT46), .C1(new_n635_), .C2(new_n623_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n633_), .A2(new_n636_), .ZN(G1329gat));
  INV_X1    g436(.A(G43gat), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n615_), .A2(new_n638_), .A3(new_n390_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n585_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n639_), .B1(new_n640_), .B2(new_n638_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT47), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OAI211_X1 g442(.A(KEYINPUT47), .B(new_n639_), .C1(new_n640_), .C2(new_n638_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(G1330gat));
  INV_X1    g444(.A(G50gat), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n615_), .A2(new_n646_), .A3(new_n253_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n254_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n647_), .B1(new_n648_), .B2(new_n646_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT110), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT110), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n651_), .B(new_n647_), .C1(new_n648_), .C2(new_n646_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(G1331gat));
  NAND4_X1  g452(.A1(new_n572_), .A2(new_n607_), .A3(new_n554_), .A4(new_n476_), .ZN(new_n654_));
  INV_X1    g453(.A(G57gat), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n654_), .A2(new_n655_), .A3(new_n377_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n418_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n476_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n658_), .A2(new_n553_), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n657_), .A2(new_n535_), .A3(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(G57gat), .B1(new_n660_), .B2(new_n376_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n656_), .A2(new_n661_), .ZN(G1332gat));
  OAI21_X1  g461(.A(G64gat), .B1(new_n654_), .B2(new_n577_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT48), .ZN(new_n664_));
  INV_X1    g463(.A(G64gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n660_), .A2(new_n665_), .A3(new_n628_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(G1333gat));
  OAI21_X1  g466(.A(G71gat), .B1(new_n654_), .B2(new_n585_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT111), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT49), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n390_), .A2(new_n444_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT112), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n660_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n670_), .A2(new_n673_), .ZN(G1334gat));
  OAI21_X1  g473(.A(G78gat), .B1(new_n654_), .B2(new_n254_), .ZN(new_n675_));
  XOR2_X1   g474(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n676_));
  XNOR2_X1  g475(.A(new_n675_), .B(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n660_), .A2(new_n445_), .A3(new_n253_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1335gat));
  NAND2_X1  g478(.A1(new_n659_), .A2(new_n499_), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n418_), .A2(new_n532_), .A3(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(G85gat), .B1(new_n681_), .B2(new_n376_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n680_), .B(KEYINPUT115), .Z(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT114), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n602_), .A2(new_n685_), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n599_), .A2(KEYINPUT114), .A3(new_n600_), .A4(new_n601_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n684_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n377_), .A2(new_n362_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n682_), .B1(new_n688_), .B2(new_n689_), .ZN(G1336gat));
  AOI21_X1  g489(.A(G92gat), .B1(new_n681_), .B2(new_n628_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n577_), .A2(new_n424_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n691_), .B1(new_n688_), .B2(new_n692_), .ZN(G1337gat));
  XNOR2_X1  g492(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n694_));
  INV_X1    g493(.A(new_n681_), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n695_), .A2(new_n426_), .A3(new_n585_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n688_), .A2(new_n390_), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n694_), .B(new_n697_), .C1(new_n698_), .C2(new_n430_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n694_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n430_), .B1(new_n688_), .B2(new_n390_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n700_), .B1(new_n701_), .B2(new_n696_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n699_), .A2(new_n702_), .ZN(G1338gat));
  NAND3_X1  g502(.A1(new_n681_), .A2(new_n431_), .A3(new_n253_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n602_), .A2(new_n253_), .A3(new_n683_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT52), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n705_), .A2(new_n706_), .A3(G106gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n705_), .B2(G106gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n704_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT53), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT53), .ZN(new_n711_));
  OAI211_X1 g510(.A(new_n711_), .B(new_n704_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(G1339gat));
  NOR2_X1   g512(.A1(new_n324_), .A2(new_n585_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT55), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n715_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT118), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n457_), .A2(new_n454_), .A3(new_n459_), .ZN(new_n719_));
  OAI211_X1 g518(.A(KEYINPUT118), .B(new_n715_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n460_), .A2(KEYINPUT55), .A3(new_n461_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n718_), .A2(new_n719_), .A3(new_n720_), .A4(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(new_n468_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT56), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT120), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n722_), .A2(KEYINPUT56), .A3(new_n468_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n725_), .A2(new_n726_), .A3(new_n727_), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n722_), .A2(KEYINPUT120), .A3(KEYINPUT56), .A4(new_n468_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n551_), .B1(new_n544_), .B2(new_n541_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT119), .ZN(new_n731_));
  INV_X1    g530(.A(new_n540_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n541_), .B2(new_n732_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n733_), .A2(new_n552_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n729_), .A2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n728_), .A2(new_n735_), .A3(new_n471_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT58), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n728_), .A2(new_n735_), .A3(KEYINPUT58), .A4(new_n471_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n738_), .A2(new_n533_), .A3(new_n534_), .A4(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n553_), .A2(new_n471_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT117), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n742_), .B1(new_n725_), .B2(new_n727_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n734_), .A2(new_n472_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n532_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT57), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT57), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n747_), .B(new_n532_), .C1(new_n743_), .C2(new_n744_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n498_), .B1(new_n740_), .B2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n535_), .A2(new_n554_), .A3(new_n658_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT54), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n751_), .B(new_n752_), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n376_), .B(new_n714_), .C1(new_n750_), .C2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(G113gat), .B1(new_n755_), .B2(new_n553_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n607_), .B1(new_n740_), .B2(new_n749_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n757_), .A2(new_n753_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT59), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n714_), .A2(new_n759_), .A3(new_n376_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n758_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n754_), .A2(KEYINPUT121), .A3(KEYINPUT59), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT121), .B1(new_n754_), .B2(KEYINPUT59), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n762_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n555_), .A2(G113gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n756_), .B1(new_n766_), .B2(new_n767_), .ZN(G1340gat));
  OAI21_X1  g567(.A(G120gat), .B1(new_n765_), .B2(new_n658_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT60), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n770_), .B1(new_n658_), .B2(G120gat), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n755_), .B(new_n771_), .C1(new_n770_), .C2(G120gat), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n769_), .A2(new_n772_), .ZN(G1341gat));
  AOI21_X1  g572(.A(G127gat), .B1(new_n755_), .B2(new_n607_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n498_), .ZN(new_n775_));
  XOR2_X1   g574(.A(KEYINPUT122), .B(G127gat), .Z(new_n776_));
  NOR2_X1   g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n774_), .B1(new_n766_), .B2(new_n777_), .ZN(G1342gat));
  AOI21_X1  g577(.A(G134gat), .B1(new_n755_), .B2(new_n571_), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n533_), .A2(G134gat), .A3(new_n534_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n766_), .B2(new_n780_), .ZN(G1343gat));
  OR2_X1    g580(.A1(new_n750_), .A2(new_n753_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n782_), .A2(new_n376_), .A3(new_n577_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n254_), .A2(new_n390_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n783_), .A2(new_n562_), .A3(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(new_n202_), .ZN(G1344gat));
  NOR3_X1   g586(.A1(new_n783_), .A2(new_n658_), .A3(new_n785_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(new_n203_), .ZN(G1345gat));
  NOR3_X1   g588(.A1(new_n783_), .A2(new_n499_), .A3(new_n785_), .ZN(new_n790_));
  XOR2_X1   g589(.A(KEYINPUT61), .B(G155gat), .Z(new_n791_));
  XNOR2_X1  g590(.A(new_n790_), .B(new_n791_), .ZN(G1346gat));
  NOR2_X1   g591(.A1(new_n783_), .A2(new_n785_), .ZN(new_n793_));
  AOI21_X1  g592(.A(G162gat), .B1(new_n793_), .B2(new_n571_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n596_), .A2(new_n520_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n793_), .B2(new_n795_), .ZN(G1347gat));
  NOR3_X1   g595(.A1(new_n577_), .A2(new_n253_), .A3(new_n391_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n553_), .B(new_n797_), .C1(new_n757_), .C2(new_n753_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(G169gat), .ZN(new_n799_));
  INV_X1    g598(.A(new_n283_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n799_), .B1(new_n800_), .B2(new_n798_), .ZN(new_n801_));
  MUX2_X1   g600(.A(new_n799_), .B(new_n801_), .S(KEYINPUT62), .Z(G1348gat));
  NAND2_X1  g601(.A1(new_n782_), .A2(new_n797_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n804_), .A2(G176gat), .A3(new_n476_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT123), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n797_), .B1(new_n757_), .B2(new_n753_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n264_), .B1(new_n808_), .B2(new_n658_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n804_), .A2(KEYINPUT123), .A3(G176gat), .A4(new_n476_), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n807_), .A2(new_n809_), .A3(new_n810_), .ZN(G1349gat));
  OAI21_X1  g610(.A(new_n257_), .B1(new_n803_), .B2(new_n499_), .ZN(new_n812_));
  OR3_X1    g611(.A1(new_n808_), .A2(new_n775_), .A3(new_n272_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT124), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT124), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n812_), .A2(new_n816_), .A3(new_n813_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(G1350gat));
  OAI21_X1  g617(.A(G190gat), .B1(new_n808_), .B2(new_n596_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n571_), .A2(new_n273_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n819_), .B1(new_n808_), .B2(new_n820_), .ZN(new_n821_));
  XOR2_X1   g620(.A(new_n821_), .B(KEYINPUT125), .Z(G1351gat));
  NOR3_X1   g621(.A1(new_n785_), .A2(KEYINPUT126), .A3(new_n376_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n823_), .A2(new_n577_), .ZN(new_n824_));
  OAI21_X1  g623(.A(KEYINPUT126), .B1(new_n785_), .B2(new_n376_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n824_), .B(new_n825_), .C1(new_n750_), .C2(new_n753_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n826_), .A2(new_n562_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(new_n232_), .ZN(G1352gat));
  INV_X1    g627(.A(new_n826_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n829_), .A2(new_n476_), .A3(new_n231_), .ZN(new_n830_));
  OAI21_X1  g629(.A(G204gat), .B1(new_n826_), .B2(new_n658_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT127), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n832_), .B(new_n833_), .ZN(G1353gat));
  NOR2_X1   g633(.A1(new_n826_), .A2(new_n775_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n836_));
  AND2_X1   g635(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n835_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n835_), .B2(new_n836_), .ZN(G1354gat));
  INV_X1    g638(.A(G218gat), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n826_), .A2(new_n840_), .A3(new_n596_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n829_), .A2(new_n571_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n841_), .B1(new_n840_), .B2(new_n842_), .ZN(G1355gat));
endmodule


