//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 1 0 1 1 1 1 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n667_, new_n668_, new_n669_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n820_,
    new_n821_, new_n822_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n832_, new_n833_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n869_, new_n870_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_;
  NOR2_X1   g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(KEYINPUT1), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(KEYINPUT1), .ZN(new_n205_));
  AOI211_X1 g004(.A(new_n202_), .B(new_n204_), .C1(KEYINPUT86), .C2(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n206_), .B1(KEYINPUT86), .B2(new_n205_), .ZN(new_n207_));
  OR2_X1    g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT2), .ZN(new_n209_));
  XOR2_X1   g008(.A(G155gat), .B(G162gat), .Z(new_n210_));
  AOI22_X1  g009(.A1(new_n207_), .A2(new_n208_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT85), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT3), .B1(new_n208_), .B2(KEYINPUT87), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n215_), .B1(new_n209_), .B2(new_n212_), .ZN(new_n216_));
  NOR3_X1   g015(.A1(new_n208_), .A2(KEYINPUT87), .A3(KEYINPUT3), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n210_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G127gat), .B(G134gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G113gat), .B(G120gat), .ZN(new_n220_));
  XOR2_X1   g019(.A(new_n219_), .B(new_n220_), .Z(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(KEYINPUT96), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n214_), .A2(new_n218_), .A3(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT97), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n214_), .A2(new_n218_), .ZN(new_n226_));
  XOR2_X1   g025(.A(new_n221_), .B(KEYINPUT83), .Z(new_n227_));
  AOI21_X1  g026(.A(KEYINPUT97), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n225_), .B(KEYINPUT4), .C1(new_n228_), .C2(new_n223_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G225gat), .A2(G233gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT4), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n226_), .A2(new_n231_), .A3(new_n227_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n229_), .A2(new_n230_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n230_), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n225_), .B(new_n234_), .C1(new_n228_), .C2(new_n223_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT99), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G1gat), .B(G29gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT0), .ZN(new_n238_));
  INV_X1    g037(.A(G57gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(G85gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n235_), .A2(new_n236_), .A3(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n236_), .B1(new_n235_), .B2(new_n242_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n233_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n242_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n230_), .B1(new_n229_), .B2(new_n232_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n225_), .B1(new_n228_), .B2(new_n223_), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n248_), .A2(new_n230_), .ZN(new_n249_));
  OAI211_X1 g048(.A(KEYINPUT33), .B(new_n246_), .C1(new_n247_), .C2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT25), .B(G183gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT26), .B(G190gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT82), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G183gat), .A2(G190gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT23), .ZN(new_n256_));
  OR2_X1    g055(.A1(G169gat), .A2(G176gat), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n257_), .A2(KEYINPUT24), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G169gat), .A2(G176gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n257_), .A2(KEYINPUT24), .A3(new_n259_), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n256_), .A2(new_n258_), .A3(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n254_), .A2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n256_), .B1(G183gat), .B2(G190gat), .ZN(new_n263_));
  XOR2_X1   g062(.A(KEYINPUT22), .B(G169gat), .Z(new_n264_));
  OAI211_X1 g063(.A(new_n263_), .B(new_n259_), .C1(G176gat), .C2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G211gat), .B(G218gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT91), .ZN(new_n268_));
  INV_X1    g067(.A(G197gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(G204gat), .ZN(new_n270_));
  INV_X1    g069(.A(G204gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(G197gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT21), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n268_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n270_), .A2(KEYINPUT89), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(new_n272_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n270_), .A2(KEYINPUT89), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT21), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(KEYINPUT90), .B(KEYINPUT21), .Z(new_n280_));
  OAI211_X1 g079(.A(new_n268_), .B(new_n279_), .C1(new_n273_), .C2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n275_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n266_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT95), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n258_), .A2(new_n260_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n253_), .A2(new_n256_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n265_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT20), .B1(new_n282_), .B2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n285_), .A2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G226gat), .A2(G233gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n290_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n282_), .A2(new_n288_), .ZN(new_n295_));
  OAI211_X1 g094(.A(new_n295_), .B(KEYINPUT20), .C1(new_n282_), .C2(new_n266_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n293_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G8gat), .B(G36gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT18), .ZN(new_n300_));
  XOR2_X1   g099(.A(G64gat), .B(G92gat), .Z(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  AND3_X1   g101(.A1(new_n294_), .A2(new_n298_), .A3(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n302_), .B1(new_n294_), .B2(new_n298_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n245_), .A2(new_n250_), .A3(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n246_), .B1(new_n247_), .B2(new_n249_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT33), .ZN(new_n308_));
  AND3_X1   g107(.A1(new_n307_), .A2(KEYINPUT98), .A3(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(KEYINPUT98), .B1(new_n307_), .B2(new_n308_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n306_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n248_), .A2(new_n230_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n229_), .A2(new_n232_), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n242_), .B(new_n312_), .C1(new_n313_), .C2(new_n230_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(new_n307_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n290_), .A2(new_n297_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n296_), .A2(new_n293_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT100), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n302_), .A2(KEYINPUT32), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n318_), .A2(new_n319_), .A3(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n316_), .A2(new_n321_), .A3(new_n317_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT100), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n294_), .A2(new_n298_), .ZN(new_n325_));
  AOI22_X1  g124(.A1(new_n322_), .A2(new_n324_), .B1(new_n325_), .B2(new_n320_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n315_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT101), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT101), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n315_), .A2(new_n326_), .A3(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n311_), .A2(new_n328_), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n282_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n332_), .B1(new_n226_), .B2(KEYINPUT29), .ZN(new_n333_));
  AOI22_X1  g132(.A1(new_n282_), .A2(KEYINPUT88), .B1(G228gat), .B2(G233gat), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  AOI211_X1 g135(.A(new_n332_), .B(new_n334_), .C1(new_n226_), .C2(KEYINPUT29), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G78gat), .B(G106gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n336_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(KEYINPUT92), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n333_), .A2(new_n335_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n341_), .B1(new_n342_), .B2(new_n337_), .ZN(new_n343_));
  OR3_X1    g142(.A1(new_n226_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT28), .B1(new_n226_), .B2(KEYINPUT29), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  XOR2_X1   g145(.A(G22gat), .B(G50gat), .Z(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n347_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n344_), .A2(new_n345_), .A3(new_n349_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n340_), .A2(new_n343_), .A3(new_n348_), .A4(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n341_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n336_), .A2(new_n338_), .A3(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(new_n343_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n348_), .A2(new_n350_), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n354_), .A2(KEYINPUT93), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT93), .B1(new_n354_), .B2(new_n355_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n351_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n266_), .B(KEYINPUT30), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G71gat), .B(G99gat), .ZN(new_n360_));
  INV_X1    g159(.A(G43gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G227gat), .A2(G233gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(G15gat), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n362_), .B(new_n364_), .Z(new_n365_));
  XNOR2_X1  g164(.A(new_n359_), .B(new_n365_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n366_), .A2(KEYINPUT84), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(KEYINPUT84), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n227_), .B(KEYINPUT31), .Z(new_n369_));
  OR3_X1    g168(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n366_), .A2(KEYINPUT84), .A3(new_n369_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n358_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n331_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n372_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n358_), .A2(new_n375_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n372_), .B(new_n351_), .C1(new_n356_), .C2(new_n357_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT27), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n303_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n318_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n380_), .B1(new_n302_), .B2(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n379_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n315_), .A2(KEYINPUT102), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT102), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n314_), .A2(new_n386_), .A3(new_n307_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n384_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n378_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n374_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G232gat), .A2(G233gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT34), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT76), .B1(new_n392_), .B2(KEYINPUT35), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT7), .ZN(new_n394_));
  INV_X1    g193(.A(G99gat), .ZN(new_n395_));
  INV_X1    g194(.A(G106gat), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G99gat), .A2(G106gat), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT6), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n397_), .A2(new_n400_), .A3(new_n401_), .A4(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(G92gat), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n241_), .A2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(G85gat), .A2(G92gat), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n403_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n403_), .A2(new_n407_), .A3(new_n409_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  XOR2_X1   g213(.A(KEYINPUT10), .B(G99gat), .Z(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n396_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n241_), .A2(KEYINPUT64), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT64), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(G85gat), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n404_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT65), .B1(new_n421_), .B2(KEYINPUT9), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT65), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT9), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT64), .B(G85gat), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n423_), .B(new_n424_), .C1(new_n425_), .C2(new_n404_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n422_), .A2(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n406_), .B1(new_n405_), .B2(KEYINPUT9), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n417_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n414_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G29gat), .B(G36gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT74), .ZN(new_n432_));
  XOR2_X1   g231(.A(G43gat), .B(G50gat), .Z(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n432_), .B(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n393_), .B1(new_n430_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT69), .ZN(new_n437_));
  AND3_X1   g236(.A1(new_n403_), .A2(new_n407_), .A3(new_n409_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n409_), .B1(new_n403_), .B2(new_n407_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n437_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n411_), .A2(KEYINPUT69), .A3(new_n412_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n428_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n442_), .B1(new_n422_), .B2(new_n426_), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n440_), .B(new_n441_), .C1(new_n443_), .C2(new_n417_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT70), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n429_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n447_), .A2(KEYINPUT70), .A3(new_n441_), .A4(new_n440_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n432_), .B(new_n433_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT15), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT15), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n435_), .A2(new_n452_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n449_), .A2(new_n454_), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n455_), .A2(KEYINPUT75), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n455_), .A2(KEYINPUT75), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n436_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n392_), .A2(KEYINPUT35), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(G190gat), .B(G218gat), .Z(new_n462_));
  XNOR2_X1  g261(.A(G134gat), .B(G162gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n465_), .A2(KEYINPUT36), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n459_), .B(new_n436_), .C1(new_n456_), .C2(new_n457_), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n461_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n464_), .B(KEYINPUT36), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n470_), .B1(new_n461_), .B2(new_n467_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n468_), .A2(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(G127gat), .B(G155gat), .Z(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT16), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G183gat), .B(G211gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT17), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT79), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT14), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT77), .B(G8gat), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n480_), .B1(new_n481_), .B2(G1gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT78), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G15gat), .B(G22gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(G1gat), .B(G8gat), .Z(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n486_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n483_), .A2(new_n484_), .A3(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  OR2_X1    g289(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n491_));
  INV_X1    g290(.A(G78gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  AND2_X1   g293(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n495_));
  NOR2_X1   g294(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n496_));
  OAI21_X1  g295(.A(G78gat), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G57gat), .B(G64gat), .ZN(new_n498_));
  AOI22_X1  g297(.A1(new_n494_), .A2(new_n497_), .B1(new_n498_), .B2(KEYINPUT11), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n494_), .A2(new_n497_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n498_), .A2(KEYINPUT11), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT11), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n239_), .A2(G64gat), .ZN(new_n504_));
  INV_X1    g303(.A(G64gat), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n505_), .A2(G57gat), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n503_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n502_), .A2(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n499_), .B1(new_n501_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G231gat), .A2(G233gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n490_), .B(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n479_), .A2(new_n512_), .ZN(new_n513_));
  OR2_X1    g312(.A1(new_n513_), .A2(KEYINPUT80), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(KEYINPUT80), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n476_), .A2(new_n477_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n512_), .A2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n514_), .A2(new_n515_), .A3(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n472_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n509_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT12), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n520_), .B1(new_n414_), .B2(new_n429_), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n413_), .B(new_n509_), .C1(new_n443_), .C2(new_n417_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT12), .ZN(new_n525_));
  AOI22_X1  g324(.A1(new_n449_), .A2(new_n522_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G230gat), .A2(G233gat), .ZN(new_n527_));
  AOI21_X1  g326(.A(KEYINPUT71), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n521_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n525_), .A2(new_n523_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT71), .ZN(new_n531_));
  INV_X1    g330(.A(new_n527_), .ZN(new_n532_));
  NOR4_X1   g331(.A1(new_n529_), .A2(new_n530_), .A3(new_n531_), .A4(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n528_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT73), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT68), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n523_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(new_n524_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n523_), .A2(new_n536_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n532_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(G120gat), .B(G148gat), .Z(new_n541_));
  XNOR2_X1  g340(.A(G176gat), .B(G204gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n543_), .B(new_n544_), .Z(new_n545_));
  NAND4_X1  g344(.A1(new_n534_), .A2(new_n535_), .A3(new_n540_), .A4(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(KEYINPUT69), .B1(new_n411_), .B2(new_n412_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n429_), .A2(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(KEYINPUT70), .B1(new_n548_), .B2(new_n441_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n444_), .A2(new_n445_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n522_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n525_), .A2(new_n523_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(new_n527_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(new_n531_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n526_), .A2(KEYINPUT71), .A3(new_n527_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n554_), .A2(new_n540_), .A3(new_n555_), .A4(new_n545_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT73), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n546_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n534_), .A2(new_n540_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n545_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n558_), .A2(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT13), .Z(new_n563_));
  NAND2_X1  g362(.A1(G229gat), .A2(G233gat), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n450_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n451_), .A2(new_n453_), .A3(new_n487_), .A4(new_n489_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n565_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n490_), .A2(new_n435_), .ZN(new_n571_));
  OR3_X1    g370(.A1(new_n571_), .A2(new_n564_), .A3(new_n566_), .ZN(new_n572_));
  XOR2_X1   g371(.A(G113gat), .B(G141gat), .Z(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT81), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G169gat), .B(G197gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n570_), .A2(new_n572_), .A3(new_n577_), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n571_), .A2(new_n564_), .A3(new_n566_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n576_), .B1(new_n579_), .B2(new_n569_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n563_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n390_), .A2(new_n519_), .A3(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n385_), .A2(new_n387_), .ZN(new_n584_));
  OAI21_X1  g383(.A(G1gat), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  AOI22_X1  g384(.A1(new_n331_), .A2(new_n373_), .B1(new_n378_), .B2(new_n388_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n582_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n472_), .A2(KEYINPUT37), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n461_), .A2(new_n467_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(new_n469_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n461_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT37), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n589_), .A2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n596_), .A2(new_n518_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n588_), .A2(new_n597_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n598_), .A2(G1gat), .A3(new_n584_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT38), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n599_), .A2(new_n600_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n585_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT103), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(G1324gat));
  INV_X1    g404(.A(new_n384_), .ZN(new_n606_));
  OR3_X1    g405(.A1(new_n598_), .A2(new_n481_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(G8gat), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n583_), .A2(new_n606_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n608_), .B1(new_n609_), .B2(KEYINPUT104), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT104), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n612_), .B1(new_n583_), .B2(new_n606_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n610_), .A2(new_n611_), .A3(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n611_), .B1(new_n610_), .B2(new_n613_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n607_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT40), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  OAI211_X1 g417(.A(KEYINPUT40), .B(new_n607_), .C1(new_n614_), .C2(new_n615_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(G1325gat));
  INV_X1    g419(.A(G15gat), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n372_), .A2(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n598_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n583_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n621_), .B1(new_n624_), .B2(new_n372_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT41), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n623_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n627_), .B1(new_n626_), .B2(new_n625_), .ZN(G1326gat));
  INV_X1    g427(.A(new_n358_), .ZN(new_n629_));
  OAI21_X1  g428(.A(G22gat), .B1(new_n583_), .B2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT42), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n629_), .A2(G22gat), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n631_), .B1(new_n598_), .B2(new_n632_), .ZN(G1327gat));
  INV_X1    g432(.A(new_n518_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n593_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n588_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n584_), .ZN(new_n638_));
  AOI21_X1  g437(.A(G29gat), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  XOR2_X1   g438(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n640_));
  INV_X1    g439(.A(KEYINPUT43), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n390_), .A2(new_n641_), .A3(new_n596_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n468_), .A2(new_n471_), .A3(new_n594_), .ZN(new_n643_));
  AOI21_X1  g442(.A(KEYINPUT37), .B1(new_n591_), .B2(new_n592_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(KEYINPUT43), .B1(new_n586_), .B2(new_n645_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n642_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n582_), .A2(new_n518_), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n648_), .A2(KEYINPUT105), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(KEYINPUT105), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n640_), .B1(new_n647_), .B2(new_n651_), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n652_), .A2(G29gat), .A3(new_n638_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n642_), .A2(new_n646_), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n654_), .A2(KEYINPUT44), .A3(new_n649_), .A4(new_n650_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n639_), .B1(new_n653_), .B2(new_n655_), .ZN(G1328gat));
  NAND3_X1  g455(.A1(new_n652_), .A2(new_n384_), .A3(new_n655_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(G36gat), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n636_), .A2(G36gat), .A3(new_n606_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT45), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n658_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT46), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n658_), .A2(new_n661_), .A3(KEYINPUT46), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1329gat));
  NAND4_X1  g465(.A1(new_n652_), .A2(G43gat), .A3(new_n372_), .A4(new_n655_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n361_), .B1(new_n636_), .B2(new_n375_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g469(.A1(new_n652_), .A2(new_n358_), .A3(new_n655_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(G50gat), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n629_), .A2(G50gat), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT107), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n672_), .B1(new_n636_), .B2(new_n674_), .ZN(G1331gat));
  INV_X1    g474(.A(new_n581_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n562_), .B(KEYINPUT13), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n586_), .A2(new_n676_), .A3(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(new_n519_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n679_), .A2(new_n239_), .A3(new_n584_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n597_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n584_), .B1(new_n681_), .B2(KEYINPUT108), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n682_), .B1(KEYINPUT108), .B2(new_n681_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n680_), .B1(new_n683_), .B2(new_n239_), .ZN(G1332gat));
  OAI21_X1  g483(.A(G64gat), .B1(new_n679_), .B2(new_n606_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT48), .ZN(new_n686_));
  INV_X1    g485(.A(new_n681_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n687_), .A2(new_n505_), .A3(new_n384_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(G1333gat));
  OAI21_X1  g488(.A(G71gat), .B1(new_n679_), .B2(new_n375_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT49), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n375_), .A2(G71gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(new_n681_), .B2(new_n692_), .ZN(G1334gat));
  OAI21_X1  g492(.A(G78gat), .B1(new_n679_), .B2(new_n629_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT50), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n687_), .A2(new_n492_), .A3(new_n358_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1335gat));
  INV_X1    g496(.A(KEYINPUT109), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n654_), .A2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n642_), .A2(new_n646_), .A3(KEYINPUT109), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n677_), .A2(new_n676_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(new_n518_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n699_), .A2(new_n700_), .A3(new_n703_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n704_), .A2(new_n584_), .A3(new_n425_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n678_), .A2(new_n635_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G85gat), .B1(new_n706_), .B2(new_n638_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n705_), .A2(new_n707_), .ZN(G1336gat));
  OAI21_X1  g507(.A(G92gat), .B1(new_n704_), .B2(new_n606_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n706_), .A2(new_n404_), .A3(new_n384_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1337gat));
  NAND4_X1  g510(.A1(new_n699_), .A2(new_n372_), .A3(new_n700_), .A4(new_n703_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(G99gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n706_), .A2(new_n415_), .A3(new_n372_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT51), .ZN(G1338gat));
  NOR2_X1   g515(.A1(new_n629_), .A2(G106gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n678_), .A2(new_n635_), .A3(new_n717_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n718_), .A2(KEYINPUT110), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n718_), .A2(KEYINPUT110), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n702_), .A2(new_n629_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n396_), .B1(new_n654_), .B2(new_n721_), .ZN(new_n722_));
  OAI22_X1  g521(.A1(new_n719_), .A2(new_n720_), .B1(new_n722_), .B2(KEYINPUT52), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n722_), .A2(KEYINPUT52), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  XOR2_X1   g524(.A(KEYINPUT111), .B(KEYINPUT53), .Z(new_n726_));
  XNOR2_X1  g525(.A(new_n725_), .B(new_n726_), .ZN(G1339gat));
  OR4_X1    g526(.A1(KEYINPUT119), .A2(new_n584_), .A3(new_n377_), .A4(new_n384_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n638_), .A2(new_n606_), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT119), .B1(new_n729_), .B2(new_n377_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT59), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n728_), .A2(new_n730_), .A3(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT54), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n634_), .A2(KEYINPUT112), .A3(new_n581_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n735_), .B1(new_n518_), .B2(new_n676_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n677_), .A2(new_n733_), .A3(new_n737_), .A4(new_n645_), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n738_), .A2(KEYINPUT113), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(KEYINPUT113), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n677_), .A2(new_n645_), .A3(new_n737_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT54), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n739_), .A2(new_n740_), .A3(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n564_), .B1(new_n571_), .B2(new_n566_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n567_), .A2(new_n565_), .A3(new_n568_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(new_n745_), .A3(new_n577_), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n580_), .A2(KEYINPUT115), .A3(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(KEYINPUT115), .B1(new_n580_), .B2(new_n746_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n558_), .B2(new_n561_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n581_), .B1(new_n546_), .B2(new_n557_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT55), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n554_), .A2(new_n752_), .A3(new_n555_), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n551_), .A2(KEYINPUT55), .A3(new_n527_), .A4(new_n552_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n532_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n545_), .B1(new_n753_), .B2(new_n756_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n757_), .A2(KEYINPUT56), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT56), .ZN(new_n759_));
  AOI211_X1 g558(.A(new_n759_), .B(new_n545_), .C1(new_n753_), .C2(new_n756_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n751_), .B1(new_n758_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT114), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n750_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n751_), .B(KEYINPUT114), .C1(new_n758_), .C2(new_n760_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n472_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n753_), .A2(new_n756_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n768_), .A2(KEYINPUT56), .A3(new_n560_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT117), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n560_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n759_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n757_), .A2(new_n773_), .A3(KEYINPUT56), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n770_), .A2(new_n772_), .A3(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n749_), .B1(new_n557_), .B2(new_n546_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(KEYINPUT58), .A3(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n596_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT58), .B1(new_n775_), .B2(new_n776_), .ZN(new_n779_));
  OAI22_X1  g578(.A1(new_n765_), .A2(new_n767_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n761_), .A2(new_n762_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n750_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(new_n764_), .A3(new_n782_), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n783_), .A2(KEYINPUT57), .A3(new_n593_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n518_), .B1(new_n780_), .B2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n732_), .B1(new_n743_), .B2(new_n785_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n728_), .A2(new_n730_), .ZN(new_n787_));
  OAI21_X1  g586(.A(KEYINPUT118), .B1(new_n780_), .B2(new_n784_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n783_), .A2(new_n593_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n766_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n765_), .A2(KEYINPUT57), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT118), .ZN(new_n792_));
  INV_X1    g591(.A(new_n779_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n793_), .A2(new_n596_), .A3(new_n777_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n790_), .A2(new_n791_), .A3(new_n792_), .A4(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n634_), .B1(new_n788_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n743_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n787_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n786_), .B1(new_n798_), .B2(KEYINPUT59), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n799_), .A2(new_n676_), .ZN(new_n800_));
  INV_X1    g599(.A(G113gat), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n676_), .A2(new_n801_), .ZN(new_n802_));
  OAI22_X1  g601(.A1(new_n800_), .A2(new_n801_), .B1(new_n798_), .B2(new_n802_), .ZN(G1340gat));
  AND2_X1   g602(.A1(new_n799_), .A2(new_n563_), .ZN(new_n804_));
  INV_X1    g603(.A(G120gat), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n677_), .A2(KEYINPUT60), .A3(G120gat), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n806_), .B1(KEYINPUT60), .B2(G120gat), .ZN(new_n807_));
  OAI22_X1  g606(.A1(new_n804_), .A2(new_n805_), .B1(new_n798_), .B2(new_n807_), .ZN(G1341gat));
  INV_X1    g607(.A(G127gat), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n518_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n799_), .A2(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n798_), .A2(new_n518_), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n811_), .B(KEYINPUT120), .C1(G127gat), .C2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n812_), .A2(G127gat), .ZN(new_n815_));
  INV_X1    g614(.A(new_n810_), .ZN(new_n816_));
  AOI211_X1 g615(.A(new_n786_), .B(new_n816_), .C1(new_n798_), .C2(KEYINPUT59), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n814_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n813_), .A2(new_n818_), .ZN(G1342gat));
  AND2_X1   g618(.A1(new_n799_), .A2(new_n596_), .ZN(new_n820_));
  INV_X1    g619(.A(G134gat), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n472_), .A2(new_n821_), .ZN(new_n822_));
  OAI22_X1  g621(.A1(new_n820_), .A2(new_n821_), .B1(new_n798_), .B2(new_n822_), .ZN(G1343gat));
  NAND2_X1  g622(.A1(new_n788_), .A2(new_n795_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n518_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n743_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n376_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n826_), .A2(new_n638_), .A3(new_n827_), .A4(new_n606_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n828_), .A2(new_n581_), .ZN(new_n829_));
  INV_X1    g628(.A(G141gat), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n829_), .B(new_n830_), .ZN(G1344gat));
  NOR2_X1   g630(.A1(new_n828_), .A2(new_n677_), .ZN(new_n832_));
  XOR2_X1   g631(.A(KEYINPUT121), .B(G148gat), .Z(new_n833_));
  XNOR2_X1  g632(.A(new_n832_), .B(new_n833_), .ZN(G1345gat));
  NOR2_X1   g633(.A1(new_n828_), .A2(new_n518_), .ZN(new_n835_));
  XOR2_X1   g634(.A(KEYINPUT61), .B(G155gat), .Z(new_n836_));
  XNOR2_X1  g635(.A(new_n835_), .B(new_n836_), .ZN(G1346gat));
  OAI21_X1  g636(.A(G162gat), .B1(new_n828_), .B2(new_n645_), .ZN(new_n838_));
  OR2_X1    g637(.A1(new_n593_), .A2(G162gat), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n828_), .B2(new_n839_), .ZN(G1347gat));
  AND2_X1   g639(.A1(new_n743_), .A2(new_n785_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n638_), .A2(new_n375_), .A3(new_n606_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n629_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  OR3_X1    g644(.A1(new_n845_), .A2(new_n581_), .A3(new_n264_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n842_), .ZN(new_n847_));
  OR3_X1    g646(.A1(new_n847_), .A2(KEYINPUT122), .A3(new_n581_), .ZN(new_n848_));
  OAI21_X1  g647(.A(KEYINPUT122), .B1(new_n847_), .B2(new_n581_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n629_), .A3(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(G169gat), .B1(new_n850_), .B2(new_n841_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n851_), .A2(KEYINPUT123), .A3(KEYINPUT62), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n852_), .B1(KEYINPUT62), .B2(new_n851_), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT123), .B1(new_n851_), .B2(KEYINPUT62), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n846_), .B1(new_n853_), .B2(new_n854_), .ZN(G1348gat));
  AOI21_X1  g654(.A(G176gat), .B1(new_n844_), .B2(new_n563_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n358_), .B1(new_n825_), .B2(new_n743_), .ZN(new_n857_));
  OR2_X1    g656(.A1(new_n857_), .A2(KEYINPUT124), .ZN(new_n858_));
  OAI211_X1 g657(.A(KEYINPUT124), .B(new_n629_), .C1(new_n796_), .C2(new_n797_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n847_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n563_), .A2(G176gat), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n856_), .B1(new_n860_), .B2(new_n861_), .ZN(G1349gat));
  NOR3_X1   g661(.A1(new_n845_), .A2(new_n518_), .A3(new_n251_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n857_), .A2(KEYINPUT124), .ZN(new_n864_));
  INV_X1    g663(.A(new_n859_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n634_), .B(new_n842_), .C1(new_n864_), .C2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(G183gat), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n863_), .B1(new_n866_), .B2(new_n867_), .ZN(G1350gat));
  OAI21_X1  g667(.A(G190gat), .B1(new_n845_), .B2(new_n645_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n844_), .A2(new_n472_), .A3(new_n252_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1351gat));
  INV_X1    g670(.A(KEYINPUT125), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n638_), .A2(new_n606_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n826_), .A2(new_n872_), .A3(new_n827_), .A4(new_n873_), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n827_), .B(new_n873_), .C1(new_n796_), .C2(new_n797_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT125), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(G197gat), .B1(new_n877_), .B2(new_n676_), .ZN(new_n878_));
  AOI211_X1 g677(.A(new_n269_), .B(new_n581_), .C1(new_n874_), .C2(new_n876_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1352gat));
  AND2_X1   g679(.A1(new_n875_), .A2(KEYINPUT125), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n875_), .A2(KEYINPUT125), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n563_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(G204gat), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n877_), .A2(new_n271_), .A3(new_n563_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1353gat));
  NOR2_X1   g685(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(KEYINPUT126), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n518_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n888_), .B1(new_n877_), .B2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n889_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n888_), .ZN(new_n892_));
  AOI211_X1 g691(.A(new_n891_), .B(new_n892_), .C1(new_n874_), .C2(new_n876_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n890_), .A2(new_n893_), .ZN(G1354gat));
  NAND2_X1  g693(.A1(new_n877_), .A2(new_n472_), .ZN(new_n895_));
  XOR2_X1   g694(.A(KEYINPUT127), .B(G218gat), .Z(new_n896_));
  NOR2_X1   g695(.A1(new_n645_), .A2(new_n896_), .ZN(new_n897_));
  AOI22_X1  g696(.A1(new_n895_), .A2(new_n896_), .B1(new_n877_), .B2(new_n897_), .ZN(G1355gat));
endmodule


