//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 1 0 0 0 0 0 0 1 1 0 0 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n761_, new_n762_, new_n763_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n891_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n928_, new_n929_, new_n930_,
    new_n932_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_;
  INV_X1    g000(.A(KEYINPUT65), .ZN(new_n202_));
  OR3_X1    g001(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT6), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n205_), .B1(G99gat), .B2(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n207_), .A2(KEYINPUT6), .ZN(new_n208_));
  OAI211_X1 g007(.A(new_n203_), .B(new_n204_), .C1(new_n206_), .C2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT8), .ZN(new_n210_));
  INV_X1    g009(.A(G85gat), .ZN(new_n211_));
  INV_X1    g010(.A(G92gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n215_), .A2(KEYINPUT64), .ZN(new_n216_));
  AND3_X1   g015(.A1(new_n209_), .A2(new_n210_), .A3(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n210_), .B1(new_n209_), .B2(new_n216_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n202_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n209_), .A2(new_n216_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT8), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n209_), .A2(new_n210_), .A3(new_n216_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(KEYINPUT65), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n219_), .A2(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(KEYINPUT10), .B(G99gat), .Z(new_n225_));
  INV_X1    g024(.A(G106gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n206_), .A2(new_n208_), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n214_), .A2(KEYINPUT9), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n213_), .A2(KEYINPUT9), .A3(new_n214_), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .A4(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n224_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G57gat), .B(G64gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT11), .ZN(new_n234_));
  XOR2_X1   g033(.A(G71gat), .B(G78gat), .Z(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n233_), .A2(KEYINPUT11), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n234_), .A2(new_n235_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(KEYINPUT12), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n232_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n221_), .A2(new_n222_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n239_), .B1(new_n237_), .B2(new_n236_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(new_n231_), .A3(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT12), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n217_), .A2(new_n218_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n231_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n239_), .B(new_n238_), .C1(new_n247_), .C2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G230gat), .A2(G233gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n242_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n251_), .B1(new_n249_), .B2(new_n245_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G120gat), .B(G148gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT5), .ZN(new_n257_));
  XOR2_X1   g056(.A(G176gat), .B(G204gat), .Z(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n255_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT67), .ZN(new_n261_));
  AOI22_X1  g060(.A1(new_n232_), .A2(new_n241_), .B1(new_n246_), .B2(new_n249_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n253_), .B1(new_n262_), .B2(new_n251_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n259_), .B1(new_n263_), .B2(KEYINPUT66), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT66), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n255_), .A2(new_n265_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n260_), .B(new_n261_), .C1(new_n264_), .C2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT13), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n263_), .A2(KEYINPUT66), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n255_), .A2(new_n265_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n269_), .A2(new_n270_), .A3(KEYINPUT67), .A4(new_n259_), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n267_), .A2(new_n268_), .A3(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n268_), .B1(new_n267_), .B2(new_n271_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT72), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G29gat), .B(G36gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G43gat), .B(G50gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n278_), .A2(new_n279_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n277_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n278_), .A2(new_n279_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n284_), .A2(new_n276_), .A3(new_n280_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT15), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n283_), .A2(new_n285_), .A3(KEYINPUT15), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(new_n232_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n247_), .A2(new_n248_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n286_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G232gat), .A2(G233gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT35), .ZN(new_n296_));
  XOR2_X1   g095(.A(KEYINPUT68), .B(KEYINPUT34), .Z(new_n297_));
  XOR2_X1   g096(.A(new_n296_), .B(new_n297_), .Z(new_n298_));
  NAND4_X1  g097(.A1(new_n292_), .A2(KEYINPUT71), .A3(new_n294_), .A4(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(KEYINPUT35), .B1(new_n292_), .B2(new_n294_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n248_), .B1(new_n219_), .B2(new_n223_), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n294_), .B(KEYINPUT71), .C1(new_n301_), .C2(new_n290_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n298_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n275_), .B(new_n299_), .C1(new_n300_), .C2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G190gat), .B(G218gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G134gat), .B(G162gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n308_), .A2(KEYINPUT36), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n305_), .A2(new_n310_), .ZN(new_n311_));
  AOI22_X1  g110(.A1(new_n291_), .A2(new_n232_), .B1(new_n286_), .B2(new_n293_), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n302_), .B(new_n303_), .C1(new_n312_), .C2(KEYINPUT35), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n313_), .A2(new_n275_), .A3(new_n299_), .A4(new_n309_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n299_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(KEYINPUT36), .A3(new_n308_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT37), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n319_), .A2(KEYINPUT73), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(KEYINPUT73), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n318_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n315_), .A2(KEYINPUT73), .A3(new_n319_), .A4(new_n317_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G231gat), .A2(G233gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n244_), .B(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G1gat), .B(G8gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT74), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G15gat), .B(G22gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G1gat), .A2(G8gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT14), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n328_), .B(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n326_), .B(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(G127gat), .B(G155gat), .Z(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G183gat), .B(G211gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT17), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n340_), .A2(new_n341_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n335_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n344_), .B1(new_n342_), .B2(new_n335_), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n345_), .B(KEYINPUT76), .Z(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n274_), .A2(new_n323_), .A3(new_n324_), .A4(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G229gat), .A2(G233gat), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n328_), .B(new_n332_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(new_n286_), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n284_), .A2(new_n276_), .A3(new_n280_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n276_), .B1(new_n284_), .B2(new_n280_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n334_), .A2(new_n356_), .ZN(new_n357_));
  AND3_X1   g156(.A1(new_n353_), .A2(new_n357_), .A3(KEYINPUT77), .ZN(new_n358_));
  AOI21_X1  g157(.A(KEYINPUT77), .B1(new_n353_), .B2(new_n357_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n351_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n288_), .A2(new_n334_), .A3(new_n289_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n361_), .A2(new_n350_), .A3(new_n353_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G113gat), .B(G141gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G169gat), .B(G197gat), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n363_), .B(new_n364_), .Z(new_n365_));
  NAND3_X1  g164(.A1(new_n360_), .A2(new_n362_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT79), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n366_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n368_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n362_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT77), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n334_), .A2(new_n356_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n352_), .A2(new_n286_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n372_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n353_), .A2(new_n357_), .A3(KEYINPUT77), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n371_), .B1(new_n377_), .B2(new_n351_), .ZN(new_n378_));
  OAI22_X1  g177(.A1(new_n369_), .A2(new_n370_), .B1(new_n378_), .B2(new_n365_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n366_), .A2(new_n367_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT79), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n378_), .A2(new_n365_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n366_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n379_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G227gat), .A2(G233gat), .ZN(new_n386_));
  INV_X1    g185(.A(G15gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT30), .ZN(new_n389_));
  INV_X1    g188(.A(G169gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT22), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT22), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(G169gat), .ZN(new_n393_));
  INV_X1    g192(.A(G176gat), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n391_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT81), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G169gat), .A2(G176gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G183gat), .A2(G190gat), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT23), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  OR2_X1    g199(.A1(G183gat), .A2(G190gat), .ZN(new_n401_));
  NAND3_X1  g200(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT81), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n391_), .A2(new_n393_), .A3(new_n404_), .A4(new_n394_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n396_), .A2(new_n397_), .A3(new_n403_), .A4(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT26), .B(G190gat), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT25), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n408_), .A2(KEYINPUT80), .A3(G183gat), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT80), .ZN(new_n410_));
  INV_X1    g209(.A(G183gat), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT25), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n407_), .A2(new_n409_), .A3(new_n412_), .ZN(new_n413_));
  AND2_X1   g212(.A1(new_n400_), .A2(new_n402_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n390_), .A2(new_n394_), .ZN(new_n415_));
  OR2_X1    g214(.A1(new_n415_), .A2(KEYINPUT24), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n415_), .A2(KEYINPUT24), .A3(new_n397_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n413_), .A2(new_n414_), .A3(new_n416_), .A4(new_n417_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n406_), .A2(new_n418_), .A3(KEYINPUT82), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT82), .B1(new_n406_), .B2(new_n418_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G71gat), .B(G99gat), .ZN(new_n422_));
  INV_X1    g221(.A(G43gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n421_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n406_), .A2(new_n418_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT82), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n406_), .A2(new_n418_), .A3(KEYINPUT82), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n424_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n389_), .B1(new_n426_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n426_), .A2(new_n432_), .A3(new_n389_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n434_), .A2(KEYINPUT83), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT83), .ZN(new_n437_));
  INV_X1    g236(.A(new_n435_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n437_), .B1(new_n438_), .B2(new_n433_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G127gat), .B(G134gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G113gat), .B(G120gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT31), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n436_), .A2(new_n439_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n443_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n437_), .B(new_n445_), .C1(new_n438_), .C2(new_n433_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n444_), .A2(KEYINPUT84), .A3(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT84), .B1(new_n444_), .B2(new_n446_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G228gat), .A2(G233gat), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT29), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G141gat), .B(G148gat), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G155gat), .A2(G162gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT1), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT86), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT86), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n455_), .A2(new_n458_), .A3(KEYINPUT1), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(G155gat), .ZN(new_n461_));
  INV_X1    g260(.A(G162gat), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(new_n462_), .A3(KEYINPUT85), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT85), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n464_), .B1(G155gat), .B2(G162gat), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT1), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(G155gat), .A3(G162gat), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n463_), .A2(new_n465_), .A3(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n454_), .B1(new_n460_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT3), .ZN(new_n470_));
  INV_X1    g269(.A(G141gat), .ZN(new_n471_));
  INV_X1    g270(.A(G148gat), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n470_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G141gat), .A2(G148gat), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT2), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n473_), .A2(new_n476_), .A3(new_n477_), .A4(new_n478_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n479_), .A2(new_n463_), .A3(new_n465_), .A4(new_n455_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n452_), .B1(new_n469_), .B2(new_n480_), .ZN(new_n481_));
  OR2_X1    g280(.A1(G197gat), .A2(G204gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G197gat), .A2(G204gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT21), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n482_), .A2(KEYINPUT21), .A3(new_n483_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G211gat), .B(G218gat), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n487_), .A2(new_n488_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n451_), .B1(new_n481_), .B2(new_n492_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n455_), .A2(new_n458_), .A3(KEYINPUT1), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n458_), .B1(new_n455_), .B2(KEYINPUT1), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n463_), .A2(new_n465_), .A3(new_n467_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n453_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n463_), .A2(new_n465_), .A3(new_n455_), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n473_), .A2(new_n478_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n476_), .A2(new_n477_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n499_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT29), .B1(new_n498_), .B2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n503_), .A2(new_n491_), .A3(new_n450_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n493_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G78gat), .B(G106gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n506_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n493_), .A2(new_n504_), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G22gat), .B(G50gat), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n469_), .A2(new_n452_), .A3(new_n480_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT87), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT87), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n469_), .A2(new_n480_), .A3(new_n515_), .A4(new_n452_), .ZN(new_n516_));
  XOR2_X1   g315(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n514_), .A2(new_n516_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n518_), .B1(new_n514_), .B2(new_n516_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n512_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n521_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n523_), .A2(new_n511_), .A3(new_n519_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n510_), .A2(new_n522_), .A3(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT89), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n510_), .A2(new_n522_), .A3(new_n524_), .A4(KEYINPUT89), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n509_), .A2(KEYINPUT91), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT91), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n493_), .A2(new_n504_), .A3(new_n531_), .A4(new_n508_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT90), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n534_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n535_));
  AOI211_X1 g334(.A(KEYINPUT90), .B(new_n508_), .C1(new_n493_), .C2(new_n504_), .ZN(new_n536_));
  NOR3_X1   g335(.A1(new_n533_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n522_), .A2(new_n524_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n529_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT33), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G1gat), .B(G29gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(G85gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT0), .B(G57gat), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n543_), .B(new_n544_), .Z(new_n545_));
  AND2_X1   g344(.A1(new_n440_), .A2(new_n441_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n440_), .A2(new_n441_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n548_), .B1(new_n498_), .B2(new_n502_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n469_), .A2(new_n442_), .A3(new_n480_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G225gat), .A2(G233gat), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n549_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n545_), .A2(new_n552_), .ZN(new_n553_));
  AND3_X1   g352(.A1(new_n549_), .A2(KEYINPUT4), .A3(new_n550_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n551_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n555_), .B1(new_n549_), .B2(KEYINPUT4), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT93), .B1(new_n554_), .B2(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n442_), .B1(new_n469_), .B2(new_n480_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT4), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n551_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT93), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n549_), .A2(new_n550_), .A3(KEYINPUT4), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n560_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n553_), .B1(new_n557_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT94), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n541_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  AOI211_X1 g365(.A(KEYINPUT94), .B(new_n553_), .C1(new_n557_), .C2(new_n563_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT95), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n553_), .ZN(new_n569_));
  NOR3_X1   g368(.A1(new_n554_), .A2(new_n556_), .A3(KEYINPUT93), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n561_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n569_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT94), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n564_), .A2(new_n565_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT95), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .A4(new_n541_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G226gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT19), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n419_), .A2(new_n420_), .A3(new_n491_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT20), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n414_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT25), .B(G183gat), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n407_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n403_), .A2(new_n397_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n395_), .ZN(new_n586_));
  OAI22_X1  g385(.A1(new_n581_), .A2(new_n584_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n580_), .B1(new_n587_), .B2(new_n491_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n578_), .B1(new_n579_), .B2(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(G8gat), .B(G36gat), .Z(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G64gat), .B(G92gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n491_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n587_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n580_), .B1(new_n597_), .B2(new_n492_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n578_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n596_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n590_), .A2(new_n595_), .A3(new_n600_), .ZN(new_n601_));
  OAI211_X1 g400(.A(KEYINPUT33), .B(new_n569_), .C1(new_n570_), .C2(new_n571_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n595_), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n596_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n429_), .A2(new_n430_), .A3(new_n492_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n599_), .B1(new_n605_), .B2(new_n588_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n603_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n545_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n549_), .A2(new_n550_), .A3(new_n555_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n551_), .B1(new_n549_), .B2(KEYINPUT4), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n608_), .B(new_n609_), .C1(new_n554_), .C2(new_n610_), .ZN(new_n611_));
  AND4_X1   g410(.A1(new_n601_), .A2(new_n602_), .A3(new_n607_), .A4(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n568_), .A2(new_n576_), .A3(new_n612_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n605_), .A2(new_n599_), .A3(new_n588_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n599_), .B1(new_n596_), .B2(new_n598_), .ZN(new_n615_));
  OAI21_X1  g414(.A(KEYINPUT96), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n605_), .A2(new_n599_), .A3(new_n588_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT96), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n616_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(KEYINPUT32), .A3(new_n595_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n552_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n622_), .B1(new_n557_), .B2(new_n563_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n572_), .B1(new_n623_), .B2(new_n545_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n595_), .A2(KEYINPUT32), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n590_), .A2(new_n625_), .A3(new_n600_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n621_), .A2(new_n624_), .A3(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n540_), .B1(new_n613_), .B2(new_n627_), .ZN(new_n628_));
  AOI22_X1  g427(.A1(new_n527_), .A2(new_n528_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT27), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n604_), .A2(new_n606_), .A3(new_n603_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n595_), .B1(new_n590_), .B2(new_n600_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n630_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n595_), .B1(new_n616_), .B2(new_n619_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n601_), .A2(KEYINPUT27), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n633_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n629_), .A2(new_n636_), .A3(new_n624_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n449_), .B1(new_n628_), .B2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n444_), .A2(new_n446_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n540_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n624_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n636_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n640_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n385_), .B1(new_n638_), .B2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n349_), .A2(new_n644_), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n641_), .A2(G1gat), .ZN(new_n646_));
  OR3_X1    g445(.A1(new_n645_), .A2(KEYINPUT97), .A3(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(KEYINPUT97), .B1(new_n645_), .B2(new_n646_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n647_), .A2(KEYINPUT38), .A3(new_n648_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT98), .Z(new_n650_));
  AOI21_X1  g449(.A(new_n318_), .B1(new_n638_), .B2(new_n643_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n385_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n651_), .A2(new_n652_), .A3(new_n347_), .A4(new_n274_), .ZN(new_n653_));
  OAI21_X1  g452(.A(G1gat), .B1(new_n653_), .B2(new_n641_), .ZN(new_n654_));
  AOI21_X1  g453(.A(KEYINPUT38), .B1(new_n647_), .B2(new_n648_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT99), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n655_), .A2(new_n656_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n650_), .B(new_n654_), .C1(new_n657_), .C2(new_n658_), .ZN(G1324gat));
  OAI21_X1  g458(.A(G8gat), .B1(new_n653_), .B2(new_n642_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT39), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n642_), .A2(G8gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n661_), .B1(new_n645_), .B2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n663_), .B(new_n664_), .Z(G1325gat));
  OAI21_X1  g464(.A(G15gat), .B1(new_n653_), .B2(new_n449_), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n666_), .B(KEYINPUT41), .Z(new_n667_));
  INV_X1    g466(.A(new_n645_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n449_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(new_n387_), .A3(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n667_), .A2(new_n670_), .ZN(G1326gat));
  OAI21_X1  g470(.A(G22gat), .B1(new_n653_), .B2(new_n629_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n672_), .B(new_n673_), .Z(new_n674_));
  NOR3_X1   g473(.A1(new_n645_), .A2(G22gat), .A3(new_n629_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1327gat));
  OR2_X1    g475(.A1(new_n272_), .A2(new_n273_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n346_), .A2(new_n318_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(new_n644_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT104), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT104), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n679_), .A2(new_n682_), .A3(new_n644_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n681_), .A2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G29gat), .B1(new_n684_), .B2(new_n624_), .ZN(new_n685_));
  XOR2_X1   g484(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n677_), .A2(new_n385_), .A3(new_n347_), .ZN(new_n688_));
  AOI221_X4 g487(.A(KEYINPUT43), .B1(new_n323_), .B2(new_n324_), .C1(new_n638_), .C2(new_n643_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n638_), .A2(new_n643_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n323_), .A2(new_n324_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n690_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n688_), .B1(new_n689_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n688_), .B(KEYINPUT102), .C1(new_n689_), .C2(new_n693_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n687_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n694_), .A2(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n624_), .A2(G29gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n685_), .B1(new_n701_), .B2(new_n702_), .ZN(G1328gat));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT46), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n636_), .B1(new_n694_), .B2(new_n699_), .ZN(new_n708_));
  OAI21_X1  g507(.A(G36gat), .B1(new_n698_), .B2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT105), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n711_));
  OAI211_X1 g510(.A(new_n711_), .B(G36gat), .C1(new_n698_), .C2(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n704_), .A2(new_n705_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n642_), .A2(KEYINPUT106), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n642_), .A2(KEYINPUT106), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n719_), .A2(G36gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n715_), .B1(new_n684_), .B2(new_n720_), .ZN(new_n721_));
  AND4_X1   g520(.A1(new_n681_), .A2(new_n683_), .A3(new_n715_), .A4(new_n720_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n714_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n707_), .B1(new_n713_), .B2(new_n724_), .ZN(new_n725_));
  AOI211_X1 g524(.A(new_n706_), .B(new_n723_), .C1(new_n710_), .C2(new_n712_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1329gat));
  INV_X1    g526(.A(new_n639_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n423_), .B1(new_n701_), .B2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT47), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n684_), .A2(new_n423_), .A3(new_n669_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  OR3_X1    g531(.A1(new_n729_), .A2(new_n730_), .A3(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n730_), .B1(new_n729_), .B2(new_n732_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1330gat));
  NAND2_X1  g534(.A1(new_n701_), .A2(new_n540_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n736_), .A2(KEYINPUT109), .A3(G50gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT109), .B1(new_n736_), .B2(G50gat), .ZN(new_n738_));
  INV_X1    g537(.A(new_n684_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n629_), .A2(G50gat), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT110), .Z(new_n741_));
  OAI22_X1  g540(.A1(new_n737_), .A2(new_n738_), .B1(new_n739_), .B2(new_n741_), .ZN(G1331gat));
  NOR2_X1   g541(.A1(new_n274_), .A2(new_n652_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(new_n691_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n744_), .A2(new_n692_), .A3(new_n346_), .ZN(new_n745_));
  INV_X1    g544(.A(G57gat), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n745_), .A2(new_n746_), .A3(new_n624_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n651_), .A2(new_n743_), .A3(new_n347_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G57gat), .B1(new_n748_), .B2(new_n641_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1332gat));
  OAI21_X1  g549(.A(G64gat), .B1(new_n748_), .B2(new_n719_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT48), .ZN(new_n752_));
  INV_X1    g551(.A(new_n745_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n719_), .A2(G64gat), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT111), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n752_), .B1(new_n753_), .B2(new_n755_), .ZN(G1333gat));
  OAI21_X1  g555(.A(G71gat), .B1(new_n748_), .B2(new_n449_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT49), .Z(new_n758_));
  NOR3_X1   g557(.A1(new_n753_), .A2(G71gat), .A3(new_n449_), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n758_), .A2(new_n759_), .ZN(G1334gat));
  OAI21_X1  g559(.A(G78gat), .B1(new_n748_), .B2(new_n629_), .ZN(new_n761_));
  XOR2_X1   g560(.A(new_n761_), .B(KEYINPUT50), .Z(new_n762_));
  NOR3_X1   g561(.A1(new_n753_), .A2(G78gat), .A3(new_n629_), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1335gat));
  NAND2_X1  g563(.A1(new_n743_), .A2(new_n346_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n691_), .A2(new_n692_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT43), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n691_), .A2(new_n690_), .A3(new_n692_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n765_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(G85gat), .B1(new_n770_), .B2(new_n641_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n744_), .A2(new_n678_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n772_), .A2(new_n211_), .A3(new_n624_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1336gat));
  OAI21_X1  g573(.A(G92gat), .B1(new_n770_), .B2(new_n719_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n772_), .A2(new_n212_), .A3(new_n636_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(G1337gat));
  NAND2_X1  g576(.A1(new_n769_), .A2(new_n669_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n728_), .A2(new_n225_), .ZN(new_n779_));
  AOI22_X1  g578(.A1(new_n778_), .A2(G99gat), .B1(new_n772_), .B2(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n780_), .B(new_n781_), .ZN(G1338gat));
  NAND3_X1  g581(.A1(new_n772_), .A2(new_n226_), .A3(new_n540_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n769_), .A2(new_n540_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(G106gat), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT113), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n784_), .A2(new_n788_), .A3(G106gat), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n786_), .A2(new_n787_), .A3(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n787_), .B1(new_n786_), .B2(new_n789_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n783_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT53), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n794_), .B(new_n783_), .C1(new_n790_), .C2(new_n791_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(G1339gat));
  NAND3_X1  g595(.A1(new_n640_), .A2(new_n624_), .A3(new_n642_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT120), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n799_), .A2(KEYINPUT59), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n361_), .A2(new_n353_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n350_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n803_), .B1(new_n802_), .B2(new_n801_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n365_), .B1(new_n377_), .B2(new_n350_), .ZN(new_n805_));
  AOI22_X1  g604(.A1(new_n804_), .A2(new_n805_), .B1(new_n378_), .B2(new_n365_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n267_), .A2(new_n271_), .A3(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n267_), .A2(KEYINPUT116), .A3(new_n271_), .A4(new_n806_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n252_), .B2(new_n812_), .ZN(new_n813_));
  OR2_X1    g612(.A1(new_n262_), .A2(new_n251_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n262_), .A2(KEYINPUT114), .A3(KEYINPUT55), .A4(new_n251_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n252_), .A2(new_n812_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n813_), .A2(new_n814_), .A3(new_n815_), .A4(new_n816_), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n817_), .A2(KEYINPUT56), .A3(new_n259_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT56), .B1(new_n817_), .B2(new_n259_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n379_), .A2(new_n384_), .A3(new_n260_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n809_), .B(new_n810_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n318_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n822_), .A2(KEYINPUT57), .A3(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n822_), .A2(new_n823_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n806_), .A2(new_n260_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n829_), .B(new_n830_), .C1(new_n818_), .C2(new_n819_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT58), .B1(new_n831_), .B2(KEYINPUT118), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT117), .B1(KEYINPUT118), .B2(KEYINPUT58), .ZN(new_n833_));
  INV_X1    g632(.A(new_n819_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n817_), .A2(KEYINPUT56), .A3(new_n259_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n833_), .B1(new_n836_), .B2(new_n829_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n692_), .B1(new_n832_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n828_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT123), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n825_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n828_), .A2(KEYINPUT123), .A3(new_n838_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n347_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT54), .B1(new_n348_), .B2(new_n652_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n692_), .A2(new_n346_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n845_), .A2(new_n846_), .A3(new_n385_), .A4(new_n274_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n844_), .A2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n800_), .B1(new_n843_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n838_), .A2(new_n850_), .ZN(new_n851_));
  OAI211_X1 g650(.A(KEYINPUT119), .B(new_n692_), .C1(new_n832_), .C2(new_n837_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n851_), .A2(new_n828_), .A3(new_n852_), .A4(new_n824_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n848_), .B1(new_n853_), .B2(new_n346_), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT59), .B1(new_n854_), .B2(new_n799_), .ZN(new_n855_));
  AND4_X1   g654(.A1(G113gat), .A2(new_n849_), .A3(new_n652_), .A4(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n853_), .A2(new_n346_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n848_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(new_n860_), .A3(new_n798_), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT121), .B1(new_n854_), .B2(new_n799_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n861_), .A2(new_n862_), .A3(new_n652_), .ZN(new_n863_));
  INV_X1    g662(.A(G113gat), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n863_), .A2(KEYINPUT122), .A3(new_n864_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n856_), .B1(new_n867_), .B2(new_n868_), .ZN(G1340gat));
  NAND2_X1  g668(.A1(new_n849_), .A2(new_n855_), .ZN(new_n870_));
  OAI21_X1  g669(.A(G120gat), .B1(new_n870_), .B2(new_n274_), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n861_), .A2(new_n862_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n274_), .A2(KEYINPUT60), .ZN(new_n873_));
  MUX2_X1   g672(.A(new_n873_), .B(KEYINPUT60), .S(G120gat), .Z(new_n874_));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n871_), .A2(new_n875_), .ZN(G1341gat));
  OAI21_X1  g675(.A(G127gat), .B1(new_n870_), .B2(new_n346_), .ZN(new_n877_));
  INV_X1    g676(.A(G127gat), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n872_), .A2(new_n878_), .A3(new_n347_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n879_), .ZN(G1342gat));
  AOI21_X1  g679(.A(G134gat), .B1(new_n872_), .B2(new_n318_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n870_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n692_), .A2(G134gat), .ZN(new_n883_));
  XOR2_X1   g682(.A(new_n883_), .B(KEYINPUT124), .Z(new_n884_));
  AOI21_X1  g683(.A(new_n881_), .B1(new_n882_), .B2(new_n884_), .ZN(G1343gat));
  NOR3_X1   g684(.A1(new_n854_), .A2(new_n669_), .A3(new_n629_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n718_), .A2(new_n641_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n886_), .A2(new_n652_), .A3(new_n887_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g688(.A1(new_n886_), .A2(new_n677_), .A3(new_n887_), .ZN(new_n890_));
  XOR2_X1   g689(.A(KEYINPUT125), .B(G148gat), .Z(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1345gat));
  NAND3_X1  g691(.A1(new_n886_), .A2(new_n347_), .A3(new_n887_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT61), .B(G155gat), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1346gat));
  AND2_X1   g694(.A1(new_n886_), .A2(new_n887_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(new_n462_), .A3(new_n318_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n896_), .A2(new_n692_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n898_), .B2(new_n462_), .ZN(G1347gat));
  NAND2_X1  g698(.A1(new_n841_), .A2(new_n842_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n848_), .B1(new_n900_), .B2(new_n346_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n719_), .A2(new_n624_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n669_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n540_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n902_), .A2(new_n905_), .ZN(new_n906_));
  OAI211_X1 g705(.A(KEYINPUT62), .B(G169gat), .C1(new_n906_), .C2(new_n385_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n908_));
  INV_X1    g707(.A(new_n905_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n901_), .A2(new_n385_), .A3(new_n909_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n908_), .B1(new_n910_), .B2(new_n390_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n910_), .A2(new_n391_), .A3(new_n393_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n907_), .A2(new_n911_), .A3(new_n912_), .ZN(G1348gat));
  NAND3_X1  g712(.A1(new_n902_), .A2(new_n677_), .A3(new_n905_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n854_), .A2(new_n540_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n904_), .A2(new_n394_), .A3(new_n274_), .ZN(new_n916_));
  AOI22_X1  g715(.A1(new_n914_), .A2(new_n394_), .B1(new_n915_), .B2(new_n916_), .ZN(G1349gat));
  NOR2_X1   g716(.A1(new_n346_), .A2(new_n582_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n902_), .A2(new_n905_), .A3(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n904_), .A2(new_n346_), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n915_), .A2(new_n920_), .ZN(new_n921_));
  OAI211_X1 g720(.A(new_n919_), .B(KEYINPUT126), .C1(G183gat), .C2(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT126), .ZN(new_n923_));
  NOR4_X1   g722(.A1(new_n901_), .A2(new_n582_), .A3(new_n346_), .A4(new_n909_), .ZN(new_n924_));
  AOI21_X1  g723(.A(G183gat), .B1(new_n915_), .B2(new_n920_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n923_), .B1(new_n924_), .B2(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n922_), .A2(new_n926_), .ZN(G1350gat));
  AND2_X1   g726(.A1(new_n323_), .A2(new_n324_), .ZN(new_n928_));
  OAI21_X1  g727(.A(G190gat), .B1(new_n906_), .B2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n318_), .A2(new_n407_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n906_), .B2(new_n930_), .ZN(G1351gat));
  NAND3_X1  g730(.A1(new_n886_), .A2(new_n652_), .A3(new_n903_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g732(.A1(new_n886_), .A2(new_n903_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n934_), .A2(new_n274_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  XOR2_X1   g736(.A(KEYINPUT127), .B(G204gat), .Z(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n935_), .B2(new_n938_), .ZN(G1353gat));
  NOR2_X1   g738(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n940_));
  INV_X1    g739(.A(new_n940_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n934_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n346_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n941_), .B1(new_n942_), .B2(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(new_n943_), .ZN(new_n945_));
  NOR3_X1   g744(.A1(new_n934_), .A2(new_n940_), .A3(new_n945_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n944_), .A2(new_n946_), .ZN(G1354gat));
  OR3_X1    g746(.A1(new_n934_), .A2(G218gat), .A3(new_n823_), .ZN(new_n948_));
  OAI21_X1  g747(.A(G218gat), .B1(new_n934_), .B2(new_n928_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n948_), .A2(new_n949_), .ZN(G1355gat));
endmodule


