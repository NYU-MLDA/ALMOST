//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 1 1 1 0 1 0 1 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n800_, new_n801_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n930_, new_n931_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n953_, new_n955_, new_n956_, new_n957_, new_n959_, new_n960_,
    new_n961_, new_n963_, new_n964_, new_n965_, new_n967_, new_n968_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n980_, new_n981_, new_n982_;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G64gat), .B(G92gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G211gat), .B(G218gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G197gat), .A2(G204gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT88), .B(G204gat), .ZN(new_n211_));
  INV_X1    g010(.A(G197gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n210_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT21), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n208_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT89), .ZN(new_n216_));
  INV_X1    g015(.A(G204gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(KEYINPUT87), .A3(G197gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT87), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n219_), .B1(new_n212_), .B2(G204gat), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n218_), .B(new_n220_), .C1(new_n211_), .C2(G197gat), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n216_), .B1(new_n221_), .B2(KEYINPUT21), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n217_), .A2(KEYINPUT88), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT88), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(G204gat), .ZN(new_n225_));
  AOI21_X1  g024(.A(G197gat), .B1(new_n223_), .B2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n220_), .A2(new_n218_), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n216_), .B(KEYINPUT21), .C1(new_n226_), .C2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n215_), .B1(new_n222_), .B2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(G183gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT25), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT25), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(G183gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT26), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n235_), .A2(G190gat), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n232_), .B(new_n234_), .C1(new_n236_), .C2(KEYINPUT78), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT78), .ZN(new_n238_));
  INV_X1    g037(.A(G190gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT26), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n235_), .A2(G190gat), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n238_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n237_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(G169gat), .ZN(new_n248_));
  INV_X1    g047(.A(G176gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G169gat), .A2(G176gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(KEYINPUT24), .A3(new_n251_), .ZN(new_n252_));
  NOR3_X1   g051(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n247_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n243_), .A2(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(new_n248_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G183gat), .A2(G190gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT23), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n231_), .A2(new_n239_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n261_), .A2(new_n244_), .A3(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT79), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n261_), .A2(new_n262_), .A3(KEYINPUT79), .A4(new_n244_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n258_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT80), .B1(new_n256_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n266_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n257_), .B(G169gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT80), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n253_), .B1(new_n274_), .B2(new_n251_), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n275_), .B(new_n247_), .C1(new_n237_), .C2(new_n242_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n271_), .A2(new_n272_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT90), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT21), .B1(new_n208_), .B2(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n207_), .A2(KEYINPUT90), .ZN(new_n280_));
  NOR3_X1   g079(.A1(new_n279_), .A2(new_n213_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n230_), .A2(new_n268_), .A3(new_n277_), .A4(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n240_), .A2(new_n241_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n232_), .A2(new_n234_), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n275_), .B(new_n247_), .C1(new_n284_), .C2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n270_), .A2(new_n263_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n287_), .A2(KEYINPUT95), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT95), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n289_), .B1(new_n270_), .B2(new_n263_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n286_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n223_), .A2(new_n225_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n209_), .B1(new_n292_), .B2(G197gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n207_), .B1(new_n293_), .B2(KEYINPUT21), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT21), .B1(new_n226_), .B2(new_n227_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT89), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n294_), .B1(new_n296_), .B2(new_n228_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n291_), .B1(new_n297_), .B2(new_n281_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n283_), .A2(KEYINPUT20), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G226gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT19), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n301_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT20), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n297_), .A2(new_n281_), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n286_), .A2(KEYINPUT99), .A3(new_n287_), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT99), .B1(new_n286_), .B2(new_n287_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n304_), .B1(new_n305_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n268_), .A2(new_n277_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n230_), .A2(new_n282_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n303_), .B1(new_n309_), .B2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n206_), .B1(new_n302_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n299_), .A2(new_n301_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n206_), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n288_), .A2(new_n290_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n317_), .A2(new_n230_), .A3(new_n282_), .A4(new_n286_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n301_), .A2(new_n304_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n312_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n315_), .A2(new_n316_), .A3(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n314_), .A2(KEYINPUT27), .A3(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G1gat), .B(G29gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(G85gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT0), .B(G57gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(G127gat), .B(G134gat), .Z(new_n327_));
  XNOR2_X1  g126(.A(G113gat), .B(G120gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n330_));
  INV_X1    g129(.A(G141gat), .ZN(new_n331_));
  INV_X1    g130(.A(G148gat), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n331_), .A2(new_n332_), .A3(KEYINPUT3), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT3), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n334_), .B1(G141gat), .B2(G148gat), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n330_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT83), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT83), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n339_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  AND3_X1   g140(.A1(new_n336_), .A2(KEYINPUT84), .A3(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(KEYINPUT84), .B1(new_n336_), .B2(new_n341_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G155gat), .B(G162gat), .ZN(new_n344_));
  NOR3_X1   g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n344_), .A2(KEYINPUT1), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n331_), .A2(new_n332_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G141gat), .A2(G148gat), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n347_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n346_), .A2(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n329_), .B1(new_n345_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n330_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n333_), .A2(new_n335_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n341_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT84), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n344_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n336_), .A2(KEYINPUT84), .A3(new_n341_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n351_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n329_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n359_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n352_), .A2(new_n362_), .B1(G225gat), .B2(G233gat), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n352_), .A2(KEYINPUT4), .A3(new_n362_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n361_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT4), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n365_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G225gat), .A2(G233gat), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n326_), .B(new_n364_), .C1(new_n369_), .C2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n326_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n370_), .B1(new_n365_), .B2(new_n368_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n372_), .B1(new_n373_), .B2(new_n363_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n371_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT100), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n304_), .B1(new_n311_), .B2(new_n291_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n303_), .B1(new_n377_), .B2(new_n283_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n319_), .B1(new_n311_), .B2(new_n291_), .ZN(new_n379_));
  AOI22_X1  g178(.A1(new_n268_), .A2(new_n277_), .B1(new_n230_), .B2(new_n282_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n206_), .B1(new_n378_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(new_n321_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT27), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n376_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  AOI211_X1 g184(.A(KEYINPUT100), .B(KEYINPUT27), .C1(new_n382_), .C2(new_n321_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n322_), .B(new_n375_), .C1(new_n385_), .C2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT91), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n351_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT29), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n388_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  OAI211_X1 g190(.A(KEYINPUT91), .B(KEYINPUT29), .C1(new_n345_), .C2(new_n351_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n392_), .A3(new_n311_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT92), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G228gat), .A2(G233gat), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  AND3_X1   g195(.A1(new_n393_), .A2(new_n394_), .A3(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n394_), .B1(new_n393_), .B2(new_n396_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n396_), .B1(new_n230_), .B2(new_n282_), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT86), .B1(new_n389_), .B2(new_n390_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT86), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n401_), .B(KEYINPUT29), .C1(new_n345_), .C2(new_n351_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n399_), .A2(new_n400_), .A3(new_n402_), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n397_), .A2(new_n398_), .A3(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G78gat), .B(G106gat), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT94), .B1(new_n404_), .B2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n389_), .A2(new_n390_), .ZN(new_n408_));
  XOR2_X1   g207(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  XOR2_X1   g209(.A(G22gat), .B(G50gat), .Z(new_n411_));
  INV_X1    g210(.A(new_n409_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n389_), .A2(new_n390_), .A3(new_n412_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n410_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n411_), .B1(new_n410_), .B2(new_n413_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n416_), .B1(new_n404_), .B2(new_n406_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n393_), .A2(new_n396_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT92), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n393_), .A2(new_n394_), .A3(new_n396_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n403_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n419_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT94), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(new_n423_), .A3(new_n405_), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n407_), .A2(new_n417_), .A3(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n403_), .B1(new_n418_), .B2(KEYINPUT92), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT93), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n426_), .A2(new_n427_), .A3(new_n406_), .A4(new_n420_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n416_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n419_), .A2(new_n406_), .A3(new_n420_), .A4(new_n421_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n427_), .B1(new_n422_), .B2(new_n405_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n429_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n387_), .B1(new_n425_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G227gat), .A2(G233gat), .ZN(new_n434_));
  INV_X1    g233(.A(G71gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(G99gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n310_), .B(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(new_n329_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G15gat), .B(G43gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT30), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT31), .ZN(new_n444_));
  XOR2_X1   g243(.A(new_n439_), .B(new_n444_), .Z(new_n445_));
  AND2_X1   g244(.A1(new_n428_), .A2(new_n416_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n422_), .A2(new_n405_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(KEYINPUT93), .A3(new_n430_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n362_), .ZN(new_n450_));
  NOR3_X1   g249(.A1(new_n450_), .A2(new_n366_), .A3(new_n370_), .ZN(new_n451_));
  AOI211_X1 g250(.A(new_n372_), .B(new_n451_), .C1(new_n369_), .C2(new_n370_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n452_), .B1(new_n383_), .B2(KEYINPUT97), .ZN(new_n453_));
  NOR2_X1   g252(.A1(KEYINPUT98), .A2(KEYINPUT33), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n374_), .A2(new_n454_), .ZN(new_n455_));
  OAI221_X1 g254(.A(new_n372_), .B1(KEYINPUT98), .B2(KEYINPUT33), .C1(new_n373_), .C2(new_n363_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT97), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n382_), .A2(new_n458_), .A3(new_n321_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n453_), .A2(new_n457_), .A3(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n407_), .A2(new_n417_), .A3(new_n424_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n316_), .A2(KEYINPUT32), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n315_), .A2(new_n320_), .A3(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n302_), .A2(new_n313_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n463_), .B1(new_n464_), .B2(new_n462_), .ZN(new_n465_));
  OR2_X1    g264(.A1(new_n375_), .A2(new_n465_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n449_), .A2(new_n460_), .A3(new_n461_), .A4(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n433_), .A2(new_n445_), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n375_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n445_), .A2(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n423_), .B1(new_n422_), .B2(new_n405_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n416_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n430_), .A2(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  AOI22_X1  g273(.A1(new_n474_), .A2(new_n424_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n322_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n315_), .A2(new_n316_), .A3(new_n320_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n316_), .B1(new_n315_), .B2(new_n320_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n384_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT100), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n383_), .A2(new_n376_), .A3(new_n384_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n476_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n470_), .A2(new_n475_), .A3(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n468_), .A2(new_n483_), .ZN(new_n484_));
  OR2_X1    g283(.A1(G85gat), .A2(G92gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G85gat), .A2(G92gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT65), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n485_), .A2(KEYINPUT65), .A3(new_n486_), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G99gat), .A2(G106gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT6), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT7), .ZN(new_n495_));
  INV_X1    g294(.A(G99gat), .ZN(new_n496_));
  INV_X1    g295(.A(G106gat), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n493_), .A2(new_n494_), .A3(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n491_), .A2(KEYINPUT66), .A3(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT66), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT6), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n492_), .B(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n498_), .A2(new_n494_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n489_), .A2(new_n490_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n501_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n500_), .A2(new_n507_), .A3(KEYINPUT8), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT9), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n493_), .B1(new_n509_), .B2(new_n487_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT10), .B(G99gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT64), .B(G92gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n509_), .A2(G85gat), .ZN(new_n513_));
  OAI22_X1  g312(.A1(G106gat), .A2(new_n511_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  OAI22_X1  g313(.A1(new_n507_), .A2(KEYINPUT8), .B1(new_n510_), .B2(new_n514_), .ZN(new_n515_));
  NOR3_X1   g314(.A1(new_n508_), .A2(new_n515_), .A3(KEYINPUT67), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT67), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n510_), .A2(new_n514_), .ZN(new_n518_));
  AOI21_X1  g317(.A(KEYINPUT66), .B1(new_n491_), .B2(new_n499_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT8), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n518_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n500_), .A2(new_n507_), .A3(KEYINPUT8), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n517_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n516_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G57gat), .B(G64gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G71gat), .B(G78gat), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n525_), .A2(new_n526_), .A3(KEYINPUT11), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(KEYINPUT11), .ZN(new_n528_));
  INV_X1    g327(.A(new_n526_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n525_), .A2(KEYINPUT11), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n527_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n532_), .B(KEYINPUT68), .Z(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT12), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n532_), .A2(KEYINPUT69), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT69), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n537_), .B(new_n527_), .C1(new_n530_), .C2(new_n531_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n535_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n539_), .B1(new_n508_), .B2(new_n515_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT70), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n521_), .A2(new_n522_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n543_), .A2(KEYINPUT70), .A3(new_n539_), .ZN(new_n544_));
  AOI22_X1  g343(.A1(new_n524_), .A2(new_n534_), .B1(new_n542_), .B2(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT67), .B1(new_n508_), .B2(new_n515_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n521_), .A2(new_n517_), .A3(new_n522_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(new_n533_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(new_n535_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G230gat), .A2(G233gat), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n545_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n534_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n549_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n551_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(G176gat), .B(G204gat), .Z(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT72), .ZN(new_n558_));
  XOR2_X1   g357(.A(KEYINPUT71), .B(KEYINPUT5), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G120gat), .B(G148gat), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n560_), .B(new_n561_), .Z(new_n562_));
  NAND3_X1  g361(.A1(new_n552_), .A2(new_n556_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n562_), .B1(new_n552_), .B2(new_n556_), .ZN(new_n565_));
  OAI21_X1  g364(.A(KEYINPUT13), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n565_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT13), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(new_n568_), .A3(new_n563_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n566_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT37), .ZN(new_n571_));
  XOR2_X1   g370(.A(G29gat), .B(G36gat), .Z(new_n572_));
  XOR2_X1   g371(.A(G43gat), .B(G50gat), .Z(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT15), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT35), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G232gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT34), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  AOI22_X1  g378(.A1(new_n543_), .A2(new_n575_), .B1(new_n576_), .B2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n574_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n580_), .B1(new_n548_), .B2(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n579_), .A2(new_n576_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  OAI221_X1 g383(.A(new_n580_), .B1(new_n576_), .B2(new_n579_), .C1(new_n548_), .C2(new_n581_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G190gat), .B(G218gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G134gat), .B(G162gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n588_), .A2(KEYINPUT36), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n584_), .A2(new_n585_), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n588_), .B(KEYINPUT36), .Z(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n593_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n594_));
  OAI211_X1 g393(.A(KEYINPUT73), .B(new_n571_), .C1(new_n591_), .C2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n594_), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n571_), .A2(KEYINPUT73), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n571_), .A2(KEYINPUT73), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n596_), .A2(new_n590_), .A3(new_n597_), .A4(new_n598_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n595_), .A2(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(G127gat), .B(G155gat), .Z(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT16), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G183gat), .B(G211gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G1gat), .A2(G8gat), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT14), .ZN(new_n606_));
  INV_X1    g405(.A(G15gat), .ZN(new_n607_));
  INV_X1    g406(.A(G22gat), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(G15gat), .A2(G22gat), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n606_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT74), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT74), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n613_), .B(new_n606_), .C1(new_n609_), .C2(new_n610_), .ZN(new_n614_));
  XOR2_X1   g413(.A(G1gat), .B(G8gat), .Z(new_n615_));
  NAND3_X1  g414(.A1(new_n612_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n615_), .B1(new_n612_), .B2(new_n614_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G231gat), .A2(G233gat), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n619_), .B(new_n620_), .Z(new_n621_));
  NAND2_X1  g420(.A1(new_n536_), .A2(new_n538_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n621_), .A2(new_n623_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n626_));
  OR4_X1    g425(.A1(new_n604_), .A2(new_n624_), .A3(new_n625_), .A4(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n621_), .B(new_n534_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n604_), .B(KEYINPUT17), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n627_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n570_), .A2(new_n600_), .A3(new_n632_), .ZN(new_n633_));
  OR3_X1    g432(.A1(new_n619_), .A2(KEYINPUT76), .A3(new_n574_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n581_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n618_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n636_), .A2(new_n616_), .A3(new_n574_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n635_), .A2(new_n637_), .A3(KEYINPUT76), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n634_), .A2(G229gat), .A3(G233gat), .A4(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n575_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(G229gat), .A2(G233gat), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(new_n641_), .A3(new_n637_), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT77), .B1(new_n639_), .B2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(G113gat), .B(G141gat), .ZN(new_n644_));
  XNOR2_X1  g443(.A(G169gat), .B(G197gat), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n644_), .B(new_n645_), .Z(new_n646_));
  NOR2_X1   g445(.A1(new_n643_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n646_), .ZN(new_n648_));
  AOI211_X1 g447(.A(KEYINPUT77), .B(new_n648_), .C1(new_n639_), .C2(new_n642_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n484_), .A2(new_n633_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT101), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n484_), .A2(new_n633_), .A3(KEYINPUT101), .A4(new_n650_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n375_), .A2(G1gat), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n653_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT38), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n445_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n375_), .A2(new_n465_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n459_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n661_), .B2(new_n453_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n659_), .B1(new_n475_), .B2(new_n662_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n482_), .A2(new_n461_), .A3(new_n449_), .ZN(new_n664_));
  AOI22_X1  g463(.A1(new_n663_), .A2(new_n433_), .B1(new_n664_), .B2(new_n470_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n596_), .A2(new_n590_), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n666_), .B(KEYINPUT102), .Z(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n665_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n570_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n650_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n670_), .A2(new_n671_), .A3(new_n631_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n669_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G1gat), .B1(new_n674_), .B2(new_n375_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n656_), .A2(new_n657_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n658_), .A2(new_n675_), .A3(new_n676_), .ZN(G1324gat));
  NOR2_X1   g476(.A1(new_n482_), .A2(G8gat), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n653_), .A2(new_n654_), .A3(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(KEYINPUT103), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n653_), .A2(new_n681_), .A3(new_n654_), .A4(new_n678_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n482_), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n672_), .A2(new_n484_), .A3(new_n684_), .A4(new_n667_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(G8gat), .ZN(new_n686_));
  XOR2_X1   g485(.A(KEYINPUT104), .B(KEYINPUT39), .Z(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n683_), .A2(new_n688_), .A3(KEYINPUT105), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT105), .B1(new_n683_), .B2(new_n688_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n689_), .A2(new_n690_), .A3(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n683_), .A2(new_n688_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n683_), .A2(new_n688_), .A3(KEYINPUT105), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n691_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n693_), .A2(new_n698_), .ZN(G1325gat));
  OAI21_X1  g498(.A(G15gat), .B1(new_n674_), .B2(new_n445_), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n700_), .A2(KEYINPUT41), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(KEYINPUT41), .ZN(new_n702_));
  INV_X1    g501(.A(new_n651_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n703_), .A2(new_n607_), .A3(new_n659_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT107), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n701_), .A2(new_n702_), .A3(new_n705_), .ZN(G1326gat));
  INV_X1    g505(.A(new_n475_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n608_), .B1(new_n673_), .B2(new_n707_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT42), .Z(new_n709_));
  NAND3_X1  g508(.A1(new_n703_), .A2(new_n608_), .A3(new_n707_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1327gat));
  INV_X1    g510(.A(G29gat), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n670_), .A2(new_n671_), .A3(new_n632_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT43), .ZN(new_n714_));
  INV_X1    g513(.A(new_n600_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n484_), .B2(new_n715_), .ZN(new_n716_));
  AOI211_X1 g515(.A(KEYINPUT43), .B(new_n600_), .C1(new_n468_), .C2(new_n483_), .ZN(new_n717_));
  OAI211_X1 g516(.A(KEYINPUT44), .B(new_n713_), .C1(new_n716_), .C2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n713_), .ZN(new_n720_));
  OAI21_X1  g519(.A(KEYINPUT43), .B1(new_n665_), .B2(new_n600_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n484_), .A2(new_n714_), .A3(new_n715_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n720_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(KEYINPUT108), .B1(new_n723_), .B2(KEYINPUT44), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n713_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n725_), .A2(new_n726_), .A3(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n719_), .B1(new_n724_), .B2(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n712_), .B1(new_n729_), .B2(new_n469_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n632_), .A2(new_n666_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n570_), .A2(new_n731_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n665_), .A2(new_n671_), .A3(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n733_), .A2(new_n712_), .A3(new_n469_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(KEYINPUT109), .B1(new_n730_), .B2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT109), .ZN(new_n737_));
  AOI211_X1 g536(.A(new_n375_), .B(new_n719_), .C1(new_n724_), .C2(new_n728_), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n737_), .B(new_n734_), .C1(new_n738_), .C2(new_n712_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n736_), .A2(new_n739_), .ZN(G1328gat));
  INV_X1    g539(.A(G36gat), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n733_), .A2(new_n741_), .A3(new_n684_), .ZN(new_n742_));
  XOR2_X1   g541(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n718_), .A2(new_n684_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n724_), .B2(new_n728_), .ZN(new_n746_));
  OAI211_X1 g545(.A(KEYINPUT111), .B(new_n744_), .C1(new_n746_), .C2(new_n741_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT112), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT46), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n744_), .B1(new_n746_), .B2(new_n741_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT112), .ZN(new_n751_));
  OAI21_X1  g550(.A(KEYINPUT111), .B1(new_n751_), .B2(new_n749_), .ZN(new_n752_));
  AOI22_X1  g551(.A1(new_n748_), .A2(new_n749_), .B1(new_n750_), .B2(new_n752_), .ZN(G1329gat));
  NAND3_X1  g552(.A1(new_n729_), .A2(G43gat), .A3(new_n659_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n733_), .A2(new_n659_), .ZN(new_n755_));
  XOR2_X1   g554(.A(KEYINPUT113), .B(G43gat), .Z(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT114), .Z(new_n758_));
  NAND2_X1  g557(.A1(new_n754_), .A2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT47), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT47), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n754_), .A2(new_n758_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1330gat));
  INV_X1    g562(.A(G50gat), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n707_), .A2(new_n764_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT115), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n733_), .A2(new_n766_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n729_), .A2(new_n707_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(new_n764_), .ZN(G1331gat));
  NAND2_X1  g568(.A1(new_n670_), .A2(new_n632_), .ZN(new_n770_));
  NOR4_X1   g569(.A1(new_n665_), .A2(new_n770_), .A3(new_n650_), .A4(new_n715_), .ZN(new_n771_));
  INV_X1    g570(.A(G57gat), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n772_), .A3(new_n469_), .ZN(new_n773_));
  NOR4_X1   g572(.A1(new_n665_), .A2(new_n770_), .A3(new_n668_), .A4(new_n650_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n774_), .A2(new_n469_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n773_), .B1(new_n775_), .B2(new_n772_), .ZN(G1332gat));
  INV_X1    g575(.A(G64gat), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n777_), .B1(new_n774_), .B2(new_n684_), .ZN(new_n778_));
  XOR2_X1   g577(.A(new_n778_), .B(KEYINPUT48), .Z(new_n779_));
  NAND3_X1  g578(.A1(new_n771_), .A2(new_n777_), .A3(new_n684_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(G1333gat));
  AOI21_X1  g580(.A(new_n435_), .B1(new_n774_), .B2(new_n659_), .ZN(new_n782_));
  XOR2_X1   g581(.A(new_n782_), .B(KEYINPUT49), .Z(new_n783_));
  NAND3_X1  g582(.A1(new_n771_), .A2(new_n435_), .A3(new_n659_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(G1334gat));
  INV_X1    g584(.A(G78gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n786_), .B1(new_n774_), .B2(new_n707_), .ZN(new_n787_));
  XOR2_X1   g586(.A(new_n787_), .B(KEYINPUT50), .Z(new_n788_));
  NAND3_X1  g587(.A1(new_n771_), .A2(new_n786_), .A3(new_n707_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(G1335gat));
  AND4_X1   g589(.A1(new_n484_), .A2(new_n671_), .A3(new_n670_), .A4(new_n731_), .ZN(new_n791_));
  INV_X1    g590(.A(G85gat), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n792_), .A3(new_n469_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n721_), .A2(new_n722_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n570_), .A2(new_n650_), .A3(new_n632_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT116), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n797_), .A2(new_n469_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n793_), .B1(new_n798_), .B2(new_n792_), .ZN(G1336gat));
  AOI21_X1  g598(.A(G92gat), .B1(new_n791_), .B2(new_n684_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n482_), .A2(new_n512_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n797_), .B2(new_n801_), .ZN(G1337gat));
  INV_X1    g601(.A(new_n511_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n791_), .A2(new_n659_), .A3(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT117), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n496_), .B1(new_n797_), .B2(new_n659_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  XOR2_X1   g606(.A(new_n807_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g607(.A1(new_n791_), .A2(new_n497_), .A3(new_n707_), .ZN(new_n809_));
  XOR2_X1   g608(.A(new_n809_), .B(KEYINPUT118), .Z(new_n810_));
  NAND3_X1  g609(.A1(new_n794_), .A2(new_n707_), .A3(new_n796_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(G106gat), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n811_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n810_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g616(.A1(new_n570_), .A2(new_n600_), .A3(new_n671_), .A4(new_n632_), .ZN(new_n818_));
  XOR2_X1   g617(.A(new_n818_), .B(KEYINPUT54), .Z(new_n819_));
  NAND2_X1  g618(.A1(new_n563_), .A2(new_n650_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT119), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n563_), .A2(new_n650_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n562_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n542_), .A2(new_n544_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n553_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT12), .B1(new_n548_), .B2(new_n533_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n827_), .A2(new_n555_), .A3(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n555_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(KEYINPUT55), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832_));
  NOR4_X1   g631(.A1(new_n827_), .A2(new_n828_), .A3(new_n832_), .A4(new_n555_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n825_), .B1(new_n831_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT56), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n551_), .B1(new_n545_), .B2(new_n550_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n552_), .B1(new_n837_), .B2(new_n832_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n833_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n562_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT56), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n824_), .B1(new_n836_), .B2(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n564_), .A2(new_n565_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n639_), .A2(new_n642_), .A3(new_n646_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n641_), .B1(new_n640_), .B2(new_n637_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n634_), .A2(new_n638_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(new_n641_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n844_), .B1(new_n847_), .B2(new_n646_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n843_), .A2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n666_), .B1(new_n842_), .B2(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n823_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n822_), .B1(new_n563_), .B2(new_n650_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n840_), .A2(KEYINPUT56), .ZN(new_n856_));
  AOI211_X1 g655(.A(new_n835_), .B(new_n562_), .C1(new_n838_), .C2(new_n839_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n855_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n849_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n851_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n666_), .A3(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n834_), .A2(KEYINPUT121), .A3(new_n835_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n864_), .B1(new_n840_), .B2(KEYINPUT56), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n863_), .A2(new_n865_), .A3(new_n841_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n564_), .A2(new_n848_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n866_), .A2(KEYINPUT58), .A3(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n715_), .ZN(new_n869_));
  AOI21_X1  g668(.A(KEYINPUT58), .B1(new_n866_), .B2(new_n867_), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n852_), .B(new_n862_), .C1(new_n869_), .C2(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n819_), .B1(new_n871_), .B2(new_n631_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n664_), .A2(new_n469_), .A3(new_n659_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(G113gat), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n874_), .A2(new_n875_), .A3(new_n650_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n874_), .A2(KEYINPUT59), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n878_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n671_), .B1(new_n877_), .B2(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n876_), .B1(new_n880_), .B2(new_n875_), .ZN(G1340gat));
  INV_X1    g680(.A(KEYINPUT60), .ZN(new_n882_));
  AOI21_X1  g681(.A(G120gat), .B1(new_n670_), .B2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(KEYINPUT122), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n885_), .B1(new_n882_), .B2(G120gat), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n874_), .B(new_n884_), .C1(new_n883_), .C2(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n570_), .B1(new_n877_), .B2(new_n879_), .ZN(new_n888_));
  INV_X1    g687(.A(G120gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n887_), .B1(new_n888_), .B2(new_n889_), .ZN(G1341gat));
  INV_X1    g689(.A(G127gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n874_), .A2(new_n891_), .A3(new_n632_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n631_), .B1(new_n877_), .B2(new_n879_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n891_), .ZN(G1342gat));
  INV_X1    g693(.A(G134gat), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n874_), .A2(new_n895_), .A3(new_n668_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n600_), .B1(new_n877_), .B2(new_n879_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n897_), .B2(new_n895_), .ZN(G1343gat));
  NOR2_X1   g697(.A1(new_n475_), .A2(new_n659_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n899_), .A2(new_n482_), .A3(new_n469_), .ZN(new_n900_));
  XOR2_X1   g699(.A(new_n900_), .B(KEYINPUT123), .Z(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(KEYINPUT124), .B1(new_n872_), .B2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT124), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n861_), .B1(new_n860_), .B2(new_n666_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n666_), .ZN(new_n906_));
  AOI211_X1 g705(.A(new_n906_), .B(new_n851_), .C1(new_n858_), .C2(new_n859_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n905_), .A2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n870_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n909_), .A2(new_n715_), .A3(new_n868_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n632_), .B1(new_n908_), .B2(new_n910_), .ZN(new_n911_));
  OAI211_X1 g710(.A(new_n904_), .B(new_n901_), .C1(new_n911_), .C2(new_n819_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n903_), .A2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n650_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(G141gat), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n913_), .A2(new_n331_), .A3(new_n650_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1344gat));
  NAND2_X1  g716(.A1(new_n913_), .A2(new_n670_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(KEYINPUT125), .B(G148gat), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n920_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n913_), .A2(new_n670_), .A3(new_n919_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1345gat));
  NAND2_X1  g722(.A1(new_n913_), .A2(new_n632_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(KEYINPUT61), .B(G155gat), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n925_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n913_), .A2(new_n632_), .A3(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n926_), .A2(new_n928_), .ZN(G1346gat));
  INV_X1    g728(.A(G162gat), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n913_), .A2(new_n930_), .A3(new_n668_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n600_), .B1(new_n903_), .B2(new_n912_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n930_), .B2(new_n932_), .ZN(G1347gat));
  NAND2_X1  g732(.A1(new_n871_), .A2(new_n631_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n819_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT126), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n482_), .A2(new_n469_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(new_n659_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n939_), .A2(new_n707_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n936_), .A2(new_n937_), .A3(new_n940_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n940_), .ZN(new_n942_));
  OAI21_X1  g741(.A(KEYINPUT126), .B1(new_n872_), .B2(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n941_), .A2(new_n943_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(KEYINPUT22), .B(G169gat), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n944_), .A2(new_n650_), .A3(new_n945_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n936_), .A2(new_n650_), .A3(new_n940_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n948_));
  AND3_X1   g747(.A1(new_n947_), .A2(new_n948_), .A3(G169gat), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n948_), .B1(new_n947_), .B2(G169gat), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n946_), .B1(new_n949_), .B2(new_n950_), .ZN(G1348gat));
  NAND3_X1  g750(.A1(new_n944_), .A2(new_n249_), .A3(new_n670_), .ZN(new_n952_));
  NOR3_X1   g751(.A1(new_n872_), .A2(new_n570_), .A3(new_n942_), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n952_), .B1(new_n249_), .B2(new_n953_), .ZN(G1349gat));
  NOR2_X1   g753(.A1(new_n872_), .A2(new_n942_), .ZN(new_n955_));
  AOI21_X1  g754(.A(G183gat), .B1(new_n955_), .B2(new_n632_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n631_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n956_), .B1(new_n944_), .B2(new_n957_), .ZN(G1350gat));
  INV_X1    g757(.A(new_n284_), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n944_), .A2(new_n959_), .A3(new_n668_), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n600_), .B1(new_n941_), .B2(new_n943_), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n960_), .B1(new_n239_), .B2(new_n961_), .ZN(G1351gat));
  NAND2_X1  g761(.A1(new_n899_), .A2(new_n938_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n872_), .A2(new_n963_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n964_), .A2(new_n650_), .ZN(new_n965_));
  XNOR2_X1  g764(.A(new_n965_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g765(.A1(new_n964_), .A2(new_n670_), .ZN(new_n967_));
  NOR2_X1   g766(.A1(new_n967_), .A2(new_n211_), .ZN(new_n968_));
  AOI21_X1  g767(.A(new_n968_), .B1(new_n217_), .B2(new_n967_), .ZN(G1353gat));
  INV_X1    g768(.A(new_n963_), .ZN(new_n970_));
  NAND3_X1  g769(.A1(new_n936_), .A2(new_n632_), .A3(new_n970_), .ZN(new_n971_));
  XOR2_X1   g770(.A(KEYINPUT63), .B(G211gat), .Z(new_n972_));
  INV_X1    g771(.A(new_n972_), .ZN(new_n973_));
  OAI21_X1  g772(.A(KEYINPUT127), .B1(new_n971_), .B2(new_n973_), .ZN(new_n974_));
  NOR2_X1   g773(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n971_), .A2(new_n975_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n974_), .A2(new_n976_), .ZN(new_n977_));
  NOR3_X1   g776(.A1(new_n971_), .A2(KEYINPUT127), .A3(new_n973_), .ZN(new_n978_));
  NOR2_X1   g777(.A1(new_n977_), .A2(new_n978_), .ZN(G1354gat));
  INV_X1    g778(.A(G218gat), .ZN(new_n980_));
  NAND3_X1  g779(.A1(new_n964_), .A2(new_n980_), .A3(new_n668_), .ZN(new_n981_));
  NOR3_X1   g780(.A1(new_n872_), .A2(new_n600_), .A3(new_n963_), .ZN(new_n982_));
  OAI21_X1  g781(.A(new_n981_), .B1(new_n982_), .B2(new_n980_), .ZN(G1355gat));
endmodule


