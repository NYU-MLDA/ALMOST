//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1 0 1 0 0 0 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n816_, new_n817_, new_n819_, new_n820_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n827_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n845_,
    new_n847_, new_n848_, new_n850_, new_n851_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_;
  XOR2_X1   g000(.A(G113gat), .B(G120gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G127gat), .B(G134gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n202_), .A2(new_n203_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT31), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n207_), .A2(KEYINPUT83), .ZN(new_n208_));
  INV_X1    g007(.A(G176gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT81), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n209_), .B1(new_n210_), .B2(KEYINPUT22), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G169gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT22), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n213_), .A2(KEYINPUT80), .ZN(new_n214_));
  INV_X1    g013(.A(G169gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n216_), .B(new_n210_), .C1(new_n214_), .C2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n219_), .B1(G183gat), .B2(G190gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(G183gat), .A3(G190gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT82), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n222_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n220_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n212_), .B(new_n218_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(G190gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n228_), .A2(KEYINPUT26), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n228_), .A2(KEYINPUT26), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT79), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n229_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT25), .B(G183gat), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n232_), .B(new_n233_), .C1(new_n231_), .C2(new_n230_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n220_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(new_n221_), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT24), .B1(new_n215_), .B2(new_n209_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n237_), .A2(new_n217_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n217_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n239_), .A2(KEYINPUT24), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n234_), .A2(new_n236_), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n227_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n208_), .B(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G227gat), .A2(G233gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(G71gat), .ZN(new_n246_));
  XOR2_X1   g045(.A(G15gat), .B(G43gat), .Z(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(KEYINPUT30), .B(G99gat), .Z(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n244_), .B(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT100), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G1gat), .B(G29gat), .ZN(new_n254_));
  INV_X1    g053(.A(G85gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT0), .B(G57gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(G155gat), .A2(G162gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT84), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G155gat), .A2(G162gat), .ZN(new_n261_));
  NOR2_X1   g060(.A1(G141gat), .A2(G148gat), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT3), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G141gat), .A2(G148gat), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT2), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n260_), .B(new_n261_), .C1(new_n264_), .C2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n262_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT84), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n259_), .B(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n261_), .B(KEYINPUT1), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n269_), .B(new_n265_), .C1(new_n271_), .C2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n268_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(new_n206_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n273_), .A2(new_n268_), .A3(new_n204_), .A4(new_n205_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(new_n276_), .A3(KEYINPUT4), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n274_), .A2(new_n278_), .A3(new_n206_), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G225gat), .A2(G233gat), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n275_), .A2(new_n276_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n281_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n258_), .B1(new_n282_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n282_), .A2(new_n286_), .A3(new_n258_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n253_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n282_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n258_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n286_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n291_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n294_), .A2(KEYINPUT100), .A3(new_n287_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n290_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT87), .ZN(new_n297_));
  INV_X1    g096(.A(G204gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(new_n298_), .A3(G197gat), .ZN(new_n299_));
  XOR2_X1   g098(.A(G197gat), .B(G204gat), .Z(new_n300_));
  OAI211_X1 g099(.A(KEYINPUT21), .B(new_n299_), .C1(new_n300_), .C2(new_n297_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT88), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n302_), .B1(new_n300_), .B2(KEYINPUT21), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT89), .ZN(new_n304_));
  AND2_X1   g103(.A1(G211gat), .A2(G218gat), .ZN(new_n305_));
  NOR2_X1   g104(.A1(G211gat), .A2(G218gat), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n304_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(G211gat), .ZN(new_n308_));
  INV_X1    g107(.A(G218gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G211gat), .A2(G218gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(KEYINPUT89), .A3(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n307_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G197gat), .B(G204gat), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT21), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(KEYINPUT88), .A3(new_n315_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n301_), .A2(new_n303_), .A3(new_n313_), .A4(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT90), .ZN(new_n318_));
  NOR3_X1   g117(.A1(new_n305_), .A2(new_n306_), .A3(new_n304_), .ZN(new_n319_));
  AOI21_X1  g118(.A(KEYINPUT89), .B1(new_n310_), .B2(new_n311_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n318_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n307_), .A2(new_n312_), .A3(KEYINPUT90), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n321_), .A2(KEYINPUT21), .A3(new_n322_), .A4(new_n300_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n323_), .A2(KEYINPUT91), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT91), .ZN(new_n325_));
  AND2_X1   g124(.A1(new_n322_), .A2(new_n300_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n315_), .B1(new_n313_), .B2(new_n318_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n325_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n317_), .B1(new_n324_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n274_), .A2(KEYINPUT29), .ZN(new_n330_));
  INV_X1    g129(.A(G233gat), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n331_), .A2(KEYINPUT86), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n331_), .A2(KEYINPUT86), .ZN(new_n333_));
  OAI21_X1  g132(.A(G228gat), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n329_), .A2(new_n330_), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n334_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n317_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n323_), .A2(KEYINPUT91), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n326_), .A2(new_n325_), .A3(new_n327_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n337_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n330_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n336_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  XOR2_X1   g141(.A(G78gat), .B(G106gat), .Z(new_n343_));
  NAND3_X1  g142(.A1(new_n335_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(G22gat), .B(G50gat), .Z(new_n345_));
  OAI21_X1  g144(.A(new_n345_), .B1(new_n274_), .B2(KEYINPUT29), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT29), .ZN(new_n347_));
  INV_X1    g146(.A(new_n345_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n273_), .A2(new_n268_), .A3(new_n347_), .A4(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n346_), .A2(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n350_), .B(new_n352_), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n344_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n343_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n334_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n356_));
  NOR3_X1   g155(.A1(new_n340_), .A2(new_n341_), .A3(new_n336_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n355_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT92), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT92), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n360_), .B(new_n355_), .C1(new_n356_), .C2(new_n357_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n354_), .A2(new_n359_), .A3(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT93), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT93), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n354_), .A2(new_n359_), .A3(new_n364_), .A4(new_n361_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n358_), .A2(new_n344_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n353_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n296_), .B1(new_n366_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n243_), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT96), .B1(new_n340_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT96), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n329_), .A2(new_n373_), .A3(new_n243_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT20), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n226_), .B1(new_n235_), .B2(new_n221_), .ZN(new_n376_));
  XOR2_X1   g175(.A(KEYINPUT22), .B(G169gat), .Z(new_n377_));
  NOR2_X1   g176(.A1(new_n377_), .A2(G176gat), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n215_), .A2(new_n209_), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n376_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT94), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n233_), .B(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n230_), .A2(new_n229_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n225_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n237_), .B(KEYINPUT95), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n240_), .B1(new_n385_), .B2(new_n239_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n380_), .B1(new_n384_), .B2(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n375_), .B1(new_n340_), .B2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G226gat), .A2(G233gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT19), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n372_), .A2(new_n374_), .A3(new_n388_), .A4(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT97), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n387_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n375_), .B1(new_n329_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n340_), .A2(new_n371_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n391_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n392_), .B1(new_n398_), .B2(new_n393_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G8gat), .B(G36gat), .ZN(new_n400_));
  INV_X1    g199(.A(G92gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT18), .B(G64gat), .ZN(new_n403_));
  XOR2_X1   g202(.A(new_n402_), .B(new_n403_), .Z(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n394_), .A2(new_n399_), .A3(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n372_), .A2(new_n374_), .A3(new_n388_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT99), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n407_), .A2(new_n408_), .A3(new_n390_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n408_), .B1(new_n407_), .B2(new_n390_), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n396_), .A2(new_n391_), .A3(new_n397_), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n409_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  OAI211_X1 g211(.A(KEYINPUT27), .B(new_n406_), .C1(new_n412_), .C2(new_n405_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT101), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n394_), .A2(new_n399_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n404_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n406_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT27), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n407_), .A2(new_n390_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT99), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n407_), .A2(new_n408_), .A3(new_n390_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n404_), .B1(new_n423_), .B2(new_n411_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT101), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n424_), .A2(new_n425_), .A3(KEYINPUT27), .A4(new_n406_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n370_), .A2(new_n414_), .A3(new_n419_), .A4(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n294_), .A2(new_n287_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n405_), .A2(KEYINPUT32), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n394_), .A2(new_n399_), .A3(new_n429_), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n428_), .B(new_n430_), .C1(new_n412_), .C2(new_n429_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n292_), .B1(new_n283_), .B2(new_n281_), .ZN(new_n432_));
  XOR2_X1   g231(.A(new_n432_), .B(KEYINPUT98), .Z(new_n433_));
  NAND2_X1  g232(.A1(new_n280_), .A2(new_n281_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n416_), .A2(new_n406_), .A3(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(new_n287_), .B(KEYINPUT33), .Z(new_n437_));
  OAI21_X1  g236(.A(new_n431_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n363_), .A2(new_n365_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n252_), .B1(new_n427_), .B2(new_n440_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n414_), .A2(new_n419_), .A3(new_n426_), .A4(new_n439_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n296_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n252_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n441_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT78), .ZN(new_n447_));
  XNOR2_X1  g246(.A(KEYINPUT72), .B(G8gat), .ZN(new_n448_));
  INV_X1    g247(.A(G1gat), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT14), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT73), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G15gat), .B(G22gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  XOR2_X1   g253(.A(G1gat), .B(G8gat), .Z(new_n455_));
  OR2_X1    g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n455_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G29gat), .B(G36gat), .ZN(new_n460_));
  INV_X1    g259(.A(G50gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT69), .B(G43gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n459_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n464_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n458_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G229gat), .A2(G233gat), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(G169gat), .B(G197gat), .Z(new_n472_));
  XNOR2_X1  g271(.A(G113gat), .B(G141gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT77), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT76), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT15), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n464_), .B(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n459_), .A2(new_n478_), .A3(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n464_), .B(KEYINPUT15), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT76), .B1(new_n458_), .B2(new_n482_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n481_), .A2(new_n483_), .A3(new_n469_), .A4(new_n467_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n471_), .A2(new_n477_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n477_), .B1(new_n471_), .B2(new_n484_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n447_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n487_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n489_), .A2(KEYINPUT78), .A3(new_n485_), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n446_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT10), .B(G99gat), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n493_), .A2(G106gat), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT65), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G99gat), .A2(G106gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT6), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G85gat), .B(G92gat), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT9), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT9), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n502_), .A2(G85gat), .A3(G92gat), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n496_), .A2(new_n498_), .A3(new_n501_), .A4(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT8), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n498_), .A2(KEYINPUT66), .ZN(new_n506_));
  NOR2_X1   g305(.A1(G99gat), .A2(G106gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT7), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n498_), .A2(KEYINPUT66), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n506_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n505_), .B1(new_n510_), .B2(new_n500_), .ZN(new_n511_));
  AOI211_X1 g310(.A(KEYINPUT8), .B(new_n499_), .C1(new_n508_), .C2(new_n498_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n504_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(KEYINPUT67), .B(G71gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(G78gat), .ZN(new_n515_));
  XOR2_X1   g314(.A(G57gat), .B(G64gat), .Z(new_n516_));
  INV_X1    g315(.A(KEYINPUT11), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n516_), .A2(new_n517_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n515_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(G78gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n514_), .B(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n518_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n513_), .A2(new_n526_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n525_), .B(new_n504_), .C1(new_n511_), .C2(new_n512_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n527_), .A2(KEYINPUT12), .A3(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT12), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n513_), .A2(new_n530_), .A3(new_n526_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G230gat), .A2(G233gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT64), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(new_n534_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n527_), .A2(new_n528_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n535_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(KEYINPUT5), .B(G176gat), .Z(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT68), .B(G204gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G120gat), .B(G148gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n537_), .B(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT13), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n492_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT37), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G232gat), .A2(G233gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT34), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n549_), .A2(KEYINPUT35), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n480_), .A2(new_n513_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT70), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n552_), .A2(KEYINPUT35), .A3(new_n549_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n513_), .A2(new_n464_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n551_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n555_), .A2(new_n552_), .A3(KEYINPUT35), .A4(new_n549_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n550_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G190gat), .B(G218gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(G162gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(KEYINPUT71), .B(G134gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT36), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n563_), .A2(new_n564_), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n559_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n565_), .B1(new_n559_), .B2(new_n566_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n547_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G231gat), .A2(G233gat), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n525_), .B(new_n570_), .Z(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(new_n458_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT17), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  XOR2_X1   g373(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n575_));
  XNOR2_X1  g374(.A(G127gat), .B(G155gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G183gat), .B(G211gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  MUX2_X1   g378(.A(new_n574_), .B(new_n573_), .S(new_n579_), .Z(new_n580_));
  INV_X1    g379(.A(KEYINPUT75), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n572_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n580_), .B(new_n582_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n557_), .A2(new_n558_), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n564_), .B(new_n563_), .C1(new_n584_), .C2(new_n550_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n559_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(KEYINPUT37), .A3(new_n586_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n569_), .A2(new_n583_), .A3(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n546_), .A2(new_n588_), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n589_), .A2(G1gat), .A3(new_n443_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n590_), .A2(KEYINPUT38), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT102), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n567_), .A2(new_n568_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n446_), .A2(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n543_), .B(KEYINPUT13), .Z(new_n595_));
  NAND2_X1  g394(.A1(new_n489_), .A2(new_n485_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n594_), .A2(new_n583_), .A3(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n449_), .B1(new_n599_), .B2(new_n296_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n600_), .B1(new_n590_), .B2(KEYINPUT38), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n592_), .A2(new_n601_), .ZN(G1324gat));
  INV_X1    g401(.A(G8gat), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n414_), .A2(new_n419_), .A3(new_n426_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n603_), .B1(new_n599_), .B2(new_n604_), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n605_), .B(KEYINPUT39), .Z(new_n606_));
  INV_X1    g405(.A(new_n589_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n607_), .A2(new_n448_), .A3(new_n604_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT40), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(G1325gat));
  INV_X1    g410(.A(G15gat), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n612_), .B1(new_n599_), .B2(new_n252_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT41), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n607_), .A2(new_n612_), .A3(new_n252_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT103), .ZN(G1326gat));
  INV_X1    g416(.A(G22gat), .ZN(new_n618_));
  INV_X1    g417(.A(new_n439_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n618_), .B1(new_n599_), .B2(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT42), .Z(new_n621_));
  NOR2_X1   g420(.A1(new_n439_), .A2(G22gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT104), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n621_), .B1(new_n589_), .B2(new_n623_), .ZN(G1327gat));
  NAND2_X1  g423(.A1(new_n427_), .A2(new_n440_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(new_n251_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n445_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT105), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT43), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n569_), .A2(new_n587_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n628_), .A2(new_n629_), .A3(new_n630_), .A4(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n631_), .ZN(new_n633_));
  OAI21_X1  g432(.A(KEYINPUT43), .B1(new_n446_), .B2(new_n633_), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n630_), .B(new_n631_), .C1(new_n441_), .C2(new_n445_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT105), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n632_), .A2(new_n634_), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n583_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(new_n638_), .A3(new_n598_), .ZN(new_n639_));
  XOR2_X1   g438(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n637_), .A2(KEYINPUT44), .A3(new_n638_), .A4(new_n598_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OAI211_X1 g442(.A(KEYINPUT107), .B(G29gat), .C1(new_n643_), .C2(new_n443_), .ZN(new_n644_));
  INV_X1    g443(.A(G29gat), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n643_), .A2(KEYINPUT107), .A3(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n593_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n545_), .A2(new_n583_), .A3(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n646_), .B1(new_n645_), .B2(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n644_), .B1(new_n649_), .B2(new_n443_), .ZN(G1328gat));
  INV_X1    g449(.A(new_n604_), .ZN(new_n651_));
  OAI21_X1  g450(.A(G36gat), .B1(new_n643_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(G36gat), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n648_), .A2(new_n653_), .A3(new_n604_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT45), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n652_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT46), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(new_n657_), .ZN(G1329gat));
  OAI21_X1  g457(.A(G43gat), .B1(new_n643_), .B2(new_n251_), .ZN(new_n659_));
  INV_X1    g458(.A(G43gat), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n648_), .A2(new_n660_), .A3(new_n252_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT47), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(G1330gat));
  NAND3_X1  g463(.A1(new_n648_), .A2(new_n461_), .A3(new_n619_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n641_), .A2(new_n619_), .A3(new_n642_), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n666_), .A2(KEYINPUT108), .A3(G50gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(KEYINPUT108), .B1(new_n666_), .B2(G50gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n665_), .B1(new_n667_), .B2(new_n668_), .ZN(G1331gat));
  NAND4_X1  g468(.A1(new_n594_), .A2(new_n583_), .A3(new_n595_), .A4(new_n491_), .ZN(new_n670_));
  INV_X1    g469(.A(G57gat), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n670_), .A2(new_n671_), .A3(new_n443_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT110), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n446_), .A2(new_n596_), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n674_), .A2(KEYINPUT109), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(KEYINPUT109), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n675_), .A2(new_n588_), .A3(new_n595_), .A4(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n671_), .B1(new_n677_), .B2(new_n443_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n673_), .A2(new_n678_), .ZN(G1332gat));
  OAI21_X1  g478(.A(G64gat), .B1(new_n670_), .B2(new_n651_), .ZN(new_n680_));
  XOR2_X1   g479(.A(KEYINPUT111), .B(KEYINPUT48), .Z(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n651_), .A2(G64gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n682_), .B1(new_n677_), .B2(new_n683_), .ZN(G1333gat));
  OAI21_X1  g483(.A(G71gat), .B1(new_n670_), .B2(new_n251_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT49), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n251_), .A2(G71gat), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n686_), .B1(new_n677_), .B2(new_n687_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT112), .ZN(G1334gat));
  OAI21_X1  g488(.A(G78gat), .B1(new_n670_), .B2(new_n439_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT50), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n619_), .A2(new_n522_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(new_n677_), .B2(new_n692_), .ZN(G1335gat));
  NOR2_X1   g492(.A1(new_n647_), .A2(new_n583_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n675_), .A2(new_n595_), .A3(new_n694_), .A4(new_n676_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n255_), .B1(new_n695_), .B2(new_n443_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n544_), .A2(new_n583_), .A3(new_n596_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n637_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n698_), .A2(G85gat), .A3(new_n296_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n696_), .A2(new_n699_), .ZN(G1336gat));
  OAI21_X1  g499(.A(new_n401_), .B1(new_n695_), .B2(new_n651_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n698_), .A2(G92gat), .A3(new_n604_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1337gat));
  OR2_X1    g502(.A1(new_n251_), .A2(new_n493_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n695_), .A2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n698_), .A2(new_n252_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(G99gat), .B2(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT114), .Z(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n709_), .B(new_n712_), .ZN(G1338gat));
  NAND3_X1  g512(.A1(new_n637_), .A2(new_n619_), .A3(new_n697_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT115), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n637_), .A2(KEYINPUT115), .A3(new_n619_), .A4(new_n697_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n716_), .A2(G106gat), .A3(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT52), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT52), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n716_), .A2(new_n720_), .A3(G106gat), .A4(new_n717_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(new_n722_));
  OR3_X1    g521(.A1(new_n695_), .A2(G106gat), .A3(new_n439_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT53), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT53), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n722_), .A2(new_n726_), .A3(new_n723_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1339gat));
  NAND4_X1  g527(.A1(new_n651_), .A2(new_n296_), .A3(new_n439_), .A4(new_n252_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n481_), .A2(new_n483_), .A3(new_n467_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(new_n470_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n465_), .A2(new_n469_), .A3(new_n467_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n474_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n471_), .A2(new_n484_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n733_), .B1(new_n474_), .B2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(new_n543_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n534_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n529_), .A2(new_n738_), .A3(new_n531_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n535_), .A2(KEYINPUT55), .A3(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT55), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n532_), .A2(new_n741_), .A3(new_n534_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n740_), .A2(new_n542_), .A3(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT56), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n740_), .A2(KEYINPUT56), .A3(new_n542_), .A4(new_n742_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT116), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n596_), .B1(new_n745_), .B2(new_n748_), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n537_), .A2(new_n542_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n743_), .A2(new_n744_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n751_), .B2(new_n747_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n737_), .B1(new_n749_), .B2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(new_n647_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT57), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n753_), .A2(KEYINPUT57), .A3(new_n647_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT117), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n751_), .A2(new_n759_), .A3(new_n746_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n743_), .A2(KEYINPUT117), .A3(new_n744_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n760_), .A2(new_n750_), .A3(new_n736_), .A4(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT118), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT58), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n762_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n765_), .A2(new_n766_), .A3(new_n633_), .ZN(new_n767_));
  OAI21_X1  g566(.A(KEYINPUT119), .B1(new_n758_), .B2(new_n767_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n753_), .A2(KEYINPUT57), .A3(new_n647_), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT57), .B1(new_n753_), .B2(new_n647_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT119), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n762_), .A2(new_n763_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT58), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n762_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(new_n631_), .A3(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n771_), .A2(new_n772_), .A3(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n768_), .A2(new_n777_), .A3(new_n638_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT54), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n588_), .A2(new_n779_), .A3(new_n544_), .A4(new_n491_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n569_), .A2(new_n491_), .A3(new_n583_), .A4(new_n587_), .ZN(new_n781_));
  OAI21_X1  g580(.A(KEYINPUT54), .B1(new_n781_), .B2(new_n595_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n780_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n729_), .B1(new_n778_), .B2(new_n784_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT120), .ZN(new_n786_));
  AOI21_X1  g585(.A(G113gat), .B1(new_n786_), .B2(new_n596_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n729_), .B(KEYINPUT122), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n638_), .B1(new_n758_), .B2(new_n767_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(new_n789_), .B2(new_n784_), .ZN(new_n790_));
  XOR2_X1   g589(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT123), .B1(new_n790_), .B2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n776_), .A2(new_n756_), .A3(new_n757_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n783_), .B1(new_n794_), .B2(new_n638_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT123), .ZN(new_n796_));
  NOR4_X1   g595(.A1(new_n795_), .A2(new_n796_), .A3(new_n791_), .A4(new_n788_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT59), .ZN(new_n798_));
  OAI22_X1  g597(.A1(new_n793_), .A2(new_n797_), .B1(new_n785_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT124), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n788_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n583_), .B1(new_n771_), .B2(new_n776_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n792_), .B(new_n802_), .C1(new_n803_), .C2(new_n783_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n796_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n790_), .A2(KEYINPUT123), .A3(new_n792_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n807_), .B(KEYINPUT124), .C1(new_n798_), .C2(new_n785_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n491_), .B1(new_n801_), .B2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n787_), .B1(new_n809_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g609(.A(G120gat), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n544_), .B2(KEYINPUT60), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n786_), .B(new_n812_), .C1(KEYINPUT60), .C2(new_n811_), .ZN(new_n813_));
  OAI21_X1  g612(.A(G120gat), .B1(new_n799_), .B2(new_n544_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(G1341gat));
  AOI21_X1  g614(.A(G127gat), .B1(new_n786_), .B2(new_n583_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n638_), .B1(new_n801_), .B2(new_n808_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n816_), .B1(new_n817_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g617(.A(G134gat), .B1(new_n786_), .B2(new_n593_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n633_), .B1(new_n801_), .B2(new_n808_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n820_), .B2(G134gat), .ZN(G1343gat));
  AOI21_X1  g620(.A(new_n252_), .B1(new_n778_), .B2(new_n784_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n822_), .A2(new_n619_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n604_), .A2(new_n443_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n596_), .A3(new_n824_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g625(.A1(new_n823_), .A2(new_n595_), .A3(new_n824_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g627(.A1(new_n823_), .A2(new_n583_), .A3(new_n824_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(KEYINPUT61), .B(G155gat), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n829_), .B(new_n830_), .ZN(G1346gat));
  AND4_X1   g630(.A1(G162gat), .A2(new_n823_), .A3(new_n631_), .A4(new_n824_), .ZN(new_n832_));
  INV_X1    g631(.A(G162gat), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n823_), .A2(new_n593_), .A3(new_n824_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n832_), .B1(new_n833_), .B2(new_n834_), .ZN(G1347gat));
  NAND4_X1  g634(.A1(new_n604_), .A2(new_n443_), .A3(new_n439_), .A4(new_n252_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n795_), .A2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n596_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(G169gat), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(KEYINPUT62), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n377_), .B2(new_n838_), .ZN(G1348gat));
  NAND3_X1  g640(.A1(new_n837_), .A2(new_n209_), .A3(new_n595_), .ZN(new_n842_));
  AOI211_X1 g641(.A(new_n544_), .B(new_n836_), .C1(new_n778_), .C2(new_n784_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n209_), .ZN(G1349gat));
  NAND2_X1  g643(.A1(new_n837_), .A2(new_n583_), .ZN(new_n845_));
  MUX2_X1   g644(.A(new_n382_), .B(G183gat), .S(new_n845_), .Z(G1350gat));
  NAND3_X1  g645(.A1(new_n837_), .A2(new_n593_), .A3(new_n383_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n795_), .A2(new_n633_), .A3(new_n836_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n228_), .B2(new_n848_), .ZN(G1351gat));
  NAND3_X1  g648(.A1(new_n822_), .A2(new_n370_), .A3(new_n604_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n850_), .A2(new_n597_), .ZN(new_n851_));
  XOR2_X1   g650(.A(new_n851_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g651(.A1(new_n850_), .A2(new_n544_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(new_n298_), .ZN(G1353gat));
  NAND2_X1  g653(.A1(new_n619_), .A2(new_n443_), .ZN(new_n855_));
  AOI211_X1 g654(.A(new_n855_), .B(new_n252_), .C1(new_n778_), .C2(new_n784_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n638_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n856_), .A2(new_n604_), .A3(new_n857_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(KEYINPUT125), .B(KEYINPUT126), .ZN(new_n859_));
  NOR2_X1   g658(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n859_), .B(new_n860_), .ZN(new_n861_));
  XOR2_X1   g660(.A(new_n858_), .B(new_n861_), .Z(G1354gat));
  NOR3_X1   g661(.A1(new_n850_), .A2(new_n309_), .A3(new_n633_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT127), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n864_), .B1(new_n850_), .B2(new_n647_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n856_), .A2(KEYINPUT127), .A3(new_n593_), .A4(new_n604_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n863_), .B1(new_n867_), .B2(new_n309_), .ZN(G1355gat));
endmodule


