//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n812_, new_n813_,
    new_n815_, new_n816_, new_n818_, new_n819_, new_n820_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n861_, new_n862_, new_n863_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  INV_X1    g001(.A(G43gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G50gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n202_), .B(G43gat), .ZN(new_n206_));
  INV_X1    g005(.A(G50gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n205_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT15), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n205_), .A2(new_n208_), .A3(KEYINPUT15), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT9), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n216_), .A2(KEYINPUT65), .ZN(new_n217_));
  INV_X1    g016(.A(G85gat), .ZN(new_n218_));
  INV_X1    g017(.A(G92gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n216_), .A2(KEYINPUT65), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n217_), .A2(new_n220_), .A3(new_n221_), .A4(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G99gat), .A2(G106gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT6), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT6), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(G99gat), .A3(G106gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT10), .B(G99gat), .ZN(new_n229_));
  OR3_X1    g028(.A1(new_n229_), .A2(KEYINPUT64), .A3(G106gat), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT64), .B1(new_n229_), .B2(G106gat), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n223_), .A2(new_n228_), .A3(new_n230_), .A4(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT8), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n220_), .A2(new_n214_), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n225_), .A2(new_n227_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT7), .ZN(new_n236_));
  INV_X1    g035(.A(G99gat), .ZN(new_n237_));
  INV_X1    g036(.A(G106gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n233_), .B(new_n234_), .C1(new_n235_), .C2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT66), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n228_), .A2(new_n240_), .A3(new_n239_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n244_), .A2(new_n245_), .A3(new_n233_), .A4(new_n234_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n228_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n225_), .A2(new_n227_), .A3(KEYINPUT67), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n249_), .A2(new_n240_), .A3(new_n239_), .A4(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n233_), .B1(new_n251_), .B2(new_n234_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n232_), .B1(new_n247_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n213_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT74), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT74), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n213_), .A2(new_n256_), .A3(new_n253_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT75), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n255_), .A2(KEYINPUT75), .A3(new_n257_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G232gat), .A2(G233gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT34), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n263_), .A2(KEYINPUT35), .ZN(new_n264_));
  INV_X1    g063(.A(new_n253_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n209_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n264_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n260_), .A2(new_n261_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n263_), .A2(KEYINPUT35), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n269_), .B(KEYINPUT73), .Z(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n268_), .A2(KEYINPUT76), .A3(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(KEYINPUT76), .B1(new_n268_), .B2(new_n271_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT36), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G190gat), .B(G218gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(G134gat), .ZN(new_n278_));
  INV_X1    g077(.A(G162gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n258_), .A2(new_n270_), .A3(new_n267_), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n275_), .A2(new_n276_), .A3(new_n280_), .A4(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n268_), .A2(new_n271_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT76), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n285_), .A2(new_n281_), .A3(new_n272_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n280_), .A2(new_n276_), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n280_), .A2(new_n276_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n286_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT77), .B(KEYINPUT37), .ZN(new_n290_));
  AND3_X1   g089(.A1(new_n282_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(KEYINPUT77), .A2(KEYINPUT37), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n292_), .B1(new_n282_), .B2(new_n289_), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G127gat), .B(G155gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT16), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G183gat), .B(G211gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT79), .B(KEYINPUT80), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n300_), .A2(new_n301_), .A3(KEYINPUT17), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G57gat), .B(G64gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT11), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G71gat), .B(G78gat), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n303_), .A2(KEYINPUT11), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n304_), .A2(new_n305_), .ZN(new_n308_));
  AND3_X1   g107(.A1(new_n306_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G231gat), .A2(G233gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G1gat), .B(G8gat), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n312_), .A2(KEYINPUT78), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(KEYINPUT78), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G15gat), .B(G22gat), .ZN(new_n316_));
  INV_X1    g115(.A(G1gat), .ZN(new_n317_));
  INV_X1    g116(.A(G8gat), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT14), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n315_), .A2(new_n320_), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n313_), .A2(new_n319_), .A3(new_n316_), .A4(new_n314_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n311_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n300_), .A2(KEYINPUT17), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n302_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n327_), .B1(new_n302_), .B2(new_n325_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n294_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT81), .ZN(new_n330_));
  XOR2_X1   g129(.A(G78gat), .B(G106gat), .Z(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G22gat), .B(G50gat), .ZN(new_n333_));
  OR2_X1    g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT89), .ZN(new_n336_));
  INV_X1    g135(.A(G141gat), .ZN(new_n337_));
  INV_X1    g136(.A(G148gat), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n336_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT2), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n337_), .A2(new_n338_), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT87), .B1(new_n341_), .B2(KEYINPUT3), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT87), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n343_), .A2(new_n344_), .A3(new_n337_), .A4(new_n338_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT2), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n336_), .B(new_n346_), .C1(new_n337_), .C2(new_n338_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n340_), .A2(new_n342_), .A3(new_n345_), .A4(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT88), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n334_), .B(new_n335_), .C1(new_n348_), .C2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n341_), .B(KEYINPUT85), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT86), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n353_), .B1(new_n335_), .B2(KEYINPUT1), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n335_), .A2(KEYINPUT1), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT1), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n356_), .A2(KEYINPUT86), .A3(G155gat), .A4(G162gat), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n354_), .A2(new_n355_), .A3(new_n334_), .A4(new_n357_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n352_), .B(new_n358_), .C1(new_n337_), .C2(new_n338_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n351_), .A2(new_n359_), .ZN(new_n360_));
  OR3_X1    g159(.A1(new_n360_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT90), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT28), .B1(new_n360_), .B2(KEYINPUT29), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n361_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n362_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n333_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n366_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n333_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n369_), .A3(new_n364_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n367_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT96), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n360_), .A2(KEYINPUT29), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT91), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G197gat), .A2(G204gat), .ZN(new_n376_));
  XOR2_X1   g175(.A(KEYINPUT92), .B(G197gat), .Z(new_n377_));
  OAI211_X1 g176(.A(KEYINPUT21), .B(new_n376_), .C1(new_n377_), .C2(G204gat), .ZN(new_n378_));
  XOR2_X1   g177(.A(G211gat), .B(G218gat), .Z(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(G204gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(G197gat), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n382_), .B1(new_n377_), .B2(new_n381_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n378_), .B(new_n380_), .C1(new_n383_), .C2(KEYINPUT21), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(KEYINPUT21), .A3(new_n379_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT93), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n384_), .A2(KEYINPUT93), .A3(new_n385_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  AND2_X1   g189(.A1(G228gat), .A2(G233gat), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n360_), .A2(KEYINPUT91), .A3(KEYINPUT29), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n375_), .A2(new_n390_), .A3(new_n392_), .A4(new_n393_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n373_), .A2(KEYINPUT94), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n386_), .B(KEYINPUT95), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n373_), .A2(KEYINPUT94), .ZN(new_n397_));
  NOR3_X1   g196(.A1(new_n395_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n372_), .B(new_n394_), .C1(new_n398_), .C2(new_n392_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n371_), .A2(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n394_), .B1(new_n398_), .B2(new_n392_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT96), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n402_), .A2(new_n399_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n332_), .B(new_n400_), .C1(new_n403_), .C2(new_n371_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n371_), .B1(new_n402_), .B2(new_n399_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n400_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n331_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n404_), .A2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G8gat), .B(G36gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT18), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(G64gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(new_n219_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT20), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G183gat), .A2(G190gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT23), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n415_), .B1(new_n416_), .B2(new_n414_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n417_), .B1(G183gat), .B2(G190gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G169gat), .A2(G176gat), .ZN(new_n419_));
  INV_X1    g218(.A(G176gat), .ZN(new_n420_));
  INV_X1    g219(.A(G169gat), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT84), .B1(new_n421_), .B2(KEYINPUT22), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT22), .B(G169gat), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n420_), .B(new_n422_), .C1(new_n423_), .C2(KEYINPUT84), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n418_), .A2(new_n419_), .A3(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(G169gat), .A2(G176gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT82), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(KEYINPUT24), .A3(new_n419_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n414_), .A2(KEYINPUT23), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n429_), .B1(new_n416_), .B2(new_n414_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT82), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n426_), .B(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT24), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT26), .B(G190gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT25), .B(G183gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n428_), .A2(new_n431_), .A3(new_n435_), .A4(new_n438_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n425_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n413_), .B1(new_n390_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G226gat), .A2(G233gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT19), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n437_), .B(KEYINPUT97), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n436_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n426_), .A2(new_n434_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n447_), .A2(new_n428_), .A3(new_n417_), .A4(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n423_), .A2(new_n420_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(G183gat), .A2(G190gat), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n450_), .B(new_n419_), .C1(new_n430_), .C2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n449_), .A2(new_n452_), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n442_), .B(new_n445_), .C1(new_n386_), .C2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n388_), .A2(new_n389_), .A3(new_n440_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n386_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n456_), .A3(KEYINPUT20), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n444_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n458_), .A2(KEYINPUT98), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT98), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n460_), .B1(new_n457_), .B2(new_n444_), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n412_), .B(new_n454_), .C1(new_n459_), .C2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n449_), .A2(KEYINPUT102), .A3(new_n452_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT102), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n453_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n396_), .A2(new_n463_), .A3(new_n465_), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n466_), .A2(new_n442_), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT103), .B1(new_n467_), .B2(new_n445_), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n457_), .A2(new_n444_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n466_), .A2(new_n442_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT103), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(new_n471_), .A3(new_n444_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n468_), .A2(new_n469_), .A3(new_n472_), .ZN(new_n473_));
  OAI211_X1 g272(.A(KEYINPUT27), .B(new_n462_), .C1(new_n473_), .C2(new_n412_), .ZN(new_n474_));
  XOR2_X1   g273(.A(KEYINPUT106), .B(KEYINPUT27), .Z(new_n475_));
  XNOR2_X1  g274(.A(new_n458_), .B(KEYINPUT98), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n412_), .B1(new_n476_), .B2(new_n454_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n462_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n475_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n474_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G127gat), .B(G134gat), .ZN(new_n481_));
  INV_X1    g280(.A(G113gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(G120gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n440_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G15gat), .B(G43gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT31), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n485_), .B(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G71gat), .B(G99gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT30), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G227gat), .A2(G233gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n488_), .B(new_n492_), .Z(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NOR3_X1   g293(.A1(new_n408_), .A2(new_n480_), .A3(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n484_), .B(new_n360_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G225gat), .A2(G233gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT4), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n484_), .A2(new_n360_), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n498_), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n501_), .B(new_n502_), .C1(new_n496_), .C2(new_n500_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n499_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G1gat), .B(G29gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(G85gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT0), .ZN(new_n507_));
  INV_X1    g306(.A(G57gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n504_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT104), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n499_), .A2(new_n503_), .A3(new_n509_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n504_), .A2(KEYINPUT104), .A3(new_n510_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n495_), .A2(new_n517_), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n404_), .A2(new_n407_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n519_), .A2(new_n480_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n468_), .A2(new_n472_), .A3(new_n469_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n412_), .A2(KEYINPUT32), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n476_), .A2(new_n522_), .A3(new_n454_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n524_), .A2(new_n516_), .A3(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT105), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n477_), .A2(new_n478_), .ZN(new_n528_));
  XOR2_X1   g327(.A(KEYINPUT100), .B(KEYINPUT33), .Z(new_n529_));
  AOI21_X1  g328(.A(KEYINPUT101), .B1(new_n514_), .B2(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n501_), .B1(new_n496_), .B2(new_n500_), .ZN(new_n531_));
  MUX2_X1   g330(.A(new_n496_), .B(new_n531_), .S(new_n498_), .Z(new_n532_));
  AOI21_X1  g331(.A(new_n530_), .B1(new_n510_), .B2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n514_), .A2(KEYINPUT101), .A3(new_n529_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n499_), .A2(new_n503_), .A3(KEYINPUT33), .A4(new_n509_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT99), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n528_), .A2(new_n533_), .A3(new_n534_), .A4(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT105), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n524_), .A2(new_n516_), .A3(new_n538_), .A4(new_n525_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n527_), .A2(new_n537_), .A3(new_n539_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n520_), .A2(new_n517_), .B1(new_n540_), .B2(new_n519_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n518_), .B1(new_n541_), .B2(new_n493_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n330_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n323_), .A2(new_n209_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n544_), .B1(new_n213_), .B2(new_n323_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G229gat), .A2(G233gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n323_), .B(new_n209_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n548_), .A2(G229gat), .A3(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G113gat), .B(G141gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(new_n421_), .ZN(new_n551_));
  INV_X1    g350(.A(G197gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n547_), .A2(new_n549_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n554_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT13), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n309_), .B(new_n232_), .C1(new_n247_), .C2(new_n252_), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n561_), .A2(KEYINPUT68), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(KEYINPUT68), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n309_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n253_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT69), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G230gat), .A2(G233gat), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n567_), .A2(new_n568_), .A3(new_n570_), .ZN(new_n571_));
  AOI22_X1  g370(.A1(new_n562_), .A2(new_n563_), .B1(new_n565_), .B2(new_n253_), .ZN(new_n572_));
  OAI21_X1  g371(.A(KEYINPUT69), .B1(new_n572_), .B2(new_n569_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n253_), .A2(KEYINPUT70), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n566_), .A2(new_n575_), .A3(KEYINPUT12), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT12), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n253_), .B(new_n565_), .C1(KEYINPUT70), .C2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n561_), .A2(new_n569_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT71), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT71), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n561_), .A2(new_n582_), .A3(new_n569_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n579_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n574_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G120gat), .B(G148gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT5), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(G176gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(new_n381_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n586_), .A2(new_n590_), .ZN(new_n591_));
  AOI22_X1  g390(.A1(new_n571_), .A2(new_n573_), .B1(new_n579_), .B2(new_n584_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n590_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n560_), .B1(new_n591_), .B2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n586_), .A2(new_n590_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n592_), .A2(new_n593_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(new_n597_), .A3(KEYINPUT13), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n595_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT72), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n543_), .A2(new_n559_), .A3(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n516_), .B(KEYINPUT107), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n602_), .A2(new_n317_), .A3(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT38), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n599_), .A2(new_n558_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n542_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n282_), .A2(new_n289_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n328_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n608_), .A2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G1gat), .B1(new_n613_), .B2(new_n517_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n606_), .A2(new_n614_), .ZN(G1324gat));
  NAND3_X1  g414(.A1(new_n602_), .A2(new_n318_), .A3(new_n480_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n480_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G8gat), .B1(new_n613_), .B2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT39), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n616_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT40), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(G1325gat));
  OAI21_X1  g421(.A(G15gat), .B1(new_n613_), .B2(new_n494_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT41), .Z(new_n624_));
  INV_X1    g423(.A(G15gat), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n602_), .A2(new_n625_), .A3(new_n493_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(G1326gat));
  OAI21_X1  g426(.A(G22gat), .B1(new_n613_), .B2(new_n519_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT108), .Z(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT42), .ZN(new_n630_));
  INV_X1    g429(.A(G22gat), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n602_), .A2(new_n631_), .A3(new_n408_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(G1327gat));
  INV_X1    g432(.A(KEYINPUT43), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n291_), .A2(new_n293_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n634_), .B1(new_n542_), .B2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n540_), .A2(new_n519_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n617_), .A2(new_n517_), .A3(new_n408_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n493_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n495_), .A2(new_n517_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n634_), .B(new_n635_), .C1(new_n639_), .C2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n611_), .B(new_n607_), .C1(new_n636_), .C2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT44), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n639_), .A2(new_n640_), .ZN(new_n646_));
  OAI21_X1  g445(.A(KEYINPUT43), .B1(new_n646_), .B2(new_n294_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(new_n641_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n648_), .A2(KEYINPUT44), .A3(new_n611_), .A4(new_n607_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n645_), .A2(new_n604_), .A3(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(G29gat), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n609_), .A2(new_n328_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT109), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n608_), .A2(new_n653_), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n517_), .A2(G29gat), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n651_), .B1(new_n654_), .B2(new_n655_), .ZN(G1328gat));
  INV_X1    g455(.A(KEYINPUT46), .ZN(new_n657_));
  INV_X1    g456(.A(G36gat), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(KEYINPUT45), .ZN(new_n659_));
  INV_X1    g458(.A(new_n654_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n660_), .B2(new_n480_), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n661_), .A2(KEYINPUT110), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n645_), .A2(KEYINPUT45), .A3(new_n649_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n660_), .A2(new_n658_), .ZN(new_n664_));
  AOI22_X1  g463(.A1(new_n663_), .A2(new_n664_), .B1(KEYINPUT45), .B2(new_n658_), .ZN(new_n665_));
  AOI211_X1 g464(.A(new_n657_), .B(new_n662_), .C1(new_n665_), .C2(new_n480_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n663_), .A2(new_n664_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n667_), .A2(new_n480_), .A3(new_n659_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n662_), .ZN(new_n669_));
  AOI21_X1  g468(.A(KEYINPUT46), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n666_), .A2(new_n670_), .ZN(G1329gat));
  NAND3_X1  g470(.A1(new_n660_), .A2(new_n203_), .A3(new_n493_), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n645_), .A2(new_n493_), .A3(new_n649_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n672_), .B1(new_n673_), .B2(new_n203_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT47), .Z(G1330gat));
  NAND3_X1  g474(.A1(new_n645_), .A2(new_n408_), .A3(new_n649_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT111), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n677_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n678_), .A2(G50gat), .A3(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n660_), .A2(new_n207_), .A3(new_n408_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1331gat));
  NAND3_X1  g481(.A1(new_n542_), .A2(new_n558_), .A3(new_n600_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(new_n612_), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n685_), .A2(new_n508_), .A3(new_n517_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n559_), .B1(new_n595_), .B2(new_n598_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n543_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n604_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n686_), .B1(new_n690_), .B2(new_n508_), .ZN(G1332gat));
  OR3_X1    g490(.A1(new_n688_), .A2(G64gat), .A3(new_n617_), .ZN(new_n692_));
  OAI21_X1  g491(.A(G64gat), .B1(new_n685_), .B2(new_n617_), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n693_), .A2(KEYINPUT112), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(KEYINPUT112), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n694_), .A2(KEYINPUT48), .A3(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(KEYINPUT48), .B1(new_n694_), .B2(new_n695_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n692_), .B1(new_n696_), .B2(new_n697_), .ZN(G1333gat));
  OR3_X1    g497(.A1(new_n688_), .A2(G71gat), .A3(new_n494_), .ZN(new_n699_));
  OAI21_X1  g498(.A(G71gat), .B1(new_n685_), .B2(new_n494_), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n700_), .A2(KEYINPUT113), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(KEYINPUT113), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n701_), .A2(KEYINPUT49), .A3(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT49), .B1(new_n701_), .B2(new_n702_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n699_), .B1(new_n703_), .B2(new_n704_), .ZN(G1334gat));
  OAI21_X1  g504(.A(G78gat), .B1(new_n685_), .B2(new_n519_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT50), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n519_), .A2(G78gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n707_), .B1(new_n688_), .B2(new_n708_), .ZN(G1335gat));
  NAND2_X1  g508(.A1(new_n684_), .A2(new_n653_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(G85gat), .B1(new_n711_), .B2(new_n604_), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n648_), .A2(new_n611_), .A3(new_n687_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n517_), .A2(new_n218_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n712_), .B1(new_n713_), .B2(new_n714_), .ZN(G1336gat));
  AOI21_X1  g514(.A(G92gat), .B1(new_n711_), .B2(new_n480_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n617_), .A2(new_n219_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n713_), .B2(new_n717_), .ZN(G1337gat));
  NOR3_X1   g517(.A1(new_n710_), .A2(new_n229_), .A3(new_n494_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n713_), .A2(new_n493_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n720_), .B2(G99gat), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT51), .Z(G1338gat));
  NAND4_X1  g521(.A1(new_n648_), .A2(new_n611_), .A3(new_n408_), .A4(new_n687_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G106gat), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT114), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT52), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n724_), .A2(new_n725_), .A3(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n711_), .A2(new_n238_), .A3(new_n408_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(KEYINPUT114), .A2(KEYINPUT52), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n725_), .A2(new_n726_), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n723_), .A2(G106gat), .A3(new_n729_), .A4(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n727_), .A2(new_n728_), .A3(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g532(.A(KEYINPUT119), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT57), .ZN(new_n735_));
  NOR2_X1   g534(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n579_), .A2(new_n584_), .A3(KEYINPUT55), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n569_), .B1(new_n579_), .B2(new_n564_), .ZN(new_n739_));
  AOI21_X1  g538(.A(KEYINPUT55), .B1(new_n579_), .B2(new_n584_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n738_), .A2(new_n739_), .A3(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n741_), .B2(new_n593_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n558_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT55), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n585_), .A2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n579_), .A2(new_n584_), .A3(KEYINPUT55), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n590_), .B(new_n736_), .C1(new_n747_), .C2(new_n739_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n742_), .A2(new_n743_), .A3(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT117), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n548_), .A2(new_n546_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n545_), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n751_), .B(new_n553_), .C1(new_n752_), .C2(new_n546_), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n555_), .B(new_n753_), .C1(new_n591_), .C2(new_n594_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT117), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n742_), .A2(new_n743_), .A3(new_n755_), .A4(new_n748_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n750_), .A2(new_n754_), .A3(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n609_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT118), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n735_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  AOI211_X1 g559(.A(KEYINPUT118), .B(KEYINPUT57), .C1(new_n757_), .C2(new_n609_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(KEYINPUT56), .B1(new_n741_), .B2(new_n593_), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n763_), .A2(new_n555_), .A3(new_n753_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT56), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n765_), .B(new_n590_), .C1(new_n747_), .C2(new_n739_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n764_), .A2(new_n597_), .A3(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT58), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n768_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n635_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n328_), .B1(new_n762_), .B2(new_n771_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n595_), .A2(new_n598_), .A3(new_n328_), .A4(new_n558_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT115), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n773_), .B(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT54), .B1(new_n775_), .B2(new_n635_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n773_), .B(KEYINPUT115), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT54), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n294_), .A2(new_n777_), .A3(new_n778_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n776_), .A2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n734_), .B1(new_n772_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n758_), .A2(new_n759_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT57), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n758_), .A2(new_n759_), .A3(new_n735_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n783_), .A2(new_n771_), .A3(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n611_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n776_), .A2(new_n779_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(KEYINPUT119), .A3(new_n787_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n495_), .A2(new_n604_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n781_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(G113gat), .B1(new_n791_), .B2(new_n559_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(KEYINPUT59), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT120), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n786_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n785_), .A2(KEYINPUT120), .A3(new_n611_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n787_), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT59), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(new_n798_), .A3(new_n789_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n793_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT121), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT121), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n793_), .A2(new_n802_), .A3(new_n799_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n558_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n792_), .B1(new_n804_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g604(.A(G120gat), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT60), .B1(new_n599_), .B2(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n790_), .A2(new_n807_), .ZN(new_n808_));
  NOR3_X1   g607(.A1(new_n800_), .A2(new_n601_), .A3(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n808_), .ZN(new_n810_));
  OAI22_X1  g609(.A1(new_n809_), .A2(new_n806_), .B1(KEYINPUT60), .B2(new_n810_), .ZN(G1341gat));
  AOI21_X1  g610(.A(G127gat), .B1(new_n791_), .B2(new_n328_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n611_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n813_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g613(.A(G134gat), .B1(new_n791_), .B2(new_n610_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n294_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n815_), .B1(new_n816_), .B2(G134gat), .ZN(G1343gat));
  NAND4_X1  g616(.A1(new_n781_), .A2(new_n788_), .A3(new_n520_), .A4(new_n494_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n818_), .A2(new_n603_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n559_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n600_), .ZN(new_n822_));
  XOR2_X1   g621(.A(KEYINPUT122), .B(G148gat), .Z(new_n823_));
  XNOR2_X1  g622(.A(new_n822_), .B(new_n823_), .ZN(G1345gat));
  INV_X1    g623(.A(KEYINPUT123), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n825_), .B1(new_n819_), .B2(new_n328_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(KEYINPUT61), .B(G155gat), .ZN(new_n828_));
  NOR4_X1   g627(.A1(new_n818_), .A2(KEYINPUT123), .A3(new_n611_), .A4(new_n603_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n827_), .A2(new_n828_), .A3(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n828_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n832_), .B1(new_n826_), .B2(new_n829_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(G1346gat));
  AOI21_X1  g633(.A(G162gat), .B1(new_n819_), .B2(new_n610_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n294_), .A2(new_n279_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n819_), .B2(new_n836_), .ZN(G1347gat));
  NOR4_X1   g636(.A1(new_n604_), .A2(new_n617_), .A3(new_n408_), .A4(new_n494_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n797_), .A2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT124), .B1(new_n839_), .B2(new_n558_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT124), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n797_), .A2(new_n841_), .A3(new_n559_), .A4(new_n838_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n840_), .A2(G169gat), .A3(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT62), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n839_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n846_), .A2(new_n559_), .A3(new_n423_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n840_), .A2(KEYINPUT62), .A3(G169gat), .A4(new_n842_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n845_), .A2(new_n847_), .A3(new_n848_), .ZN(G1348gat));
  AOI21_X1  g648(.A(G176gat), .B1(new_n846_), .B2(new_n599_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n781_), .A2(new_n788_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n851_), .A2(new_n838_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n601_), .A2(new_n420_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n850_), .B1(new_n852_), .B2(new_n853_), .ZN(G1349gat));
  OR3_X1    g653(.A1(new_n839_), .A2(new_n611_), .A3(new_n446_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n855_), .A2(KEYINPUT125), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n855_), .A2(KEYINPUT125), .ZN(new_n857_));
  AOI21_X1  g656(.A(G183gat), .B1(new_n852_), .B2(new_n328_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n856_), .A2(new_n857_), .A3(new_n858_), .ZN(G1350gat));
  NAND3_X1  g658(.A1(new_n846_), .A2(new_n610_), .A3(new_n436_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n846_), .A2(new_n635_), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n861_), .A2(KEYINPUT126), .A3(G190gat), .ZN(new_n862_));
  AOI21_X1  g661(.A(KEYINPUT126), .B1(new_n861_), .B2(G190gat), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n860_), .B1(new_n862_), .B2(new_n863_), .ZN(G1351gat));
  NAND3_X1  g663(.A1(new_n851_), .A2(new_n480_), .A3(new_n494_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n408_), .A2(new_n517_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n865_), .A2(new_n558_), .A3(new_n866_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(new_n552_), .ZN(G1352gat));
  NOR3_X1   g667(.A1(new_n865_), .A2(new_n601_), .A3(new_n866_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(new_n381_), .ZN(G1353gat));
  XNOR2_X1  g669(.A(KEYINPUT63), .B(G211gat), .ZN(new_n871_));
  NOR4_X1   g670(.A1(new_n865_), .A2(new_n611_), .A3(new_n866_), .A4(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n865_), .A2(new_n866_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n328_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n872_), .B1(new_n874_), .B2(new_n875_), .ZN(G1354gat));
  NAND2_X1  g675(.A1(new_n873_), .A2(new_n610_), .ZN(new_n877_));
  INV_X1    g676(.A(G218gat), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n294_), .A2(new_n878_), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n877_), .A2(new_n878_), .B1(new_n873_), .B2(new_n879_), .ZN(G1355gat));
endmodule


