//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 1 1 1 0 1 1 0 1 0 1 0 1 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n615_, new_n616_, new_n617_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n885_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT18), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G64gat), .B(G92gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G226gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT21), .ZN(new_n210_));
  AND2_X1   g009(.A1(G197gat), .A2(G204gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G197gat), .A2(G204gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n210_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT90), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  OAI211_X1 g014(.A(KEYINPUT90), .B(new_n210_), .C1(new_n211_), .C2(new_n212_), .ZN(new_n216_));
  INV_X1    g015(.A(G197gat), .ZN(new_n217_));
  INV_X1    g016(.A(G204gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT89), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G197gat), .A2(G204gat), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n219_), .A2(new_n220_), .A3(KEYINPUT21), .A4(new_n221_), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n215_), .A2(new_n216_), .A3(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G211gat), .B(G218gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n219_), .A2(KEYINPUT21), .A3(new_n221_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n225_), .B1(KEYINPUT89), .B2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT91), .B1(new_n226_), .B2(new_n224_), .ZN(new_n228_));
  OR3_X1    g027(.A1(new_n226_), .A2(new_n224_), .A3(KEYINPUT91), .ZN(new_n229_));
  AOI22_X1  g028(.A1(new_n223_), .A2(new_n227_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G183gat), .A2(G190gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT81), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT81), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n234_), .A2(G183gat), .A3(G190gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n231_), .B1(new_n236_), .B2(KEYINPUT23), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n237_), .B1(G183gat), .B2(G190gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT83), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT22), .ZN(new_n240_));
  INV_X1    g039(.A(G176gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT83), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(G169gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n238_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT23), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n247_), .B1(G183gat), .B2(G190gat), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n248_), .B1(new_n236_), .B2(new_n247_), .ZN(new_n249_));
  NOR3_X1   g048(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT82), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT82), .ZN(new_n252_));
  INV_X1    g051(.A(new_n250_), .ZN(new_n253_));
  AOI21_X1  g052(.A(KEYINPUT23), .B1(new_n233_), .B2(new_n235_), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n252_), .B(new_n253_), .C1(new_n254_), .C2(new_n248_), .ZN(new_n255_));
  OAI21_X1  g054(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n256_));
  AND2_X1   g055(.A1(G169gat), .A2(G176gat), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT25), .ZN(new_n259_));
  AOI21_X1  g058(.A(KEYINPUT79), .B1(new_n259_), .B2(G183gat), .ZN(new_n260_));
  INV_X1    g059(.A(G183gat), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n260_), .B1(KEYINPUT25), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(KEYINPUT80), .A2(G190gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT26), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT26), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(KEYINPUT80), .A3(G190gat), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n259_), .A2(KEYINPUT79), .A3(G183gat), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n264_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n258_), .B1(new_n262_), .B2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n251_), .A2(new_n255_), .A3(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n230_), .A2(new_n246_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT95), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(new_n272_), .A3(KEYINPUT20), .ZN(new_n273_));
  INV_X1    g072(.A(new_n230_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT22), .B(G169gat), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n257_), .B1(new_n275_), .B2(new_n241_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(G183gat), .A2(G190gat), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n276_), .B1(new_n249_), .B2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT26), .B(G190gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n261_), .A2(KEYINPUT25), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n259_), .A2(G183gat), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n258_), .A2(new_n250_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n237_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n278_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n274_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n273_), .A2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n272_), .B1(new_n271_), .B2(KEYINPUT20), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n209_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT96), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT96), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n291_), .B(new_n209_), .C1(new_n287_), .C2(new_n288_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n270_), .A2(new_n246_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(new_n274_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT20), .ZN(new_n296_));
  INV_X1    g095(.A(new_n209_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n297_), .B1(new_n274_), .B2(new_n285_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n206_), .B1(new_n293_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n206_), .ZN(new_n302_));
  AOI211_X1 g101(.A(new_n302_), .B(new_n299_), .C1(new_n290_), .C2(new_n292_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n202_), .B1(new_n301_), .B2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n293_), .A2(new_n206_), .A3(new_n300_), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n278_), .A2(KEYINPUT97), .A3(new_n284_), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT97), .B1(new_n278_), .B2(new_n284_), .ZN(new_n307_));
  NOR3_X1   g106(.A1(new_n274_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n209_), .B1(new_n296_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n271_), .A2(KEYINPUT20), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT95), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n311_), .A2(new_n286_), .A3(new_n273_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n309_), .B1(new_n312_), .B2(new_n209_), .ZN(new_n313_));
  AOI21_X1  g112(.A(KEYINPUT99), .B1(new_n313_), .B2(new_n302_), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n313_), .A2(KEYINPUT99), .A3(new_n302_), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n305_), .B(KEYINPUT27), .C1(new_n314_), .C2(new_n315_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n304_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n294_), .B(KEYINPUT30), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n318_), .A2(KEYINPUT85), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n318_), .A2(KEYINPUT85), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G227gat), .A2(G233gat), .ZN(new_n322_));
  INV_X1    g121(.A(G71gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(G99gat), .ZN(new_n325_));
  XOR2_X1   g124(.A(G15gat), .B(G43gat), .Z(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT84), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n325_), .B(new_n327_), .Z(new_n328_));
  NOR2_X1   g127(.A1(new_n321_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n328_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n319_), .A2(new_n330_), .ZN(new_n331_));
  XOR2_X1   g130(.A(G127gat), .B(G134gat), .Z(new_n332_));
  XOR2_X1   g131(.A(G113gat), .B(G120gat), .Z(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT86), .B(KEYINPUT31), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  OR3_X1    g136(.A1(new_n329_), .A2(new_n331_), .A3(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n337_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n332_), .B(new_n333_), .Z(new_n340_));
  OR2_X1    g139(.A1(G155gat), .A2(G162gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G155gat), .A2(G162gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT87), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT3), .ZN(new_n346_));
  INV_X1    g145(.A(G141gat), .ZN(new_n347_));
  INV_X1    g146(.A(G148gat), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G141gat), .A2(G148gat), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT2), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n349_), .A2(new_n352_), .A3(new_n353_), .A4(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n341_), .A2(KEYINPUT87), .A3(new_n342_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n345_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n347_), .A2(new_n348_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n342_), .A2(KEYINPUT1), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n341_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n342_), .A2(KEYINPUT1), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n350_), .B(new_n358_), .C1(new_n360_), .C2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n357_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n340_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n334_), .A2(new_n362_), .A3(new_n357_), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n364_), .A2(KEYINPUT4), .A3(new_n365_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT4), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n340_), .A2(new_n363_), .A3(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n367_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G1gat), .B(G29gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(G85gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT0), .B(G57gat), .ZN(new_n376_));
  XOR2_X1   g175(.A(new_n375_), .B(new_n376_), .Z(new_n377_));
  OR3_X1    g176(.A1(new_n369_), .A2(new_n373_), .A3(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n377_), .B1(new_n369_), .B2(new_n373_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n378_), .A2(new_n379_), .A3(KEYINPUT98), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT98), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n381_), .B(new_n377_), .C1(new_n369_), .C2(new_n373_), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n363_), .A2(KEYINPUT29), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G228gat), .A2(G233gat), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n274_), .B(new_n385_), .C1(KEYINPUT92), .C2(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n230_), .B1(KEYINPUT29), .B2(new_n363_), .ZN(new_n388_));
  XOR2_X1   g187(.A(new_n386_), .B(KEYINPUT92), .Z(new_n389_));
  OAI21_X1  g188(.A(new_n387_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G78gat), .B(G106gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n391_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n387_), .B(new_n393_), .C1(new_n388_), .C2(new_n389_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  OR2_X1    g194(.A1(new_n363_), .A2(KEYINPUT29), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XOR2_X1   g197(.A(G22gat), .B(G50gat), .Z(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n398_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT93), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n402_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n395_), .B1(new_n401_), .B2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n398_), .B(new_n399_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n405_), .A2(new_n402_), .A3(new_n392_), .A4(new_n394_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  AND4_X1   g206(.A1(new_n338_), .A2(new_n339_), .A3(new_n384_), .A4(new_n407_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n317_), .A2(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n383_), .A2(new_n407_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n304_), .A2(new_n316_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT100), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT100), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n304_), .A2(new_n316_), .A3(new_n413_), .A4(new_n410_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n292_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n291_), .B1(new_n312_), .B2(new_n209_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n300_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n302_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n377_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n370_), .A2(new_n367_), .A3(new_n372_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT33), .ZN(new_n422_));
  MUX2_X1   g221(.A(KEYINPUT33), .B(new_n422_), .S(new_n379_), .Z(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n418_), .A2(new_n305_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n206_), .A2(KEYINPUT32), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n313_), .A2(new_n427_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n383_), .B(new_n428_), .C1(new_n417_), .C2(new_n427_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n425_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n407_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n412_), .A2(new_n414_), .A3(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n338_), .A2(new_n339_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n409_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G29gat), .B(G36gat), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(G43gat), .B(G50gat), .Z(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT15), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G15gat), .B(G22gat), .ZN(new_n440_));
  INV_X1    g239(.A(G1gat), .ZN(new_n441_));
  INV_X1    g240(.A(G8gat), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT14), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n440_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G1gat), .B(G8gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n439_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n438_), .ZN(new_n448_));
  OR2_X1    g247(.A1(new_n448_), .A2(new_n446_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G229gat), .A2(G233gat), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n447_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n448_), .B(new_n446_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n450_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n451_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G113gat), .B(G141gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G169gat), .B(G197gat), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n456_), .B(new_n457_), .Z(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n455_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n451_), .A2(new_n454_), .A3(new_n458_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n434_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G99gat), .A2(G106gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT6), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT6), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n467_), .A2(G99gat), .A3(G106gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G85gat), .A2(G92gat), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n469_), .B1(KEYINPUT9), .B2(new_n470_), .ZN(new_n471_));
  OR2_X1    g270(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n472_));
  INV_X1    g271(.A(G106gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(G85gat), .ZN(new_n476_));
  INV_X1    g275(.A(G92gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(KEYINPUT9), .A3(new_n470_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n475_), .A2(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT65), .B1(new_n471_), .B2(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n470_), .A2(KEYINPUT9), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n482_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT65), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n483_), .A2(new_n484_), .A3(new_n475_), .A4(new_n479_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n481_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT66), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n469_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT67), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NOR3_X1   g290(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n489_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n466_), .A2(new_n468_), .A3(KEYINPUT66), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT7), .ZN(new_n495_));
  INV_X1    g294(.A(G99gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(new_n496_), .A3(new_n473_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n497_), .A2(KEYINPUT67), .A3(new_n490_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n488_), .A2(new_n493_), .A3(new_n494_), .A4(new_n498_), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n478_), .A2(new_n470_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n500_), .A2(KEYINPUT8), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT70), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n469_), .A2(new_n497_), .A3(new_n490_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n500_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT8), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n502_), .A2(new_n503_), .A3(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n503_), .B1(new_n502_), .B2(new_n507_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n486_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(new_n439_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT72), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n510_), .A2(KEYINPUT72), .A3(new_n439_), .ZN(new_n514_));
  AOI21_X1  g313(.A(KEYINPUT73), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G232gat), .A2(G233gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT34), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT35), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n515_), .A2(new_n518_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n502_), .A2(new_n507_), .A3(new_n485_), .A4(new_n481_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT68), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n486_), .A2(KEYINPUT68), .A3(new_n507_), .A4(new_n502_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n513_), .A2(new_n514_), .B1(new_n438_), .B2(new_n524_), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n517_), .A2(KEYINPUT35), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n519_), .A2(new_n527_), .ZN(new_n528_));
  NOR3_X1   g327(.A1(new_n525_), .A2(new_n515_), .A3(new_n518_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT36), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G134gat), .B(G162gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT76), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G190gat), .B(G218gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n528_), .A2(new_n530_), .A3(new_n531_), .A4(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n531_), .ZN(new_n539_));
  OR2_X1    g338(.A1(new_n537_), .A2(new_n531_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n519_), .A2(new_n527_), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n539_), .B(new_n540_), .C1(new_n541_), .C2(new_n529_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n538_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT37), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G57gat), .B(G64gat), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n545_), .A2(KEYINPUT11), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G71gat), .B(G78gat), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT69), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n547_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT69), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n549_), .B(new_n550_), .C1(KEYINPUT11), .C2(new_n545_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n548_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n545_), .A2(KEYINPUT11), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n548_), .A2(KEYINPUT11), .A3(new_n551_), .A4(new_n545_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n524_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n522_), .A2(new_n523_), .A3(new_n556_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G230gat), .A2(G233gat), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n561_), .B(KEYINPUT64), .Z(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n560_), .A2(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n563_), .B1(new_n524_), .B2(new_n557_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT12), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n559_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n510_), .A2(KEYINPUT12), .A3(new_n556_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n565_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n564_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G120gat), .B(G148gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT5), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G176gat), .B(G204gat), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n572_), .B(new_n573_), .Z(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n575_), .A2(KEYINPUT71), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n570_), .B(new_n576_), .Z(new_n577_));
  OR2_X1    g376(.A1(new_n577_), .A2(KEYINPUT13), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(KEYINPUT13), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n446_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(new_n556_), .ZN(new_n583_));
  XOR2_X1   g382(.A(G127gat), .B(G155gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(G183gat), .B(G211gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(KEYINPUT17), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n583_), .A2(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n588_), .B(KEYINPUT17), .Z(new_n591_));
  OAI21_X1  g390(.A(new_n590_), .B1(new_n591_), .B2(new_n583_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n592_), .A2(KEYINPUT78), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(KEYINPUT78), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n544_), .A2(new_n580_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n464_), .A2(new_n598_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n599_), .A2(G1gat), .A3(new_n384_), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n600_), .A2(KEYINPUT38), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(KEYINPUT38), .ZN(new_n602_));
  INV_X1    g401(.A(new_n543_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n434_), .A2(new_n603_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n604_), .A2(new_n462_), .A3(new_n580_), .A4(new_n596_), .ZN(new_n605_));
  OAI21_X1  g404(.A(G1gat), .B1(new_n605_), .B2(new_n384_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n601_), .A2(new_n602_), .A3(new_n606_), .ZN(G1324gat));
  OAI21_X1  g406(.A(G8gat), .B1(new_n605_), .B2(new_n317_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT39), .ZN(new_n609_));
  INV_X1    g408(.A(new_n317_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(new_n442_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n609_), .B1(new_n599_), .B2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(G1325gat));
  OAI21_X1  g413(.A(G15gat), .B1(new_n605_), .B2(new_n433_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT41), .ZN(new_n616_));
  NOR3_X1   g415(.A1(new_n599_), .A2(G15gat), .A3(new_n433_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1326gat));
  OAI21_X1  g417(.A(G22gat), .B1(new_n605_), .B2(new_n407_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT42), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n407_), .A2(G22gat), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n621_), .B(KEYINPUT102), .Z(new_n622_));
  OAI21_X1  g421(.A(new_n620_), .B1(new_n599_), .B2(new_n622_), .ZN(G1327gat));
  INV_X1    g422(.A(new_n580_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n603_), .A2(new_n595_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n464_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  OR3_X1    g427(.A1(new_n628_), .A2(G29gat), .A3(new_n384_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n624_), .A2(new_n463_), .A3(new_n596_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT103), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n631_), .B(KEYINPUT43), .C1(new_n434_), .C2(new_n544_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT37), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n543_), .B(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n433_), .ZN(new_n636_));
  AOI22_X1  g435(.A1(new_n411_), .A2(KEYINPUT100), .B1(new_n430_), .B2(new_n407_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n636_), .B1(new_n637_), .B2(new_n414_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n635_), .B1(new_n638_), .B2(new_n409_), .ZN(new_n639_));
  AOI21_X1  g438(.A(KEYINPUT43), .B1(new_n639_), .B2(new_n631_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n630_), .B1(new_n633_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT44), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n641_), .A2(new_n642_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(new_n383_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n646_), .A2(KEYINPUT104), .ZN(new_n647_));
  OAI21_X1  g446(.A(G29gat), .B1(new_n646_), .B2(KEYINPUT104), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n629_), .B1(new_n647_), .B2(new_n648_), .ZN(G1328gat));
  INV_X1    g448(.A(G36gat), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n627_), .A2(new_n650_), .A3(new_n610_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n651_), .B(new_n652_), .Z(new_n653_));
  NOR3_X1   g452(.A1(new_n643_), .A2(new_n644_), .A3(new_n317_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n653_), .B1(new_n654_), .B2(new_n650_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(KEYINPUT106), .B(KEYINPUT46), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n653_), .B(new_n656_), .C1(new_n654_), .C2(new_n650_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1329gat));
  NAND3_X1  g459(.A1(new_n645_), .A2(G43gat), .A3(new_n636_), .ZN(new_n661_));
  INV_X1    g460(.A(G43gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n662_), .B1(new_n628_), .B2(new_n433_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n661_), .A2(KEYINPUT47), .A3(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT47), .B1(new_n661_), .B2(new_n663_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1330gat));
  INV_X1    g465(.A(new_n407_), .ZN(new_n667_));
  AOI21_X1  g466(.A(G50gat), .B1(new_n627_), .B2(new_n667_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n667_), .A2(G50gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n645_), .B2(new_n669_), .ZN(G1331gat));
  NOR2_X1   g469(.A1(new_n434_), .A2(new_n462_), .ZN(new_n671_));
  AND4_X1   g470(.A1(new_n624_), .A2(new_n671_), .A3(new_n596_), .A4(new_n544_), .ZN(new_n672_));
  INV_X1    g471(.A(G57gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n672_), .A2(new_n673_), .A3(new_n383_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n604_), .A2(new_n463_), .A3(new_n624_), .A4(new_n596_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT107), .Z(new_n676_));
  AND2_X1   g475(.A1(new_n676_), .A2(new_n383_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n674_), .B1(new_n677_), .B2(new_n673_), .ZN(G1332gat));
  NOR2_X1   g477(.A1(new_n317_), .A2(G64gat), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT109), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n672_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n676_), .A2(new_n610_), .ZN(new_n682_));
  XOR2_X1   g481(.A(KEYINPUT108), .B(KEYINPUT48), .Z(new_n683_));
  AND3_X1   g482(.A1(new_n682_), .A2(G64gat), .A3(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n682_), .B2(G64gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n681_), .B1(new_n684_), .B2(new_n685_), .ZN(G1333gat));
  NAND3_X1  g485(.A1(new_n672_), .A2(new_n323_), .A3(new_n636_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT49), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n676_), .A2(new_n636_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(G71gat), .ZN(new_n690_));
  AOI211_X1 g489(.A(KEYINPUT49), .B(new_n323_), .C1(new_n676_), .C2(new_n636_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n687_), .B1(new_n690_), .B2(new_n691_), .ZN(G1334gat));
  INV_X1    g491(.A(G78gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n672_), .A2(new_n693_), .A3(new_n667_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT50), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n676_), .A2(new_n667_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n696_), .B2(G78gat), .ZN(new_n697_));
  AOI211_X1 g496(.A(KEYINPUT50), .B(new_n693_), .C1(new_n676_), .C2(new_n667_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n694_), .B1(new_n697_), .B2(new_n698_), .ZN(G1335gat));
  NOR2_X1   g498(.A1(new_n625_), .A2(new_n580_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n671_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n702_), .A2(new_n476_), .A3(new_n383_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n624_), .A2(new_n463_), .A3(new_n595_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n631_), .B1(new_n434_), .B2(new_n544_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n704_), .B1(new_n707_), .B2(new_n632_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n708_), .A2(KEYINPUT110), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n708_), .A2(KEYINPUT110), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n709_), .A2(new_n710_), .A3(new_n384_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n703_), .B1(new_n711_), .B2(new_n476_), .ZN(G1336gat));
  NAND3_X1  g511(.A1(new_n702_), .A2(new_n477_), .A3(new_n610_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n709_), .A2(new_n710_), .A3(new_n317_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n713_), .B1(new_n714_), .B2(new_n477_), .ZN(G1337gat));
  AND2_X1   g514(.A1(new_n708_), .A2(new_n636_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n472_), .A2(new_n474_), .ZN(new_n717_));
  OR2_X1    g516(.A1(new_n433_), .A2(new_n717_), .ZN(new_n718_));
  OAI22_X1  g517(.A1(new_n716_), .A2(new_n496_), .B1(new_n701_), .B2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g519(.A1(new_n702_), .A2(new_n473_), .A3(new_n667_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT52), .ZN(new_n722_));
  AOI211_X1 g521(.A(new_n407_), .B(new_n704_), .C1(new_n707_), .C2(new_n632_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n473_), .B1(new_n723_), .B2(KEYINPUT111), .ZN(new_n724_));
  INV_X1    g523(.A(new_n704_), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n667_), .B(new_n725_), .C1(new_n633_), .C2(new_n640_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT111), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n722_), .B1(new_n724_), .B2(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G106gat), .B1(new_n726_), .B2(new_n727_), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT111), .B1(new_n708_), .B2(new_n667_), .ZN(new_n731_));
  NOR3_X1   g530(.A1(new_n730_), .A2(new_n731_), .A3(KEYINPUT52), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n721_), .B1(new_n729_), .B2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT53), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT53), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n735_), .B(new_n721_), .C1(new_n729_), .C2(new_n732_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(G1339gat));
  NOR3_X1   g536(.A1(new_n610_), .A2(new_n433_), .A3(new_n384_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT117), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT114), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT55), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n567_), .A2(new_n558_), .A3(new_n568_), .ZN(new_n742_));
  AOI22_X1  g541(.A1(new_n741_), .A2(new_n569_), .B1(new_n742_), .B2(new_n563_), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n565_), .A2(new_n567_), .A3(KEYINPUT55), .A4(new_n568_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n575_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n740_), .B1(new_n745_), .B2(KEYINPUT56), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n569_), .A2(new_n741_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n742_), .A2(new_n563_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n747_), .A2(new_n748_), .A3(new_n744_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n749_), .A2(KEYINPUT56), .A3(new_n574_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT113), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n574_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT56), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(KEYINPUT114), .A3(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT113), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n749_), .A2(new_n755_), .A3(KEYINPUT56), .A4(new_n574_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n746_), .A2(new_n751_), .A3(new_n754_), .A4(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT115), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n447_), .A2(new_n449_), .A3(new_n453_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n452_), .A2(new_n450_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n759_), .A2(new_n459_), .A3(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n762_), .A2(KEYINPUT112), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(KEYINPUT112), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n763_), .A2(new_n461_), .A3(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n564_), .A2(new_n569_), .A3(new_n575_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n765_), .A2(new_n767_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n757_), .A2(new_n758_), .A3(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n758_), .B1(new_n757_), .B2(new_n768_), .ZN(new_n770_));
  XOR2_X1   g569(.A(KEYINPUT116), .B(KEYINPUT58), .Z(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n769_), .A2(new_n770_), .A3(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n739_), .B1(new_n773_), .B2(new_n544_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n757_), .A2(new_n768_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT58), .ZN(new_n777_));
  INV_X1    g576(.A(new_n770_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n757_), .A2(new_n758_), .A3(new_n768_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(new_n779_), .A3(new_n771_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n780_), .A2(KEYINPUT117), .A3(new_n635_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n774_), .A2(new_n777_), .A3(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n752_), .A2(new_n753_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n750_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n784_), .A2(new_n462_), .A3(new_n766_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(new_n577_), .B2(new_n765_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT118), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT57), .ZN(new_n788_));
  AOI22_X1  g587(.A1(new_n538_), .A2(new_n542_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n786_), .A2(new_n789_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n787_), .A2(new_n788_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n790_), .B(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n596_), .B1(new_n782_), .B2(new_n794_), .ZN(new_n795_));
  OR3_X1    g594(.A1(new_n597_), .A2(KEYINPUT54), .A3(new_n462_), .ZN(new_n796_));
  OAI21_X1  g595(.A(KEYINPUT54), .B1(new_n597_), .B2(new_n462_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n407_), .B(new_n738_), .C1(new_n795_), .C2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT59), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n796_), .A2(new_n797_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n770_), .A2(new_n772_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n544_), .B1(new_n803_), .B2(new_n779_), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n804_), .A2(KEYINPUT117), .B1(KEYINPUT58), .B2(new_n776_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n793_), .B1(new_n805_), .B2(new_n774_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n802_), .B1(new_n806_), .B2(new_n596_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n807_), .A2(KEYINPUT59), .A3(new_n407_), .A4(new_n738_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n801_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n462_), .A2(G113gat), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(KEYINPUT119), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT120), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n807_), .A2(new_n407_), .A3(new_n462_), .A4(new_n738_), .ZN(new_n814_));
  INV_X1    g613(.A(G113gat), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n812_), .A2(new_n813_), .A3(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n811_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n818_), .B1(new_n801_), .B2(new_n808_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n799_), .ZN(new_n820_));
  AOI21_X1  g619(.A(G113gat), .B1(new_n820_), .B2(new_n462_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT120), .B1(new_n819_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n817_), .A2(new_n822_), .ZN(G1340gat));
  AOI21_X1  g622(.A(new_n580_), .B1(new_n801_), .B2(new_n808_), .ZN(new_n824_));
  INV_X1    g623(.A(G120gat), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n825_), .B1(new_n580_), .B2(KEYINPUT60), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(KEYINPUT60), .B2(new_n825_), .ZN(new_n827_));
  OAI22_X1  g626(.A1(new_n824_), .A2(new_n825_), .B1(new_n799_), .B2(new_n827_), .ZN(G1341gat));
  INV_X1    g627(.A(G127gat), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n820_), .A2(new_n829_), .A3(new_n596_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n595_), .B1(new_n801_), .B2(new_n808_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n831_), .B2(new_n829_), .ZN(G1342gat));
  INV_X1    g631(.A(G134gat), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n820_), .A2(new_n833_), .A3(new_n603_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n544_), .B1(new_n801_), .B2(new_n808_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(new_n833_), .ZN(G1343gat));
  NOR2_X1   g635(.A1(new_n636_), .A2(new_n407_), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n837_), .A2(new_n317_), .A3(new_n383_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n807_), .A2(new_n838_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(new_n463_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(new_n347_), .ZN(G1344gat));
  AND2_X1   g640(.A1(new_n807_), .A2(new_n838_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT122), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n843_), .A3(new_n624_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT122), .B1(new_n839_), .B2(new_n580_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(KEYINPUT121), .B(G148gat), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n844_), .A2(new_n845_), .A3(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1345gat));
  NAND3_X1  g648(.A1(new_n842_), .A2(KEYINPUT123), .A3(new_n596_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT123), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n839_), .B2(new_n595_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(KEYINPUT61), .B(G155gat), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n850_), .A2(new_n852_), .A3(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n853_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(G1346gat));
  OR3_X1    g655(.A1(new_n839_), .A2(G162gat), .A3(new_n543_), .ZN(new_n857_));
  OAI21_X1  g656(.A(G162gat), .B1(new_n839_), .B2(new_n544_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(G1347gat));
  NOR4_X1   g658(.A1(new_n317_), .A2(new_n433_), .A3(new_n383_), .A4(new_n463_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n807_), .A2(new_n407_), .A3(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(KEYINPUT124), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n782_), .A2(new_n794_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n595_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n667_), .B1(new_n864_), .B2(new_n802_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT124), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n866_), .A3(new_n860_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n862_), .A2(new_n867_), .A3(G169gat), .ZN(new_n868_));
  XOR2_X1   g667(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n865_), .A2(new_n275_), .A3(new_n860_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n869_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n862_), .A2(new_n867_), .A3(G169gat), .A4(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n870_), .A2(new_n871_), .A3(new_n873_), .ZN(G1348gat));
  AOI21_X1  g673(.A(new_n317_), .B1(new_n864_), .B2(new_n802_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n408_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n580_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(new_n241_), .ZN(G1349gat));
  INV_X1    g677(.A(new_n876_), .ZN(new_n879_));
  AOI21_X1  g678(.A(G183gat), .B1(new_n879_), .B2(new_n596_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n280_), .A2(new_n281_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n876_), .A2(new_n595_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n880_), .B1(new_n881_), .B2(new_n882_), .ZN(G1350gat));
  OAI21_X1  g682(.A(G190gat), .B1(new_n876_), .B2(new_n544_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n603_), .A2(new_n279_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n876_), .B2(new_n885_), .ZN(G1351gat));
  NAND2_X1  g685(.A1(new_n837_), .A2(new_n384_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n875_), .A2(new_n888_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(new_n463_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(new_n217_), .ZN(G1352gat));
  NOR2_X1   g690(.A1(new_n889_), .A2(new_n580_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(new_n218_), .ZN(G1353gat));
  NOR3_X1   g692(.A1(KEYINPUT126), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(KEYINPUT126), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n595_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n875_), .A2(new_n888_), .A3(new_n898_), .ZN(new_n899_));
  MUX2_X1   g698(.A(new_n894_), .B(new_n897_), .S(new_n899_), .Z(G1354gat));
  NAND4_X1  g699(.A1(new_n807_), .A2(new_n610_), .A3(new_n635_), .A4(new_n888_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(G218gat), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n543_), .A2(G218gat), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n902_), .B1(new_n889_), .B2(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT127), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n902_), .B(KEYINPUT127), .C1(new_n889_), .C2(new_n904_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1355gat));
endmodule


