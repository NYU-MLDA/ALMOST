//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 1 1 0 0 1 1 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n583_, new_n584_, new_n585_, new_n586_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n645_, new_n646_, new_n647_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n654_, new_n655_, new_n656_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n796_,
    new_n797_, new_n799_, new_n800_, new_n801_, new_n802_, new_n804_,
    new_n805_, new_n806_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n825_, new_n826_,
    new_n827_, new_n829_, new_n830_, new_n831_, new_n833_, new_n834_,
    new_n836_, new_n838_, new_n839_, new_n841_, new_n842_, new_n844_,
    new_n845_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT88), .ZN(new_n203_));
  XOR2_X1   g002(.A(G113gat), .B(G120gat), .Z(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT89), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208_));
  XOR2_X1   g007(.A(new_n208_), .B(KEYINPUT92), .Z(new_n209_));
  AOI21_X1  g008(.A(new_n207_), .B1(new_n209_), .B2(KEYINPUT1), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n210_), .B1(KEYINPUT1), .B2(new_n209_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  OR2_X1    g011(.A1(G141gat), .A2(G148gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n216_), .B1(KEYINPUT3), .B2(new_n213_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n217_), .B1(KEYINPUT3), .B2(new_n213_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n212_), .A2(new_n215_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT93), .ZN(new_n220_));
  OAI221_X1 g019(.A(new_n209_), .B1(G155gat), .B2(G162gat), .C1(new_n218_), .C2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n214_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n206_), .A2(new_n222_), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n223_), .A2(KEYINPUT4), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT103), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G225gat), .A2(G233gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n214_), .A2(new_n221_), .A3(new_n205_), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n223_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT4), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n225_), .A2(new_n227_), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n229_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n231_), .B1(new_n227_), .B2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G1gat), .B(G29gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT0), .ZN(new_n235_));
  INV_X1    g034(.A(G57gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(G85gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n233_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT33), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n241_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n225_), .A2(new_n226_), .A3(new_n230_), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n244_), .B(new_n239_), .C1(new_n226_), .C2(new_n232_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n242_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT102), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G183gat), .A2(G190gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT23), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT83), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT23), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n251_), .A2(G183gat), .A3(G190gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n253_), .B1(G183gat), .B2(G190gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G169gat), .A2(G176gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT22), .B(G169gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT99), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n254_), .B(new_n255_), .C1(G176gat), .C2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT85), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n249_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n252_), .B(KEYINPUT86), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n255_), .A2(KEYINPUT24), .ZN(new_n264_));
  NOR2_X1   g063(.A1(G169gat), .A2(G176gat), .ZN(new_n265_));
  MUX2_X1   g064(.A(new_n264_), .B(KEYINPUT24), .S(new_n265_), .Z(new_n266_));
  XOR2_X1   g065(.A(KEYINPUT25), .B(G183gat), .Z(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT26), .B(G190gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n263_), .B(new_n266_), .C1(new_n267_), .C2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n259_), .A2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT96), .B(G204gat), .ZN(new_n272_));
  MUX2_X1   g071(.A(G204gat), .B(new_n272_), .S(G197gat), .Z(new_n273_));
  NOR2_X1   g072(.A1(new_n273_), .A2(KEYINPUT21), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G211gat), .B(G218gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT97), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n272_), .A2(G197gat), .ZN(new_n278_));
  INV_X1    g077(.A(G197gat), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n279_), .A2(G204gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT21), .B1(new_n278_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n277_), .A2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n276_), .A2(new_n273_), .A3(KEYINPUT21), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n271_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT84), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n256_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT22), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n286_), .B1(new_n288_), .B2(G169gat), .ZN(new_n289_));
  INV_X1    g088(.A(G176gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n255_), .B1(new_n287_), .B2(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n263_), .B1(G183gat), .B2(G190gat), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n292_), .B1(new_n293_), .B2(KEYINPUT87), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n294_), .B1(KEYINPUT87), .B2(new_n293_), .ZN(new_n295_));
  INV_X1    g094(.A(G190gat), .ZN(new_n296_));
  NOR3_X1   g095(.A1(new_n296_), .A2(KEYINPUT82), .A3(KEYINPUT26), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n297_), .B1(new_n268_), .B2(KEYINPUT82), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n253_), .B(new_n266_), .C1(new_n267_), .C2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n295_), .A2(new_n299_), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n285_), .B(KEYINPUT20), .C1(new_n300_), .C2(new_n284_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G226gat), .A2(G233gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT19), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT100), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n300_), .A2(new_n284_), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n306_), .B(KEYINPUT101), .Z(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT20), .B1(new_n271_), .B2(new_n284_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n308_), .A2(new_n303_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n305_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(G8gat), .B(G36gat), .Z(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT18), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G64gat), .B(G92gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n247_), .B1(new_n310_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n310_), .A2(new_n314_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n317_), .B1(KEYINPUT102), .B2(new_n316_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n314_), .A2(KEYINPUT32), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n319_), .B(KEYINPUT104), .Z(new_n320_));
  NAND2_X1  g119(.A1(new_n310_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT105), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n233_), .A2(new_n239_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n240_), .A2(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n301_), .A2(new_n303_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n308_), .B(KEYINPUT106), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n307_), .A2(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n325_), .B1(new_n327_), .B2(new_n303_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n324_), .B1(new_n328_), .B2(new_n319_), .ZN(new_n329_));
  OAI22_X1  g128(.A1(new_n246_), .A2(new_n318_), .B1(new_n322_), .B2(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n222_), .A2(KEYINPUT29), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT28), .ZN(new_n332_));
  XOR2_X1   g131(.A(G22gat), .B(G50gat), .Z(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n222_), .A2(KEYINPUT29), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n284_), .ZN(new_n336_));
  INV_X1    g135(.A(G228gat), .ZN(new_n337_));
  INV_X1    g136(.A(G233gat), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n338_), .A2(KEYINPUT94), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(KEYINPUT94), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n337_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT95), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n336_), .B(new_n342_), .Z(new_n343_));
  XNOR2_X1  g142(.A(G78gat), .B(G106gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n334_), .B1(new_n345_), .B2(KEYINPUT98), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n346_), .B1(KEYINPUT98), .B2(new_n345_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n345_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT98), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(new_n349_), .A3(new_n334_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n347_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n300_), .B(KEYINPUT30), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G71gat), .B(G99gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(G43gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G227gat), .A2(G233gat), .ZN(new_n356_));
  INV_X1    g155(.A(G15gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n355_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n353_), .B(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n206_), .B(KEYINPUT31), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT90), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT91), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n364_), .A2(new_n365_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT91), .B1(new_n361_), .B2(new_n363_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n352_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n330_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT27), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n318_), .A2(new_n371_), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n316_), .B(KEYINPUT27), .C1(new_n314_), .C2(new_n328_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n368_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n352_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n351_), .A2(new_n368_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n324_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n374_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n370_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G230gat), .A2(G233gat), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT67), .ZN(new_n383_));
  INV_X1    g182(.A(G64gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(G57gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n236_), .A2(G64gat), .ZN(new_n386_));
  AOI21_X1  g185(.A(KEYINPUT11), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G71gat), .B(G78gat), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n383_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  AND2_X1   g188(.A1(G71gat), .A2(G78gat), .ZN(new_n390_));
  NOR2_X1   g189(.A1(G71gat), .A2(G78gat), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G57gat), .B(G64gat), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n392_), .B(KEYINPUT67), .C1(new_n393_), .C2(KEYINPUT11), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(KEYINPUT11), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n389_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n395_), .B1(new_n389_), .B2(new_n394_), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT68), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n395_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT11), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n236_), .A2(G64gat), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n384_), .A2(G57gat), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n400_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(KEYINPUT67), .B1(new_n403_), .B2(new_n392_), .ZN(new_n404_));
  NOR3_X1   g203(.A1(new_n387_), .A2(new_n383_), .A3(new_n388_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n399_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT68), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n389_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n406_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n398_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(G99gat), .ZN(new_n411_));
  INV_X1    g210(.A(G106gat), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n412_), .A3(KEYINPUT65), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT65), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n414_), .B1(G99gat), .B2(G106gat), .ZN(new_n415_));
  OR2_X1    g214(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n416_));
  NAND2_X1  g215(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n413_), .A2(new_n415_), .A3(new_n416_), .A4(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n419_));
  OR2_X1    g218(.A1(KEYINPUT64), .A2(KEYINPUT6), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G99gat), .A2(G106gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(KEYINPUT64), .A2(KEYINPUT6), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n420_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n421_), .B1(new_n420_), .B2(new_n422_), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n418_), .B(new_n419_), .C1(new_n423_), .C2(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(G85gat), .B(G92gat), .Z(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(KEYINPUT8), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(G92gat), .ZN(new_n428_));
  NOR3_X1   g227(.A1(new_n238_), .A2(new_n428_), .A3(KEYINPUT9), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n429_), .B1(new_n426_), .B2(KEYINPUT9), .ZN(new_n430_));
  XNOR2_X1  g229(.A(KEYINPUT10), .B(G99gat), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n431_), .A2(G106gat), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n430_), .B(new_n432_), .C1(new_n424_), .C2(new_n423_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n427_), .A2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT8), .B1(new_n425_), .B2(new_n426_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n410_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n410_), .A2(new_n436_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n382_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  XOR2_X1   g239(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n441_));
  OAI21_X1  g240(.A(new_n441_), .B1(new_n410_), .B2(new_n436_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n396_), .A2(new_n397_), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n443_), .B(KEYINPUT12), .C1(new_n434_), .C2(new_n435_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n442_), .A2(new_n381_), .A3(new_n437_), .A4(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n440_), .A2(new_n445_), .ZN(new_n446_));
  XOR2_X1   g245(.A(G120gat), .B(G148gat), .Z(new_n447_));
  XNOR2_X1  g246(.A(G176gat), .B(G204gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n449_), .B(new_n450_), .Z(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT70), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n446_), .B(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT13), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT13), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n454_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  OR2_X1    g258(.A1(new_n357_), .A2(G22gat), .ZN(new_n460_));
  INV_X1    g259(.A(G1gat), .ZN(new_n461_));
  INV_X1    g260(.A(G8gat), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT14), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n357_), .A2(G22gat), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n460_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  OR2_X1    g264(.A1(new_n465_), .A2(KEYINPUT78), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(KEYINPUT78), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(G1gat), .B(G8gat), .Z(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n466_), .A2(new_n469_), .A3(new_n467_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G29gat), .B(G36gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G43gat), .B(G50gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n473_), .B(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n477_), .A2(G229gat), .A3(G233gat), .ZN(new_n478_));
  XOR2_X1   g277(.A(new_n476_), .B(KEYINPUT15), .Z(new_n479_));
  OR2_X1    g278(.A1(new_n479_), .A2(new_n473_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n473_), .A2(new_n476_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G229gat), .A2(G233gat), .ZN(new_n482_));
  XOR2_X1   g281(.A(new_n482_), .B(KEYINPUT81), .Z(new_n483_));
  NAND3_X1  g282(.A1(new_n480_), .A2(new_n481_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n478_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G113gat), .B(G141gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G169gat), .B(G197gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n485_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n488_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n478_), .A2(new_n484_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n459_), .A2(new_n492_), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n380_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G232gat), .A2(G233gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT34), .ZN(new_n496_));
  OAI22_X1  g295(.A1(new_n436_), .A2(new_n479_), .B1(KEYINPUT35), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n435_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n498_), .A2(new_n476_), .A3(new_n427_), .A4(new_n433_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT72), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT72), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n436_), .A2(new_n501_), .A3(new_n476_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n497_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n496_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT35), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n503_), .A2(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT74), .B1(new_n503_), .B2(new_n507_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n497_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n502_), .A2(new_n500_), .ZN(new_n511_));
  AND4_X1   g310(.A1(KEYINPUT74), .A2(new_n510_), .A3(new_n511_), .A4(new_n507_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n508_), .B1(new_n509_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT76), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G190gat), .B(G218gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT73), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G134gat), .B(G162gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT36), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n503_), .A2(new_n507_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n510_), .A2(new_n511_), .A3(new_n507_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT74), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n503_), .A2(KEYINPUT74), .A3(new_n507_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n521_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT76), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n520_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n518_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n529_), .A2(KEYINPUT36), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n508_), .B(new_n530_), .C1(new_n509_), .C2(new_n512_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT75), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n526_), .A2(KEYINPUT75), .A3(new_n530_), .ZN(new_n534_));
  AOI22_X1  g333(.A1(new_n514_), .A2(new_n528_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(KEYINPUT77), .B(KEYINPUT37), .Z(new_n536_));
  NAND2_X1  g335(.A1(new_n513_), .A2(new_n519_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n531_), .A2(new_n532_), .ZN(new_n538_));
  AOI21_X1  g337(.A(KEYINPUT75), .B1(new_n526_), .B2(new_n530_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n537_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n535_), .A2(new_n536_), .B1(new_n540_), .B2(KEYINPUT37), .ZN(new_n541_));
  AND2_X1   g340(.A1(G231gat), .A2(G233gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n473_), .B(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n443_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n544_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n407_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT80), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n545_), .A2(KEYINPUT68), .A3(new_n546_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n548_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G127gat), .B(G155gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT16), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT79), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G183gat), .B(G211gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT17), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n551_), .A2(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n549_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n560_));
  OAI22_X1  g359(.A1(new_n559_), .A2(new_n560_), .B1(new_n557_), .B2(new_n556_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n556_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n547_), .A2(KEYINPUT17), .A3(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n541_), .A2(new_n565_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n494_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n567_), .A2(new_n461_), .A3(new_n324_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT38), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n565_), .A2(new_n535_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n494_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n324_), .ZN(new_n572_));
  OAI21_X1  g371(.A(G1gat), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n569_), .A2(new_n573_), .ZN(G1324gat));
  NAND2_X1  g373(.A1(new_n372_), .A2(new_n373_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n567_), .A2(new_n462_), .A3(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(G8gat), .B1(new_n571_), .B2(new_n374_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n577_), .A2(KEYINPUT39), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n577_), .A2(KEYINPUT39), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n576_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT40), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(G1325gat));
  OAI21_X1  g381(.A(G15gat), .B1(new_n571_), .B2(new_n375_), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n583_), .A2(KEYINPUT41), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(KEYINPUT41), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n567_), .A2(new_n357_), .A3(new_n368_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n584_), .A2(new_n585_), .A3(new_n586_), .ZN(G1326gat));
  OAI21_X1  g386(.A(G22gat), .B1(new_n571_), .B2(new_n351_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT42), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n351_), .A2(G22gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT107), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n567_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n589_), .A2(new_n592_), .ZN(G1327gat));
  INV_X1    g392(.A(new_n535_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n564_), .A2(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n494_), .A2(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(G29gat), .B1(new_n596_), .B2(new_n324_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT109), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT44), .ZN(new_n599_));
  OAI21_X1  g398(.A(KEYINPUT108), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT43), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n380_), .A2(new_n601_), .A3(new_n541_), .ZN(new_n602_));
  AOI22_X1  g401(.A1(new_n330_), .A2(new_n369_), .B1(new_n374_), .B2(new_n378_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n535_), .A2(new_n536_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n540_), .A2(KEYINPUT37), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(KEYINPUT43), .B1(new_n603_), .B2(new_n606_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n602_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n565_), .A2(new_n493_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n600_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n609_), .B1(new_n602_), .B2(new_n607_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n598_), .B1(new_n611_), .B2(KEYINPUT108), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n610_), .B1(new_n612_), .B2(KEYINPUT44), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n324_), .A2(G29gat), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n597_), .B1(new_n613_), .B2(new_n614_), .ZN(G1328gat));
  INV_X1    g414(.A(G36gat), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n596_), .A2(new_n616_), .A3(new_n575_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT45), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n613_), .A2(new_n575_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n618_), .B(KEYINPUT46), .C1(new_n619_), .C2(new_n616_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT46), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n617_), .B(KEYINPUT45), .Z(new_n622_));
  AOI21_X1  g421(.A(new_n616_), .B1(new_n613_), .B2(new_n575_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n621_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n620_), .A2(new_n624_), .ZN(G1329gat));
  AOI21_X1  g424(.A(G43gat), .B1(new_n596_), .B2(new_n368_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n368_), .A2(G43gat), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n626_), .B1(new_n613_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT47), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(G1330gat));
  INV_X1    g429(.A(G50gat), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n596_), .A2(new_n631_), .A3(new_n352_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n613_), .A2(new_n352_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n633_), .A2(KEYINPUT110), .ZN(new_n634_));
  OAI21_X1  g433(.A(G50gat), .B1(new_n633_), .B2(KEYINPUT110), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n632_), .B1(new_n634_), .B2(new_n635_), .ZN(G1331gat));
  NOR3_X1   g435(.A1(new_n603_), .A2(new_n492_), .A3(new_n459_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(new_n570_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n638_), .A2(new_n236_), .A3(new_n572_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT112), .Z(new_n640_));
  NAND2_X1  g439(.A1(new_n637_), .A2(new_n566_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n236_), .B1(new_n641_), .B2(new_n572_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT111), .Z(new_n643_));
  NOR2_X1   g442(.A1(new_n640_), .A2(new_n643_), .ZN(G1332gat));
  OAI21_X1  g443(.A(G64gat), .B1(new_n638_), .B2(new_n374_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT48), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n575_), .A2(new_n384_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n646_), .B1(new_n641_), .B2(new_n647_), .ZN(G1333gat));
  OAI21_X1  g447(.A(G71gat), .B1(new_n638_), .B2(new_n375_), .ZN(new_n649_));
  XOR2_X1   g448(.A(KEYINPUT113), .B(KEYINPUT49), .Z(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n375_), .A2(G71gat), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n651_), .B1(new_n641_), .B2(new_n652_), .ZN(G1334gat));
  OAI21_X1  g452(.A(G78gat), .B1(new_n638_), .B2(new_n351_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT50), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n351_), .A2(G78gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n655_), .B1(new_n641_), .B2(new_n656_), .ZN(G1335gat));
  NOR3_X1   g456(.A1(new_n564_), .A2(new_n492_), .A3(new_n459_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT114), .Z(new_n659_));
  AOI21_X1  g458(.A(new_n659_), .B1(new_n602_), .B2(new_n607_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G85gat), .B1(new_n661_), .B2(new_n572_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n637_), .A2(new_n595_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n664_), .A2(new_n238_), .A3(new_n324_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n662_), .A2(new_n665_), .ZN(G1336gat));
  OAI21_X1  g465(.A(G92gat), .B1(new_n661_), .B2(new_n374_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n664_), .A2(new_n428_), .A3(new_n575_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1337gat));
  AOI21_X1  g468(.A(new_n411_), .B1(new_n660_), .B2(new_n368_), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n663_), .A2(new_n431_), .A3(new_n375_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g472(.A1(new_n664_), .A2(new_n412_), .A3(new_n352_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n412_), .B1(new_n660_), .B2(new_n352_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT52), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n675_), .A2(new_n676_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n674_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g479(.A1(new_n575_), .A2(new_n572_), .A3(new_n377_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n477_), .A2(new_n483_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n480_), .A2(new_n481_), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n683_), .B(new_n488_), .C1(new_n684_), .C2(new_n483_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n685_), .A2(new_n491_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n455_), .A2(new_n686_), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n442_), .A2(new_n437_), .A3(new_n444_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n688_), .A2(KEYINPUT116), .A3(KEYINPUT55), .A4(new_n381_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT116), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT55), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n690_), .B1(new_n445_), .B2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n689_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n445_), .A2(new_n691_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT115), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n437_), .A2(new_n444_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n696_), .B2(new_n442_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n442_), .A2(new_n695_), .A3(new_n437_), .A4(new_n444_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n382_), .B1(new_n697_), .B2(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n693_), .A2(new_n694_), .A3(new_n700_), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n701_), .A2(KEYINPUT56), .A3(new_n452_), .ZN(new_n702_));
  AOI21_X1  g501(.A(KEYINPUT56), .B1(new_n701_), .B2(new_n452_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n702_), .A2(new_n703_), .A3(KEYINPUT117), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n701_), .A2(new_n452_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT56), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n705_), .A2(KEYINPUT117), .A3(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n440_), .A2(new_n445_), .A3(new_n451_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n492_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n707_), .A2(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n687_), .B1(new_n704_), .B2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n712_), .A2(KEYINPUT57), .A3(new_n594_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n686_), .A2(new_n708_), .ZN(new_n714_));
  OAI211_X1 g513(.A(KEYINPUT58), .B(new_n714_), .C1(new_n702_), .C2(new_n703_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT118), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n705_), .A2(new_n706_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n701_), .A2(KEYINPUT56), .A3(new_n452_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n720_), .A2(KEYINPUT118), .A3(KEYINPUT58), .A4(new_n714_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n714_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT58), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n717_), .A2(new_n721_), .A3(new_n541_), .A4(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n713_), .A2(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT57), .B1(new_n712_), .B2(new_n594_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n565_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n492_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n528_), .A2(new_n514_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n533_), .A2(new_n534_), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n730_), .A2(new_n731_), .A3(new_n536_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT37), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n731_), .B2(new_n537_), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n564_), .B(new_n729_), .C1(new_n732_), .C2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT54), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n606_), .A2(KEYINPUT54), .A3(new_n564_), .A4(new_n729_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n728_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT119), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT119), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n728_), .A2(new_n740_), .A3(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n682_), .B1(new_n742_), .B2(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(G113gat), .B1(new_n745_), .B2(new_n492_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT120), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT59), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n745_), .B2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n743_), .B1(new_n728_), .B2(new_n740_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT57), .ZN(new_n751_));
  INV_X1    g550(.A(new_n687_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT117), .ZN(new_n753_));
  AOI211_X1 g552(.A(new_n753_), .B(KEYINPUT56), .C1(new_n701_), .C2(new_n452_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n754_), .A2(new_n709_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n718_), .A2(new_n753_), .A3(new_n719_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n752_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n751_), .B1(new_n757_), .B2(new_n535_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(new_n713_), .A3(new_n725_), .ZN(new_n759_));
  AOI211_X1 g558(.A(KEYINPUT119), .B(new_n739_), .C1(new_n759_), .C2(new_n565_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n681_), .B1(new_n750_), .B2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(KEYINPUT120), .A3(KEYINPUT59), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n749_), .A2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n741_), .A2(new_n748_), .A3(new_n681_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n492_), .A2(KEYINPUT121), .A3(G113gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n767_), .B1(KEYINPUT121), .B2(G113gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n746_), .B1(new_n766_), .B2(new_n768_), .ZN(G1340gat));
  INV_X1    g568(.A(new_n459_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n761_), .A2(KEYINPUT120), .A3(KEYINPUT59), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT120), .B1(new_n761_), .B2(KEYINPUT59), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n770_), .B(new_n764_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT122), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n763_), .A2(KEYINPUT122), .A3(new_n770_), .A4(new_n764_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(G120gat), .A3(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT60), .ZN(new_n778_));
  INV_X1    g577(.A(G120gat), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n770_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n780_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n745_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n777_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT123), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT123), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n777_), .A2(new_n785_), .A3(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1341gat));
  OAI21_X1  g586(.A(G127gat), .B1(new_n765_), .B2(new_n565_), .ZN(new_n788_));
  INV_X1    g587(.A(G127gat), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n745_), .A2(new_n789_), .A3(new_n564_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT124), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n788_), .A2(KEYINPUT124), .A3(new_n790_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(G1342gat));
  OAI21_X1  g594(.A(G134gat), .B1(new_n765_), .B2(new_n606_), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n594_), .A2(G134gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n761_), .B2(new_n797_), .ZN(G1343gat));
  AOI21_X1  g597(.A(new_n376_), .B1(new_n742_), .B2(new_n744_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n575_), .A2(new_n572_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(new_n492_), .A3(new_n800_), .ZN(new_n801_));
  XOR2_X1   g600(.A(KEYINPUT125), .B(G141gat), .Z(new_n802_));
  XNOR2_X1  g601(.A(new_n801_), .B(new_n802_), .ZN(G1344gat));
  NAND2_X1  g602(.A1(new_n799_), .A2(new_n800_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n804_), .A2(new_n459_), .ZN(new_n805_));
  XOR2_X1   g604(.A(KEYINPUT126), .B(G148gat), .Z(new_n806_));
  XNOR2_X1  g605(.A(new_n805_), .B(new_n806_), .ZN(G1345gat));
  NOR2_X1   g606(.A1(new_n804_), .A2(new_n565_), .ZN(new_n808_));
  XOR2_X1   g607(.A(KEYINPUT61), .B(G155gat), .Z(new_n809_));
  XNOR2_X1  g608(.A(new_n808_), .B(new_n809_), .ZN(G1346gat));
  OAI21_X1  g609(.A(G162gat), .B1(new_n804_), .B2(new_n606_), .ZN(new_n811_));
  OR2_X1    g610(.A1(new_n594_), .A2(G162gat), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n804_), .B2(new_n812_), .ZN(G1347gat));
  INV_X1    g612(.A(KEYINPUT127), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n374_), .A2(new_n324_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n368_), .ZN(new_n816_));
  AOI211_X1 g615(.A(new_n352_), .B(new_n816_), .C1(new_n728_), .C2(new_n740_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n492_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(G169gat), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n814_), .B1(new_n819_), .B2(KEYINPUT62), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(KEYINPUT62), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n819_), .A2(new_n814_), .A3(KEYINPUT62), .ZN(new_n823_));
  OAI22_X1  g622(.A1(new_n822_), .A2(new_n823_), .B1(new_n258_), .B2(new_n818_), .ZN(G1348gat));
  AOI21_X1  g623(.A(G176gat), .B1(new_n817_), .B2(new_n770_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n352_), .B1(new_n742_), .B2(new_n744_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n816_), .A2(new_n290_), .A3(new_n459_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n825_), .B1(new_n826_), .B2(new_n827_), .ZN(G1349gat));
  NAND4_X1  g627(.A1(new_n826_), .A2(new_n368_), .A3(new_n564_), .A4(new_n815_), .ZN(new_n829_));
  INV_X1    g628(.A(G183gat), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n564_), .A2(new_n267_), .ZN(new_n831_));
  AOI22_X1  g630(.A1(new_n829_), .A2(new_n830_), .B1(new_n817_), .B2(new_n831_), .ZN(G1350gat));
  NAND3_X1  g631(.A1(new_n817_), .A2(new_n268_), .A3(new_n535_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n817_), .A2(new_n541_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n834_), .B2(new_n296_), .ZN(G1351gat));
  NAND3_X1  g634(.A1(new_n799_), .A2(new_n492_), .A3(new_n815_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g636(.A1(new_n799_), .A2(new_n815_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n838_), .A2(new_n459_), .ZN(new_n839_));
  MUX2_X1   g638(.A(G204gat), .B(new_n272_), .S(new_n839_), .Z(G1353gat));
  AOI211_X1 g639(.A(new_n565_), .B(new_n838_), .C1(KEYINPUT63), .C2(G211gat), .ZN(new_n841_));
  NOR2_X1   g640(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n841_), .B(new_n842_), .ZN(G1354gat));
  OAI21_X1  g642(.A(G218gat), .B1(new_n838_), .B2(new_n606_), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n594_), .A2(G218gat), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n838_), .B2(new_n845_), .ZN(G1355gat));
endmodule


