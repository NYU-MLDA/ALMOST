//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n845_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n879_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n204_));
  XOR2_X1   g003(.A(G71gat), .B(G78gat), .Z(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n204_), .A2(new_n205_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(KEYINPUT10), .B(G99gat), .Z(new_n209_));
  INV_X1    g008(.A(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(G85gat), .B(G92gat), .Z(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT9), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G99gat), .A3(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G85gat), .ZN(new_n219_));
  INV_X1    g018(.A(G92gat), .ZN(new_n220_));
  OR3_X1    g019(.A1(new_n219_), .A2(new_n220_), .A3(KEYINPUT9), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n211_), .A2(new_n213_), .A3(new_n218_), .A4(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT8), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n218_), .A2(KEYINPUT64), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G99gat), .A2(G106gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT7), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT64), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n215_), .A2(new_n217_), .A3(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n224_), .A2(new_n226_), .A3(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n223_), .B1(new_n229_), .B2(new_n212_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n212_), .A2(new_n223_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n231_), .B1(new_n218_), .B2(new_n226_), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n208_), .B(new_n222_), .C1(new_n230_), .C2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(new_n233_), .B(KEYINPUT65), .Z(new_n234_));
  OAI21_X1  g033(.A(new_n222_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n208_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n234_), .A2(new_n237_), .ZN(new_n238_));
  AND2_X1   g037(.A1(G230gat), .A2(G233gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n235_), .A2(KEYINPUT66), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n242_), .B(new_n222_), .C1(new_n230_), .C2(new_n232_), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n241_), .A2(KEYINPUT12), .A3(new_n236_), .A4(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT12), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n237_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n233_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n247_), .A2(new_n239_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n244_), .A2(new_n246_), .A3(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n240_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G120gat), .B(G148gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT5), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G176gat), .B(G204gat), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n252_), .B(new_n253_), .Z(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT67), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n250_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n254_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n240_), .A2(new_n249_), .A3(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(KEYINPUT68), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n250_), .A2(new_n260_), .A3(new_n255_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT13), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT13), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n259_), .A2(new_n264_), .A3(new_n261_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G29gat), .B(G36gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT71), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G43gat), .B(G50gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT15), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G15gat), .B(G22gat), .ZN(new_n274_));
  INV_X1    g073(.A(G1gat), .ZN(new_n275_));
  INV_X1    g074(.A(G8gat), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT14), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n274_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G1gat), .B(G8gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n273_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n280_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n272_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G229gat), .A2(G233gat), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n281_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n272_), .B(new_n280_), .ZN(new_n286_));
  NOR3_X1   g085(.A1(new_n286_), .A2(KEYINPUT77), .A3(new_n284_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT77), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n272_), .B(new_n282_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n284_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n288_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n285_), .B1(new_n287_), .B2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G113gat), .B(G141gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT78), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G169gat), .B(G197gat), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n294_), .B(new_n295_), .Z(new_n296_));
  NAND2_X1  g095(.A1(new_n292_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n296_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n285_), .B(new_n298_), .C1(new_n287_), .C2(new_n291_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n263_), .A2(KEYINPUT69), .A3(new_n265_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n268_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT25), .B(G183gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT26), .B(G190gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307_));
  AOI22_X1  g106(.A1(new_n303_), .A2(new_n304_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  NOR3_X1   g107(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G183gat), .A2(G190gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT23), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT23), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n312_), .A2(G183gat), .A3(G190gat), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n309_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n308_), .A2(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(G183gat), .A2(G190gat), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n316_), .B1(new_n312_), .B2(new_n310_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n317_), .B1(new_n312_), .B2(new_n310_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(G169gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n315_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT30), .ZN(new_n323_));
  INV_X1    g122(.A(G99gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(KEYINPUT79), .B(G43gat), .Z(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n323_), .B(G99gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n326_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G227gat), .A2(G233gat), .ZN(new_n332_));
  INV_X1    g131(.A(G15gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(G71gat), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n331_), .A2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n328_), .A2(new_n330_), .A3(new_n335_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n337_), .A2(KEYINPUT80), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT31), .ZN(new_n340_));
  XOR2_X1   g139(.A(G127gat), .B(G134gat), .Z(new_n341_));
  XOR2_X1   g140(.A(G113gat), .B(G120gat), .Z(new_n342_));
  XOR2_X1   g141(.A(new_n341_), .B(new_n342_), .Z(new_n343_));
  INV_X1    g142(.A(KEYINPUT31), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n337_), .A2(KEYINPUT80), .A3(new_n344_), .A4(new_n338_), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n340_), .A2(new_n343_), .A3(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n343_), .B1(new_n340_), .B2(new_n345_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT27), .ZN(new_n349_));
  NOR2_X1   g148(.A1(G197gat), .A2(G204gat), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT86), .ZN(new_n351_));
  INV_X1    g150(.A(G204gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(KEYINPUT86), .A2(G204gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n350_), .B1(new_n355_), .B2(G197gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G211gat), .B(G218gat), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n356_), .A2(KEYINPUT21), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(G197gat), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n353_), .A2(new_n360_), .A3(new_n354_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT87), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT21), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n363_), .B1(G197gat), .B2(G204gat), .ZN(new_n364_));
  AND3_X1   g163(.A1(new_n361_), .A2(new_n362_), .A3(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n362_), .B1(new_n361_), .B2(new_n364_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n357_), .B1(new_n356_), .B2(KEYINPUT21), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n359_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(new_n322_), .ZN(new_n370_));
  AOI22_X1  g169(.A1(new_n314_), .A2(new_n308_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n371_), .B(new_n359_), .C1(new_n367_), .C2(new_n368_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(KEYINPUT20), .A3(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G226gat), .A2(G233gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n373_), .A2(new_n376_), .ZN(new_n377_));
  XOR2_X1   g176(.A(G8gat), .B(G36gat), .Z(new_n378_));
  XNOR2_X1  g177(.A(G64gat), .B(G92gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n376_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n370_), .A2(KEYINPUT20), .A3(new_n372_), .A4(new_n383_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n377_), .A2(new_n382_), .A3(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n382_), .B1(new_n377_), .B2(new_n384_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n349_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT100), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT100), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n389_), .B(new_n349_), .C1(new_n385_), .C2(new_n386_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n382_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT98), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n370_), .A2(new_n392_), .A3(new_n372_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n373_), .A2(new_n393_), .A3(new_n376_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n373_), .B1(new_n376_), .B2(new_n393_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n391_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n396_), .A2(KEYINPUT27), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n377_), .A2(new_n382_), .A3(new_n384_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT99), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  AOI22_X1  g199(.A1(new_n388_), .A2(new_n390_), .B1(new_n397_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G22gat), .B(G50gat), .ZN(new_n403_));
  XOR2_X1   g202(.A(G141gat), .B(G148gat), .Z(new_n404_));
  NAND2_X1  g203(.A1(G155gat), .A2(G162gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT81), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT81), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n407_), .A2(G155gat), .A3(G162gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT1), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT82), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT1), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n406_), .A2(new_n408_), .A3(new_n411_), .A4(new_n412_), .ZN(new_n413_));
  OR2_X1    g212(.A1(G155gat), .A2(G162gat), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n410_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n406_), .A2(new_n408_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n411_), .B1(new_n416_), .B2(new_n412_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n404_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(G141gat), .ZN(new_n419_));
  INV_X1    g218(.A(G148gat), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT83), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT2), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT2), .ZN(new_n423_));
  OAI211_X1 g222(.A(KEYINPUT83), .B(new_n423_), .C1(new_n419_), .C2(new_n420_), .ZN(new_n424_));
  OR3_X1    g223(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n422_), .A2(new_n424_), .A3(new_n425_), .A4(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(new_n409_), .A3(new_n414_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n418_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT84), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT84), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n418_), .A2(new_n431_), .A3(new_n428_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT28), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT29), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n433_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n434_), .B1(new_n433_), .B2(new_n435_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n403_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n438_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n403_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(new_n436_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n429_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n369_), .B1(new_n444_), .B2(new_n435_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT88), .ZN(new_n446_));
  INV_X1    g245(.A(G233gat), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n447_), .A2(KEYINPUT85), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(KEYINPUT85), .ZN(new_n449_));
  OAI21_X1  g248(.A(G228gat), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n445_), .A2(new_n446_), .A3(new_n451_), .ZN(new_n452_));
  OAI221_X1 g251(.A(new_n357_), .B1(new_n356_), .B2(KEYINPUT21), .C1(new_n365_), .C2(new_n366_), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n429_), .A2(KEYINPUT29), .B1(new_n453_), .B2(new_n359_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT88), .B1(new_n454_), .B2(new_n450_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n452_), .A2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G78gat), .B(G106gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT89), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n369_), .B(new_n450_), .C1(new_n433_), .C2(new_n435_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n456_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n459_), .B1(new_n456_), .B2(new_n460_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n443_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n456_), .A2(new_n460_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(new_n458_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n466_), .A2(new_n442_), .A3(new_n439_), .A4(new_n461_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n464_), .A2(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n402_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n430_), .A2(new_n432_), .A3(new_n343_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n470_), .A2(KEYINPUT4), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G225gat), .A2(G233gat), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT93), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT4), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT92), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n476_), .B1(new_n429_), .B2(new_n343_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n470_), .A2(new_n478_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n430_), .A2(KEYINPUT92), .A3(new_n432_), .A4(new_n343_), .ZN(new_n480_));
  AOI211_X1 g279(.A(new_n474_), .B(new_n475_), .C1(new_n479_), .C2(new_n480_), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n418_), .A2(new_n431_), .A3(new_n428_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n431_), .B1(new_n418_), .B2(new_n428_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n343_), .ZN(new_n484_));
  NOR3_X1   g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n480_), .B1(new_n485_), .B2(new_n477_), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT93), .B1(new_n486_), .B2(KEYINPUT4), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n473_), .B1(new_n481_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n472_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G1gat), .B(G29gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(G85gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT0), .B(G57gat), .ZN(new_n493_));
  XOR2_X1   g292(.A(new_n492_), .B(new_n493_), .Z(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n489_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n496_), .A2(new_n495_), .ZN(new_n497_));
  AOI22_X1  g296(.A1(new_n490_), .A2(new_n495_), .B1(new_n488_), .B2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n348_), .A2(new_n469_), .A3(new_n498_), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n346_), .A2(new_n347_), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n385_), .A2(new_n386_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n488_), .A2(new_n497_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT33), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n501_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n472_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n471_), .A2(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n506_), .B1(new_n481_), .B2(new_n487_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT96), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n494_), .B1(new_n486_), .B2(new_n505_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT95), .ZN(new_n511_));
  OAI211_X1 g310(.A(KEYINPUT96), .B(new_n506_), .C1(new_n481_), .C2(new_n487_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n509_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n488_), .A2(KEYINPUT33), .A3(new_n497_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT94), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n488_), .A2(new_n497_), .A3(KEYINPUT94), .A4(KEYINPUT33), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n504_), .A2(new_n513_), .A3(new_n516_), .A4(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n473_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n486_), .A2(KEYINPUT4), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(new_n474_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n486_), .A2(KEYINPUT93), .A3(KEYINPUT4), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n519_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n495_), .B1(new_n523_), .B2(new_n496_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(new_n502_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n382_), .A2(KEYINPUT32), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n377_), .A2(new_n384_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT97), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n526_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  OR3_X1    g328(.A1(new_n394_), .A2(new_n395_), .A3(new_n526_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n527_), .A2(KEYINPUT97), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n529_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n525_), .A2(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n468_), .B1(new_n518_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n388_), .A2(new_n390_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n385_), .A2(new_n399_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n398_), .A2(KEYINPUT99), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n536_), .A2(new_n396_), .A3(KEYINPUT27), .A4(new_n537_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n535_), .A2(new_n467_), .A3(new_n464_), .A4(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT101), .B1(new_n525_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT101), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n498_), .A2(new_n468_), .A3(new_n541_), .A4(new_n401_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n500_), .B1(new_n534_), .B2(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n302_), .B1(new_n499_), .B2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n273_), .A2(new_n241_), .A3(new_n243_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n272_), .B(new_n222_), .C1(new_n230_), .C2(new_n232_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT35), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G190gat), .B(G218gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT73), .ZN(new_n551_));
  XOR2_X1   g350(.A(G134gat), .B(G162gat), .Z(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  AOI22_X1  g353(.A1(new_n548_), .A2(new_n549_), .B1(KEYINPUT36), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G232gat), .A2(G233gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT35), .ZN(new_n557_));
  XOR2_X1   g356(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n558_));
  XOR2_X1   g357(.A(new_n557_), .B(new_n558_), .Z(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT72), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n560_), .B1(new_n548_), .B2(new_n561_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n546_), .A2(KEYINPUT72), .A3(new_n547_), .A4(new_n559_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n555_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n554_), .A2(KEYINPUT36), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n565_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n555_), .A2(new_n562_), .A3(new_n567_), .A4(new_n563_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT74), .B(KEYINPUT37), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n566_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n569_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT17), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n280_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(new_n208_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n576_), .A2(KEYINPUT75), .ZN(new_n577_));
  XOR2_X1   g376(.A(G127gat), .B(G155gat), .Z(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT16), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G183gat), .B(G211gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n576_), .A2(KEYINPUT75), .ZN(new_n582_));
  OR4_X1    g381(.A1(new_n573_), .A2(new_n577_), .A3(new_n581_), .A4(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n581_), .B(KEYINPUT17), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n576_), .A2(new_n584_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n585_), .A2(KEYINPUT76), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(KEYINPUT76), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n583_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n572_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n545_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(KEYINPUT102), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT102), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n545_), .A2(new_n592_), .A3(new_n589_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n498_), .A2(G1gat), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(KEYINPUT103), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT103), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n595_), .A2(new_n599_), .A3(new_n596_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT38), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n302_), .A2(KEYINPUT104), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT104), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n268_), .A2(new_n605_), .A3(new_n300_), .A4(new_n301_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n588_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n566_), .A2(new_n568_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT105), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n609_), .B1(new_n544_), .B2(new_n499_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n607_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(new_n525_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(G1gat), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n598_), .A2(KEYINPUT38), .A3(new_n600_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n603_), .A2(new_n613_), .A3(new_n614_), .ZN(G1324gat));
  NAND3_X1  g414(.A1(new_n607_), .A2(new_n402_), .A3(new_n610_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT39), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n616_), .A2(new_n617_), .A3(G8gat), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n617_), .B1(new_n616_), .B2(G8gat), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n402_), .A2(new_n276_), .ZN(new_n620_));
  OAI22_X1  g419(.A1(new_n618_), .A2(new_n619_), .B1(new_n594_), .B2(new_n620_), .ZN(new_n621_));
  XOR2_X1   g420(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(G1325gat));
  NAND3_X1  g422(.A1(new_n595_), .A2(new_n333_), .A3(new_n348_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n611_), .A2(new_n348_), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n625_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT41), .B1(new_n625_), .B2(G15gat), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n624_), .B1(new_n626_), .B2(new_n627_), .ZN(G1326gat));
  INV_X1    g427(.A(new_n468_), .ZN(new_n629_));
  OR3_X1    g428(.A1(new_n594_), .A2(G22gat), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n611_), .A2(new_n468_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(G22gat), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n632_), .A2(KEYINPUT42), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(KEYINPUT42), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n630_), .B1(new_n633_), .B2(new_n634_), .ZN(G1327gat));
  INV_X1    g434(.A(new_n588_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n636_), .A2(new_n608_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n637_), .B(KEYINPUT107), .Z(new_n638_));
  NAND2_X1  g437(.A1(new_n545_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(G29gat), .B1(new_n640_), .B2(new_n525_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n636_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT43), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n544_), .A2(new_n499_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n643_), .B1(new_n644_), .B2(new_n572_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n572_), .ZN(new_n646_));
  AOI211_X1 g445(.A(KEYINPUT43), .B(new_n646_), .C1(new_n544_), .C2(new_n499_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n642_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  OAI211_X1 g449(.A(KEYINPUT44), .B(new_n642_), .C1(new_n645_), .C2(new_n647_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n525_), .A2(G29gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n641_), .B1(new_n652_), .B2(new_n653_), .ZN(G1328gat));
  NOR2_X1   g453(.A1(new_n401_), .A2(G36gat), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n545_), .A2(new_n638_), .A3(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n650_), .A2(new_n402_), .A3(new_n651_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n659_), .B2(G36gat), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT109), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT46), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n660_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n661_), .A2(new_n662_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n660_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n663_), .A2(new_n666_), .ZN(G1329gat));
  NAND4_X1  g466(.A1(new_n650_), .A2(G43gat), .A3(new_n348_), .A4(new_n651_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n639_), .A2(new_n500_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(G43gat), .B2(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g470(.A1(new_n652_), .A2(new_n468_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(G50gat), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n629_), .A2(G50gat), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT110), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n673_), .B1(new_n639_), .B2(new_n675_), .ZN(G1331gat));
  INV_X1    g475(.A(new_n268_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n301_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n679_), .A2(new_n300_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n680_), .A2(new_n644_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n681_), .A2(new_n589_), .ZN(new_n682_));
  INV_X1    g481(.A(G57gat), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(new_n683_), .A3(new_n525_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n680_), .A2(new_n636_), .A3(new_n610_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n685_), .A2(new_n525_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n684_), .B1(new_n683_), .B2(new_n686_), .ZN(G1332gat));
  NOR2_X1   g486(.A1(new_n401_), .A2(G64gat), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT111), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n682_), .A2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n685_), .A2(new_n402_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(G64gat), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n692_), .A2(KEYINPUT48), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(KEYINPUT48), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n690_), .B1(new_n693_), .B2(new_n694_), .ZN(G1333gat));
  INV_X1    g494(.A(G71gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n682_), .A2(new_n696_), .A3(new_n348_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n685_), .A2(new_n348_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(G71gat), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n699_), .A2(KEYINPUT49), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(KEYINPUT49), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n697_), .B1(new_n700_), .B2(new_n701_), .ZN(G1334gat));
  INV_X1    g501(.A(G78gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n682_), .A2(new_n703_), .A3(new_n468_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n685_), .A2(new_n468_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(G78gat), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n706_), .A2(KEYINPUT50), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(KEYINPUT50), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n704_), .B1(new_n707_), .B2(new_n708_), .ZN(G1335gat));
  AND2_X1   g508(.A1(new_n681_), .A2(new_n638_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n710_), .A2(new_n219_), .A3(new_n525_), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n645_), .A2(new_n647_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n679_), .A2(new_n636_), .A3(new_n300_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n525_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n711_), .B1(new_n716_), .B2(new_n219_), .ZN(G1336gat));
  NAND3_X1  g516(.A1(new_n710_), .A2(new_n220_), .A3(new_n402_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n714_), .A2(new_n402_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n718_), .B1(new_n720_), .B2(new_n220_), .ZN(G1337gat));
  INV_X1    g520(.A(KEYINPUT112), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n713_), .B(new_n348_), .C1(new_n645_), .C2(new_n647_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n722_), .B1(new_n724_), .B2(new_n324_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n723_), .A2(KEYINPUT112), .A3(G99gat), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n681_), .A2(new_n209_), .A3(new_n348_), .A4(new_n638_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n725_), .A2(new_n726_), .A3(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT113), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT51), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n729_), .A2(KEYINPUT51), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n728_), .A2(new_n730_), .A3(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n730_), .B1(new_n728_), .B2(new_n731_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1338gat));
  NAND3_X1  g533(.A1(new_n710_), .A2(new_n210_), .A3(new_n468_), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n713_), .B(new_n468_), .C1(new_n645_), .C2(new_n647_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT52), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n736_), .A2(new_n737_), .A3(G106gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n736_), .B2(G106gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g540(.A(KEYINPUT119), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n281_), .A2(new_n283_), .A3(new_n290_), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n743_), .B(new_n296_), .C1(new_n286_), .C2(new_n290_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n299_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT118), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n299_), .A2(new_n744_), .A3(KEYINPUT118), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(new_n258_), .ZN(new_n750_));
  XOR2_X1   g549(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n751_));
  NAND2_X1  g550(.A1(new_n249_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT116), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n234_), .A2(new_n246_), .A3(new_n244_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(new_n239_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT116), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n249_), .A2(new_n756_), .A3(new_n751_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n753_), .A2(new_n755_), .A3(new_n757_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n244_), .A2(new_n248_), .A3(KEYINPUT55), .A4(new_n246_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT117), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n255_), .B1(new_n758_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT56), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  OAI211_X1 g562(.A(KEYINPUT56), .B(new_n255_), .C1(new_n758_), .C2(new_n760_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n750_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n572_), .B(new_n742_), .C1(new_n765_), .C2(KEYINPUT58), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(KEYINPUT58), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT58), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n763_), .A2(new_n764_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(new_n770_), .B2(new_n750_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n742_), .B1(new_n771_), .B2(new_n572_), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT120), .B1(new_n768_), .B2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n572_), .B1(new_n765_), .B2(KEYINPUT58), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT119), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT120), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n767_), .A4(new_n766_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n300_), .A2(new_n258_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n778_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n749_), .A2(new_n259_), .A3(new_n261_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n608_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT57), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n773_), .A2(new_n777_), .A3(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n588_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n266_), .A2(new_n300_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n589_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n787_), .B2(KEYINPUT54), .ZN(new_n788_));
  XNOR2_X1  g587(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n785_), .B2(new_n589_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n788_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n784_), .A2(new_n792_), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n348_), .A2(new_n469_), .A3(new_n525_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT59), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n775_), .A2(new_n767_), .A3(new_n766_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n636_), .B1(new_n797_), .B2(new_n782_), .ZN(new_n798_));
  OR2_X1    g597(.A1(new_n798_), .A2(new_n791_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n794_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n800_), .A2(KEYINPUT121), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n800_), .A2(KEYINPUT121), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n801_), .A2(new_n802_), .A3(KEYINPUT59), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n799_), .A2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n796_), .A2(new_n300_), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(G113gat), .ZN(new_n806_));
  INV_X1    g605(.A(new_n300_), .ZN(new_n807_));
  OR3_X1    g606(.A1(new_n795_), .A2(G113gat), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(G1340gat));
  INV_X1    g608(.A(new_n679_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n796_), .A2(new_n810_), .A3(new_n804_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(G120gat), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n800_), .B1(new_n784_), .B2(new_n792_), .ZN(new_n813_));
  INV_X1    g612(.A(G120gat), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n679_), .B2(KEYINPUT60), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n813_), .B(new_n815_), .C1(KEYINPUT60), .C2(new_n814_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n812_), .A2(new_n816_), .ZN(G1341gat));
  NAND2_X1  g616(.A1(new_n636_), .A2(G127gat), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(KEYINPUT122), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT59), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n804_), .B(new_n819_), .C1(new_n813_), .C2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n781_), .B(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n823_), .B1(new_n797_), .B2(KEYINPUT120), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n636_), .B1(new_n824_), .B2(new_n777_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n636_), .B(new_n794_), .C1(new_n825_), .C2(new_n791_), .ZN(new_n826_));
  INV_X1    g625(.A(G127gat), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n821_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT123), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT123), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n821_), .A2(new_n831_), .A3(new_n828_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1342gat));
  AOI21_X1  g632(.A(G134gat), .B1(new_n813_), .B2(new_n609_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n796_), .A2(new_n804_), .ZN(new_n835_));
  XOR2_X1   g634(.A(KEYINPUT124), .B(G134gat), .Z(new_n836_));
  NOR2_X1   g635(.A1(new_n646_), .A2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n834_), .B1(new_n835_), .B2(new_n837_), .ZN(G1343gat));
  AOI21_X1  g637(.A(new_n791_), .B1(new_n783_), .B2(new_n588_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n348_), .A2(new_n498_), .A3(new_n539_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n839_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n300_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n810_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g645(.A1(new_n793_), .A2(new_n636_), .A3(new_n840_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT125), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT125), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n842_), .A2(new_n849_), .A3(new_n636_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(KEYINPUT61), .B(G155gat), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n848_), .A2(new_n850_), .A3(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n851_), .B1(new_n848_), .B2(new_n850_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n852_), .A2(new_n853_), .ZN(G1346gat));
  INV_X1    g653(.A(new_n842_), .ZN(new_n855_));
  OAI21_X1  g654(.A(G162gat), .B1(new_n855_), .B2(new_n646_), .ZN(new_n856_));
  INV_X1    g655(.A(G162gat), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n842_), .A2(new_n857_), .A3(new_n609_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(G1347gat));
  NAND3_X1  g658(.A1(new_n348_), .A2(new_n402_), .A3(new_n498_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(new_n468_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n799_), .A2(new_n300_), .A3(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT62), .B1(new_n862_), .B2(KEYINPUT22), .ZN(new_n863_));
  OAI21_X1  g662(.A(G169gat), .B1(new_n862_), .B2(KEYINPUT62), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(G169gat), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(new_n863_), .ZN(G1348gat));
  NAND3_X1  g666(.A1(new_n799_), .A2(new_n810_), .A3(new_n861_), .ZN(new_n868_));
  INV_X1    g667(.A(G176gat), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n839_), .A2(new_n468_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n679_), .A2(new_n869_), .A3(new_n860_), .ZN(new_n871_));
  AOI22_X1  g670(.A1(new_n868_), .A2(new_n869_), .B1(new_n870_), .B2(new_n871_), .ZN(G1349gat));
  NOR2_X1   g671(.A1(new_n860_), .A2(new_n588_), .ZN(new_n873_));
  AOI21_X1  g672(.A(G183gat), .B1(new_n870_), .B2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n799_), .A2(new_n861_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n875_), .A2(new_n588_), .A3(new_n303_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n874_), .A2(new_n876_), .ZN(G1350gat));
  OAI21_X1  g676(.A(G190gat), .B1(new_n875_), .B2(new_n646_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n609_), .A2(new_n304_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n875_), .B2(new_n879_), .ZN(G1351gat));
  NOR3_X1   g679(.A1(new_n348_), .A2(new_n629_), .A3(new_n525_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n881_), .A2(KEYINPUT126), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n881_), .A2(KEYINPUT126), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n882_), .A2(new_n883_), .A3(new_n401_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n793_), .A2(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n807_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(new_n360_), .ZN(G1352gat));
  INV_X1    g686(.A(KEYINPUT127), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n885_), .A2(new_n679_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(new_n352_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n889_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n891_));
  OAI211_X1 g690(.A(KEYINPUT127), .B(G204gat), .C1(new_n885_), .C2(new_n679_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n890_), .A2(new_n891_), .A3(new_n892_), .ZN(G1353gat));
  AND2_X1   g692(.A1(new_n793_), .A2(new_n884_), .ZN(new_n894_));
  AOI211_X1 g693(.A(KEYINPUT63), .B(G211gat), .C1(new_n894_), .C2(new_n636_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT63), .B(G211gat), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n885_), .A2(new_n588_), .A3(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n895_), .A2(new_n897_), .ZN(G1354gat));
  INV_X1    g697(.A(G218gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n894_), .A2(new_n899_), .A3(new_n609_), .ZN(new_n900_));
  OAI21_X1  g699(.A(G218gat), .B1(new_n885_), .B2(new_n646_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(G1355gat));
endmodule


