//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 0 1 1 1 1 0 1 0 0 1 1 1 1 1 0 1 0 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 1 0 0 1 1 1 0 0 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n927_, new_n928_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n940_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n954_;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G85gat), .B(G92gat), .ZN(new_n203_));
  AOI21_X1  g002(.A(new_n203_), .B1(KEYINPUT64), .B2(KEYINPUT8), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT6), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT7), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n204_), .B1(new_n207_), .B2(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(KEYINPUT64), .A2(KEYINPUT8), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT9), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n203_), .A2(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(KEYINPUT10), .B(G99gat), .Z(new_n216_));
  INV_X1    g015(.A(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n214_), .A2(G85gat), .A3(G92gat), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n215_), .A2(new_n218_), .A3(new_n219_), .A4(new_n206_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n213_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT65), .ZN(new_n222_));
  INV_X1    g021(.A(new_n220_), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n211_), .A2(new_n212_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n211_), .A2(new_n212_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n223_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT65), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n222_), .A2(new_n228_), .ZN(new_n229_));
  XOR2_X1   g028(.A(G29gat), .B(G36gat), .Z(new_n230_));
  XOR2_X1   g029(.A(G43gat), .B(G50gat), .Z(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n202_), .B1(new_n229_), .B2(new_n233_), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n222_), .A2(KEYINPUT71), .A3(new_n228_), .A4(new_n232_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n232_), .B(KEYINPUT15), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT35), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G232gat), .A2(G233gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT34), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  AOI22_X1  g040(.A1(new_n221_), .A2(new_n237_), .B1(new_n238_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n236_), .A2(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n241_), .A2(new_n238_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G190gat), .B(G218gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G134gat), .B(G162gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n248_), .A2(KEYINPUT36), .ZN(new_n249_));
  INV_X1    g048(.A(new_n244_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n236_), .A2(new_n250_), .A3(new_n242_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n245_), .A2(new_n249_), .A3(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n248_), .B(KEYINPUT36), .Z(new_n253_));
  AOI21_X1  g052(.A(new_n250_), .B1(new_n236_), .B2(new_n242_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n242_), .ZN(new_n255_));
  AOI211_X1 g054(.A(new_n244_), .B(new_n255_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n253_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT37), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n252_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n258_), .B1(new_n252_), .B2(new_n257_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G15gat), .B(G22gat), .ZN(new_n262_));
  INV_X1    g061(.A(G1gat), .ZN(new_n263_));
  INV_X1    g062(.A(G8gat), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT14), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G1gat), .B(G8gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G231gat), .A2(G233gat), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n269_), .B(KEYINPUT72), .Z(new_n270_));
  XNOR2_X1  g069(.A(new_n268_), .B(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G57gat), .B(G64gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT11), .ZN(new_n273_));
  OR2_X1    g072(.A1(new_n273_), .A2(KEYINPUT66), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(KEYINPUT66), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n272_), .A2(KEYINPUT11), .ZN(new_n277_));
  XOR2_X1   g076(.A(G71gat), .B(G78gat), .Z(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n276_), .A2(new_n279_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n274_), .A2(new_n277_), .A3(new_n278_), .A4(new_n275_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n271_), .B(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G183gat), .B(G211gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT74), .ZN(new_n285_));
  XOR2_X1   g084(.A(G127gat), .B(G155gat), .Z(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n283_), .A2(KEYINPUT17), .A3(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT75), .ZN(new_n291_));
  XOR2_X1   g090(.A(new_n289_), .B(KEYINPUT17), .Z(new_n292_));
  AND3_X1   g091(.A1(new_n280_), .A2(KEYINPUT67), .A3(new_n281_), .ZN(new_n293_));
  AOI21_X1  g092(.A(KEYINPUT67), .B1(new_n280_), .B2(new_n281_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(new_n271_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n292_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n291_), .A2(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n261_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G230gat), .A2(G233gat), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT68), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n226_), .A2(new_n227_), .ZN(new_n303_));
  AOI211_X1 g102(.A(KEYINPUT65), .B(new_n223_), .C1(new_n224_), .C2(new_n225_), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n295_), .B(new_n302_), .C1(new_n303_), .C2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT67), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n282_), .A2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n280_), .A2(KEYINPUT67), .A3(new_n281_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n222_), .A2(new_n309_), .A3(new_n228_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n305_), .A2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n302_), .B1(new_n229_), .B2(new_n295_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n301_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n303_), .A2(new_n304_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT69), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n280_), .A2(KEYINPUT12), .A3(new_n281_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n315_), .B1(new_n226_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n316_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(new_n221_), .A3(KEYINPUT69), .ZN(new_n319_));
  AOI22_X1  g118(.A1(new_n314_), .A2(new_n309_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT12), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n321_), .B1(new_n314_), .B2(new_n309_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(new_n322_), .A3(new_n300_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G120gat), .B(G148gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT5), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G176gat), .B(G204gat), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n325_), .B(new_n326_), .Z(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n313_), .A2(new_n323_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n327_), .B(KEYINPUT70), .Z(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n332_), .B1(new_n313_), .B2(new_n323_), .ZN(new_n333_));
  OR3_X1    g132(.A1(new_n330_), .A2(KEYINPUT13), .A3(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT13), .B1(new_n330_), .B2(new_n333_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n299_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT76), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G227gat), .A2(G233gat), .ZN(new_n339_));
  INV_X1    g138(.A(G71gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT25), .B(G183gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT80), .B(G190gat), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT26), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n343_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G183gat), .A2(G190gat), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n349_), .A2(KEYINPUT81), .A3(KEYINPUT23), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(KEYINPUT23), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT81), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n349_), .B(KEYINPUT82), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n350_), .B(new_n353_), .C1(new_n354_), .C2(KEYINPUT23), .ZN(new_n355_));
  NOR3_X1   g154(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT24), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n357_), .B1(G169gat), .B2(G176gat), .ZN(new_n358_));
  INV_X1    g157(.A(G169gat), .ZN(new_n359_));
  INV_X1    g158(.A(G176gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n356_), .B1(new_n358_), .B2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n348_), .A2(new_n355_), .A3(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT83), .B(G169gat), .ZN(new_n364_));
  NOR2_X1   g163(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT23), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n349_), .A2(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n368_), .B1(new_n354_), .B2(new_n367_), .ZN(new_n369_));
  INV_X1    g168(.A(G183gat), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n344_), .A2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n366_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n372_));
  AND3_X1   g171(.A1(new_n363_), .A2(new_n372_), .A3(KEYINPUT30), .ZN(new_n373_));
  AOI21_X1  g172(.A(KEYINPUT30), .B1(new_n363_), .B2(new_n372_), .ZN(new_n374_));
  OAI21_X1  g173(.A(G99gat), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n363_), .A2(new_n372_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT30), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(G99gat), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n363_), .A2(new_n372_), .A3(KEYINPUT30), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n378_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G15gat), .B(G43gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT84), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n375_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n383_), .B1(new_n375_), .B2(new_n381_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n342_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n375_), .A2(new_n381_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n383_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n375_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(new_n341_), .A3(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT85), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n386_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT31), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT31), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n386_), .A2(new_n391_), .A3(new_n392_), .A4(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G127gat), .B(G134gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G113gat), .B(G120gat), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n398_), .B(new_n399_), .Z(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n397_), .A2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n394_), .A2(new_n400_), .A3(new_n396_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(G197gat), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n405_), .A2(G204gat), .ZN(new_n406_));
  INV_X1    g205(.A(G204gat), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n407_), .A2(G197gat), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT21), .B1(new_n406_), .B2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G211gat), .B(G218gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n408_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT90), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n405_), .B2(G204gat), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n407_), .A2(KEYINPUT90), .A3(G197gat), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n411_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n409_), .B(new_n410_), .C1(new_n415_), .C2(KEYINPUT21), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT91), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n411_), .A2(KEYINPUT91), .A3(new_n413_), .A4(new_n414_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT21), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n410_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n418_), .A2(new_n419_), .A3(new_n421_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n363_), .A2(new_n372_), .A3(new_n416_), .A4(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT26), .B(G190gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n343_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n362_), .A2(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n369_), .A2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n359_), .A2(new_n360_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT22), .B(G169gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT92), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n428_), .B1(new_n430_), .B2(new_n360_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n355_), .B1(G183gat), .B2(G190gat), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n427_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n422_), .A2(new_n416_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  OAI211_X1 g234(.A(KEYINPUT20), .B(new_n423_), .C1(new_n433_), .C2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G226gat), .A2(G233gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT19), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G8gat), .B(G36gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT18), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G64gat), .B(G92gat), .ZN(new_n442_));
  XOR2_X1   g241(.A(new_n441_), .B(new_n442_), .Z(new_n443_));
  NAND2_X1  g242(.A1(new_n433_), .A2(new_n435_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n376_), .A2(new_n434_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n438_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n444_), .A2(new_n445_), .A3(KEYINPUT20), .A4(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n439_), .A2(new_n443_), .A3(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n436_), .A2(new_n438_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n444_), .A2(KEYINPUT20), .A3(new_n445_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n449_), .B1(new_n438_), .B2(new_n450_), .ZN(new_n451_));
  OAI211_X1 g250(.A(KEYINPUT27), .B(new_n448_), .C1(new_n451_), .C2(new_n443_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT27), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n439_), .A2(new_n443_), .A3(new_n447_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n443_), .B1(new_n439_), .B2(new_n447_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n453_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n452_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(G141gat), .ZN(new_n459_));
  INV_X1    g258(.A(G148gat), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(G141gat), .A2(G148gat), .ZN(new_n462_));
  AND2_X1   g261(.A1(G155gat), .A2(G162gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT1), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT86), .ZN(new_n465_));
  INV_X1    g264(.A(G155gat), .ZN(new_n466_));
  INV_X1    g265(.A(G162gat), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT86), .B1(G155gat), .B2(G162gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  AOI211_X1 g269(.A(new_n461_), .B(new_n462_), .C1(new_n464_), .C2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n463_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n469_), .ZN(new_n474_));
  NOR3_X1   g273(.A1(KEYINPUT86), .A2(G155gat), .A3(G162gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n473_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT87), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT87), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n470_), .A2(new_n478_), .A3(new_n473_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT2), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n481_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT3), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n462_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n482_), .A2(new_n484_), .A3(new_n485_), .A4(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT88), .B1(new_n480_), .B2(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n478_), .B1(new_n470_), .B2(new_n473_), .ZN(new_n489_));
  AOI211_X1 g288(.A(KEYINPUT87), .B(new_n463_), .C1(new_n468_), .C2(new_n469_), .ZN(new_n490_));
  OAI211_X1 g289(.A(KEYINPUT88), .B(new_n487_), .C1(new_n489_), .C2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n472_), .B1(new_n488_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT89), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n487_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT88), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n471_), .B1(new_n498_), .B2(new_n491_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT89), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n495_), .A2(new_n500_), .A3(new_n400_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n493_), .A2(new_n400_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G225gat), .A2(G233gat), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n501_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  AND3_X1   g304(.A1(new_n501_), .A2(KEYINPUT4), .A3(new_n503_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT4), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n495_), .A2(new_n500_), .A3(new_n507_), .A4(new_n400_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n504_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n505_), .B1(new_n506_), .B2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G1gat), .B(G29gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(G85gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(KEYINPUT0), .B(G57gat), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n513_), .B(new_n514_), .Z(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n498_), .A2(new_n491_), .ZN(new_n517_));
  AOI21_X1  g316(.A(KEYINPUT89), .B1(new_n517_), .B2(new_n472_), .ZN(new_n518_));
  AOI211_X1 g317(.A(new_n494_), .B(new_n471_), .C1(new_n498_), .C2(new_n491_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n502_), .B1(new_n520_), .B2(new_n400_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n516_), .B1(new_n521_), .B2(new_n504_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n501_), .A2(KEYINPUT4), .A3(new_n503_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n523_), .A2(new_n509_), .A3(new_n508_), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n511_), .A2(new_n516_), .B1(new_n522_), .B2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G22gat), .B(G50gat), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT28), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n495_), .A2(new_n500_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT29), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n527_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  AOI211_X1 g329(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n495_), .C2(new_n500_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n526_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  XOR2_X1   g331(.A(G78gat), .B(G106gat), .Z(new_n533_));
  INV_X1    g332(.A(G228gat), .ZN(new_n534_));
  INV_X1    g333(.A(G233gat), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n434_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n536_), .B1(new_n520_), .B2(KEYINPUT29), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n434_), .B1(new_n499_), .B2(new_n529_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n534_), .A2(new_n535_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n533_), .B1(new_n537_), .B2(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT28), .B1(new_n520_), .B2(KEYINPUT29), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n528_), .A2(new_n527_), .A3(new_n529_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n526_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n495_), .A2(KEYINPUT29), .A3(new_n500_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n536_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n533_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(new_n550_), .A3(new_n540_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n532_), .A2(new_n542_), .A3(new_n546_), .A4(new_n551_), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n543_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n545_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n554_));
  AOI221_X4 g353(.A(new_n533_), .B1(new_n539_), .B2(new_n538_), .C1(new_n547_), .C2(new_n548_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n550_), .B1(new_n549_), .B2(new_n540_), .ZN(new_n556_));
  OAI22_X1  g355(.A1(new_n553_), .A2(new_n554_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n458_), .A2(new_n525_), .A3(new_n552_), .A4(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n404_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n552_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n560_), .A2(new_n525_), .A3(new_n458_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n443_), .A2(KEYINPUT32), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n439_), .A2(new_n447_), .A3(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n563_), .B1(new_n451_), .B2(new_n562_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n511_), .A2(new_n516_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n522_), .A2(new_n524_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n564_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n508_), .A2(new_n504_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n515_), .B1(new_n568_), .B2(new_n523_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT96), .ZN(new_n570_));
  NOR3_X1   g369(.A1(new_n518_), .A2(new_n519_), .A3(new_n401_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n570_), .B1(new_n571_), .B2(new_n502_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n501_), .A2(KEYINPUT96), .A3(new_n503_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n572_), .A2(new_n509_), .A3(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n569_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT93), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n576_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n439_), .A2(new_n447_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n443_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n580_), .A2(KEYINPUT93), .A3(new_n448_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n577_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n522_), .A2(KEYINPUT33), .A3(new_n524_), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n575_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n566_), .A2(KEYINPUT94), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT94), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n522_), .A2(new_n586_), .A3(new_n524_), .ZN(new_n587_));
  XOR2_X1   g386(.A(KEYINPUT95), .B(KEYINPUT33), .Z(new_n588_));
  NAND3_X1  g387(.A1(new_n585_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n567_), .B1(new_n584_), .B2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n561_), .B1(new_n590_), .B2(new_n560_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n559_), .B1(new_n591_), .B2(new_n404_), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n266_), .B(new_n267_), .Z(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(new_n232_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n233_), .A2(new_n268_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT77), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G229gat), .A2(G233gat), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n594_), .A2(new_n595_), .A3(KEYINPUT77), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n598_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n237_), .A2(new_n268_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(new_n599_), .A3(new_n594_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G113gat), .B(G141gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G169gat), .B(G197gat), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n606_), .B(new_n607_), .Z(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(KEYINPUT79), .B1(new_n605_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT79), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n602_), .A2(new_n604_), .A3(new_n611_), .A4(new_n608_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n608_), .B(KEYINPUT78), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n605_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n592_), .A2(new_n617_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n338_), .A2(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n525_), .A2(G1gat), .ZN(new_n620_));
  AOI22_X1  g419(.A1(new_n619_), .A2(new_n620_), .B1(KEYINPUT98), .B2(KEYINPUT38), .ZN(new_n621_));
  NOR2_X1   g420(.A1(KEYINPUT98), .A2(KEYINPUT38), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n253_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n624_), .B1(new_n245_), .B2(new_n251_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n249_), .ZN(new_n626_));
  NOR3_X1   g425(.A1(new_n254_), .A2(new_n256_), .A3(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n336_), .A2(new_n616_), .ZN(new_n629_));
  NOR4_X1   g428(.A1(new_n592_), .A2(new_n628_), .A3(new_n629_), .A4(new_n298_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n565_), .A2(new_n566_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n263_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n632_), .B(KEYINPUT97), .Z(new_n633_));
  NAND2_X1  g432(.A1(new_n621_), .A2(new_n622_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n623_), .A2(new_n633_), .A3(new_n634_), .ZN(G1324gat));
  NAND3_X1  g434(.A1(new_n619_), .A2(new_n264_), .A3(new_n457_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n630_), .A2(new_n457_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(KEYINPUT99), .B(KEYINPUT39), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n637_), .A2(G8gat), .A3(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n637_), .B2(G8gat), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n636_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g441(.A(G15gat), .ZN(new_n643_));
  INV_X1    g442(.A(new_n404_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n619_), .A2(new_n643_), .A3(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n643_), .B1(new_n630_), .B2(new_n644_), .ZN(new_n646_));
  XOR2_X1   g445(.A(KEYINPUT100), .B(KEYINPUT41), .Z(new_n647_));
  OR2_X1    g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n647_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n645_), .A2(new_n648_), .A3(new_n649_), .ZN(G1326gat));
  INV_X1    g449(.A(G22gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n630_), .B2(new_n560_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT42), .Z(new_n653_));
  NAND3_X1  g452(.A1(new_n619_), .A2(new_n651_), .A3(new_n560_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1327gat));
  INV_X1    g454(.A(new_n628_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n298_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n658_), .A2(new_n336_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n618_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(G29gat), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n631_), .A2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT102), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n660_), .A2(new_n663_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n629_), .A2(new_n657_), .ZN(new_n665_));
  OAI21_X1  g464(.A(KEYINPUT37), .B1(new_n625_), .B2(new_n627_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n252_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n592_), .A2(KEYINPUT43), .A3(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT43), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n404_), .A2(new_n558_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n560_), .A2(new_n525_), .A3(new_n458_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n564_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n631_), .A2(new_n673_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n522_), .A2(new_n586_), .A3(new_n524_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n586_), .B1(new_n522_), .B2(new_n524_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n588_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n675_), .A2(new_n676_), .A3(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n575_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n674_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n560_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n672_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n671_), .B1(new_n682_), .B2(new_n644_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n670_), .B1(new_n683_), .B2(new_n261_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n665_), .B1(new_n669_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n685_), .A2(new_n686_), .A3(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n665_), .ZN(new_n689_));
  OAI21_X1  g488(.A(KEYINPUT43), .B1(new_n592_), .B2(new_n668_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n680_), .A2(new_n681_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n644_), .B1(new_n691_), .B2(new_n561_), .ZN(new_n692_));
  OAI211_X1 g491(.A(new_n670_), .B(new_n261_), .C1(new_n692_), .C2(new_n559_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n689_), .B1(new_n690_), .B2(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(KEYINPUT101), .B1(new_n694_), .B2(KEYINPUT44), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n688_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(KEYINPUT44), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n696_), .A2(new_n631_), .A3(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n664_), .B1(new_n698_), .B2(new_n661_), .ZN(G1328gat));
  AOI21_X1  g498(.A(new_n458_), .B1(new_n694_), .B2(KEYINPUT44), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n686_), .B1(new_n685_), .B2(new_n687_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n694_), .A2(KEYINPUT101), .A3(KEYINPUT44), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n700_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(G36gat), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT46), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n458_), .A2(G36gat), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n618_), .A2(new_n659_), .A3(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT103), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT103), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n618_), .A2(new_n709_), .A3(new_n659_), .A4(new_n706_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT45), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n708_), .A2(new_n710_), .A3(KEYINPUT45), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n704_), .A2(KEYINPUT104), .A3(new_n705_), .A4(new_n715_), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n705_), .A2(KEYINPUT104), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n705_), .A2(KEYINPUT104), .ZN(new_n718_));
  INV_X1    g517(.A(G36gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n719_), .B1(new_n696_), .B2(new_n700_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n713_), .A2(new_n714_), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n717_), .B(new_n718_), .C1(new_n720_), .C2(new_n721_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n716_), .A2(new_n722_), .ZN(G1329gat));
  NAND4_X1  g522(.A1(new_n696_), .A2(G43gat), .A3(new_n644_), .A4(new_n697_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n660_), .A2(new_n644_), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n725_), .A2(G43gat), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT47), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n724_), .A2(new_n729_), .A3(new_n726_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1330gat));
  INV_X1    g530(.A(KEYINPUT105), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n560_), .B(new_n697_), .C1(new_n701_), .C2(new_n702_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(G50gat), .ZN(new_n734_));
  INV_X1    g533(.A(G50gat), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n660_), .A2(new_n735_), .A3(new_n560_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n732_), .B1(new_n734_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n736_), .ZN(new_n738_));
  AOI211_X1 g537(.A(KEYINPUT105), .B(new_n738_), .C1(new_n733_), .C2(G50gat), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n737_), .A2(new_n739_), .ZN(G1331gat));
  NOR2_X1   g539(.A1(new_n336_), .A2(new_n616_), .ZN(new_n741_));
  AND4_X1   g540(.A1(new_n683_), .A2(new_n656_), .A3(new_n657_), .A4(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n742_), .A2(G57gat), .A3(new_n631_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT106), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n592_), .A2(new_n616_), .A3(new_n336_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n745_), .A2(new_n299_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(new_n631_), .ZN(new_n747_));
  INV_X1    g546(.A(G57gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  AOI211_X1 g548(.A(KEYINPUT106), .B(G57gat), .C1(new_n746_), .C2(new_n631_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n743_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT107), .ZN(G1332gat));
  INV_X1    g551(.A(G64gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n746_), .A2(new_n753_), .A3(new_n457_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n742_), .A2(new_n457_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(G64gat), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n756_), .A2(KEYINPUT48), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n756_), .A2(KEYINPUT48), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT108), .ZN(G1333gat));
  AOI21_X1  g559(.A(new_n340_), .B1(new_n742_), .B2(new_n644_), .ZN(new_n761_));
  XOR2_X1   g560(.A(new_n761_), .B(KEYINPUT49), .Z(new_n762_));
  NAND3_X1  g561(.A1(new_n746_), .A2(new_n340_), .A3(new_n644_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1334gat));
  INV_X1    g563(.A(G78gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n742_), .B2(new_n560_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n766_), .B(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n560_), .A2(new_n765_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT110), .Z(new_n770_));
  NAND2_X1  g569(.A1(new_n746_), .A2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n768_), .A2(new_n771_), .ZN(G1335gat));
  INV_X1    g571(.A(G85gat), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n745_), .A2(new_n658_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n774_), .B2(new_n525_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT111), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n690_), .A2(new_n693_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n777_), .A2(new_n298_), .A3(new_n741_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n778_), .A2(new_n773_), .A3(new_n525_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n776_), .A2(new_n779_), .ZN(G1336gat));
  OAI21_X1  g579(.A(G92gat), .B1(new_n778_), .B2(new_n458_), .ZN(new_n781_));
  OR3_X1    g580(.A1(new_n774_), .A2(G92gat), .A3(new_n458_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(G1337gat));
  INV_X1    g582(.A(new_n774_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n784_), .A2(new_n644_), .A3(new_n216_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n777_), .A2(new_n644_), .A3(new_n298_), .A4(new_n741_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n786_), .A2(new_n787_), .A3(G99gat), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n786_), .B2(G99gat), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n785_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n791_), .A2(KEYINPUT113), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n790_), .B(new_n792_), .ZN(G1338gat));
  NAND3_X1  g592(.A1(new_n784_), .A2(new_n217_), .A3(new_n560_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n777_), .A2(new_n560_), .A3(new_n298_), .A4(new_n741_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n795_), .A2(new_n796_), .A3(G106gat), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n795_), .B2(G106gat), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n794_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g599(.A1(new_n329_), .A2(new_n616_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT115), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n329_), .A2(new_n803_), .A3(new_n616_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n300_), .B1(new_n320_), .B2(new_n322_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n323_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n320_), .A2(new_n322_), .A3(KEYINPUT55), .A4(new_n300_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n331_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT56), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n810_), .A2(KEYINPUT56), .A3(new_n331_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n805_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n330_), .A2(new_n333_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n603_), .A2(new_n600_), .A3(new_n594_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n598_), .A2(new_n599_), .A3(new_n601_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n609_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n819_), .A2(KEYINPUT116), .A3(new_n609_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n818_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  OR2_X1    g623(.A1(new_n824_), .A2(KEYINPUT117), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(KEYINPUT117), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n613_), .A3(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n816_), .A2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n656_), .B1(new_n815_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n827_), .A2(new_n330_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT56), .B1(new_n810_), .B2(new_n331_), .ZN(new_n832_));
  AOI211_X1 g631(.A(new_n812_), .B(new_n332_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n831_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT58), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n668_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n831_), .B(KEYINPUT58), .C1(new_n832_), .C2(new_n833_), .ZN(new_n837_));
  AOI22_X1  g636(.A1(new_n829_), .A2(new_n830_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  OAI211_X1 g637(.A(KEYINPUT57), .B(new_n656_), .C1(new_n815_), .C2(new_n828_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n298_), .ZN(new_n841_));
  XOR2_X1   g640(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n843_), .B1(new_n337_), .B2(new_n616_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n299_), .A2(new_n617_), .A3(new_n336_), .A4(new_n842_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n560_), .B1(new_n841_), .B2(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n525_), .A2(new_n457_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n644_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n847_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(G113gat), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(new_n853_), .A3(new_n616_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n851_), .A2(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n847_), .A2(KEYINPUT59), .A3(new_n850_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n617_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n854_), .B1(new_n858_), .B2(new_n853_), .ZN(G1340gat));
  INV_X1    g658(.A(G120gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n336_), .B2(KEYINPUT60), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n852_), .B(new_n861_), .C1(KEYINPUT60), .C2(new_n860_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n336_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(new_n860_), .ZN(G1341gat));
  AOI21_X1  g663(.A(G127gat), .B1(new_n852_), .B2(new_n657_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n856_), .A2(new_n857_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n657_), .A2(G127gat), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(KEYINPUT118), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n865_), .B1(new_n866_), .B2(new_n868_), .ZN(G1342gat));
  AOI21_X1  g668(.A(G134gat), .B1(new_n852_), .B2(new_n628_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n261_), .A2(G134gat), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(KEYINPUT119), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n870_), .B1(new_n866_), .B2(new_n872_), .ZN(G1343gat));
  NOR3_X1   g672(.A1(new_n681_), .A2(new_n525_), .A3(new_n457_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n657_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n844_), .A2(new_n845_), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n404_), .B(new_n874_), .C1(new_n875_), .C2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n877_), .A2(new_n878_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n616_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(G141gat), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n644_), .B1(new_n841_), .B2(new_n846_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n884_), .A2(KEYINPUT120), .A3(new_n874_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n879_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n886_), .A2(new_n459_), .A3(new_n616_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n883_), .A2(new_n887_), .ZN(G1344gat));
  XNOR2_X1  g687(.A(KEYINPUT121), .B(G148gat), .ZN(new_n889_));
  INV_X1    g688(.A(new_n336_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n886_), .B2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n889_), .ZN(new_n892_));
  AOI211_X1 g691(.A(new_n336_), .B(new_n892_), .C1(new_n885_), .C2(new_n879_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n891_), .A2(new_n893_), .ZN(G1345gat));
  OAI21_X1  g693(.A(new_n657_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT61), .B(G155gat), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n896_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n886_), .A2(new_n657_), .A3(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n899_), .ZN(G1346gat));
  NAND3_X1  g699(.A1(new_n886_), .A2(new_n467_), .A3(new_n628_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n668_), .B1(new_n885_), .B2(new_n879_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n467_), .B2(new_n902_), .ZN(G1347gat));
  NAND2_X1  g702(.A1(new_n525_), .A2(new_n457_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n404_), .A2(new_n904_), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n847_), .A2(new_n430_), .A3(new_n616_), .A4(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n616_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(KEYINPUT122), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n681_), .B(new_n908_), .C1(new_n875_), .C2(new_n876_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT62), .ZN(new_n910_));
  AND3_X1   g709(.A1(new_n909_), .A2(new_n910_), .A3(G169gat), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n910_), .B1(new_n909_), .B2(G169gat), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n906_), .B1(new_n911_), .B2(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  OAI211_X1 g714(.A(KEYINPUT123), .B(new_n906_), .C1(new_n911_), .C2(new_n912_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1348gat));
  OAI211_X1 g716(.A(new_n681_), .B(new_n905_), .C1(new_n875_), .C2(new_n876_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n336_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(new_n360_), .ZN(G1349gat));
  OR3_X1    g719(.A1(new_n918_), .A2(new_n343_), .A3(new_n298_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n370_), .B1(new_n918_), .B2(new_n298_), .ZN(new_n923_));
  AND3_X1   g722(.A1(new_n921_), .A2(new_n922_), .A3(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n922_), .B1(new_n921_), .B2(new_n923_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n924_), .A2(new_n925_), .ZN(G1350gat));
  OAI21_X1  g725(.A(G190gat), .B1(new_n918_), .B2(new_n668_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n628_), .A2(new_n424_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n927_), .B1(new_n918_), .B2(new_n928_), .ZN(G1351gat));
  NOR2_X1   g728(.A1(new_n681_), .A2(new_n904_), .ZN(new_n930_));
  NAND4_X1  g729(.A1(new_n884_), .A2(G197gat), .A3(new_n616_), .A4(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n932_));
  AND2_X1   g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n841_), .A2(new_n846_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n934_), .A2(new_n404_), .A3(new_n930_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n935_), .ZN(new_n936_));
  AOI21_X1  g735(.A(G197gat), .B1(new_n936_), .B2(new_n616_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n931_), .A2(new_n932_), .ZN(new_n938_));
  NOR3_X1   g737(.A1(new_n933_), .A2(new_n937_), .A3(new_n938_), .ZN(G1352gat));
  NOR2_X1   g738(.A1(new_n935_), .A2(new_n336_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(new_n407_), .ZN(G1353gat));
  NOR2_X1   g740(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n942_), .B1(new_n935_), .B2(new_n298_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n943_), .A2(new_n944_), .ZN(new_n945_));
  OAI211_X1 g744(.A(KEYINPUT127), .B(new_n942_), .C1(new_n935_), .C2(new_n298_), .ZN(new_n946_));
  XOR2_X1   g745(.A(KEYINPUT63), .B(G211gat), .Z(new_n947_));
  NAND4_X1  g746(.A1(new_n936_), .A2(KEYINPUT126), .A3(new_n657_), .A4(new_n947_), .ZN(new_n948_));
  NAND4_X1  g747(.A1(new_n884_), .A2(new_n657_), .A3(new_n930_), .A4(new_n947_), .ZN(new_n949_));
  INV_X1    g748(.A(KEYINPUT126), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n949_), .A2(new_n950_), .ZN(new_n951_));
  AOI22_X1  g750(.A1(new_n945_), .A2(new_n946_), .B1(new_n948_), .B2(new_n951_), .ZN(G1354gat));
  OR3_X1    g751(.A1(new_n935_), .A2(G218gat), .A3(new_n656_), .ZN(new_n953_));
  OAI21_X1  g752(.A(G218gat), .B1(new_n935_), .B2(new_n668_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n953_), .A2(new_n954_), .ZN(G1355gat));
endmodule


