//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_, new_n934_;
  XOR2_X1   g000(.A(G57gat), .B(G64gat), .Z(new_n202_));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT68), .ZN(new_n205_));
  XOR2_X1   g004(.A(G71gat), .B(G78gat), .Z(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n205_), .B1(new_n204_), .B2(new_n206_), .ZN(new_n209_));
  OAI22_X1  g008(.A1(new_n208_), .A2(new_n209_), .B1(new_n203_), .B2(new_n202_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n209_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n202_), .A2(new_n203_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n211_), .A2(new_n212_), .A3(new_n207_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G15gat), .B(G22gat), .ZN(new_n215_));
  INV_X1    g014(.A(G1gat), .ZN(new_n216_));
  INV_X1    g015(.A(G8gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT14), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n215_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G1gat), .B(G8gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n219_), .B(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n214_), .B(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G231gat), .A2(G233gat), .ZN(new_n223_));
  XOR2_X1   g022(.A(new_n222_), .B(new_n223_), .Z(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n224_), .A2(new_n226_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT76), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(G183gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G127gat), .B(G155gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(G211gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n231_), .B(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT17), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n227_), .A2(new_n228_), .A3(new_n235_), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n227_), .A2(new_n228_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT17), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n234_), .A2(new_n238_), .ZN(new_n239_));
  OAI211_X1 g038(.A(KEYINPUT77), .B(new_n236_), .C1(new_n237_), .C2(new_n239_), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n236_), .A2(KEYINPUT77), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G99gat), .A2(G106gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT6), .ZN(new_n245_));
  XOR2_X1   g044(.A(new_n245_), .B(KEYINPUT64), .Z(new_n246_));
  NOR2_X1   g045(.A1(G99gat), .A2(G106gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n248_));
  XOR2_X1   g047(.A(new_n247_), .B(new_n248_), .Z(new_n249_));
  INV_X1    g048(.A(KEYINPUT8), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT9), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n252_), .A2(G85gat), .A3(G92gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G85gat), .B(G92gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT10), .B(G99gat), .ZN(new_n255_));
  OAI221_X1 g054(.A(new_n253_), .B1(new_n254_), .B2(new_n252_), .C1(G106gat), .C2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n251_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n246_), .A2(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n254_), .B(KEYINPUT66), .Z(new_n259_));
  INV_X1    g058(.A(KEYINPUT67), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n245_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n249_), .A2(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n245_), .A2(new_n260_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n259_), .B(KEYINPUT8), .C1(new_n262_), .C2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n254_), .B(KEYINPUT66), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(new_n250_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n258_), .A2(new_n264_), .A3(new_n266_), .ZN(new_n267_));
  XOR2_X1   g066(.A(G43gat), .B(G50gat), .Z(new_n268_));
  XNOR2_X1  g067(.A(G29gat), .B(G36gat), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n269_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT15), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT35), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G232gat), .A2(G233gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT34), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  AOI22_X1  g077(.A1(new_n267_), .A2(new_n274_), .B1(new_n275_), .B2(new_n278_), .ZN(new_n279_));
  AOI22_X1  g078(.A1(new_n246_), .A2(new_n257_), .B1(new_n250_), .B2(new_n265_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n280_), .A2(new_n270_), .A3(new_n271_), .A4(new_n264_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n278_), .A2(new_n275_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n283_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n279_), .A2(new_n285_), .A3(new_n281_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G190gat), .B(G218gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G134gat), .B(G162gat), .ZN(new_n288_));
  XOR2_X1   g087(.A(new_n287_), .B(new_n288_), .Z(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n290_), .A2(KEYINPUT36), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n284_), .A2(new_n286_), .A3(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n289_), .B(KEYINPUT36), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n294_), .B1(new_n284_), .B2(new_n286_), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT37), .B1(new_n292_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT71), .ZN(new_n297_));
  INV_X1    g096(.A(new_n286_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n285_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n293_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT72), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n295_), .A2(KEYINPUT72), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT37), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n284_), .A2(new_n286_), .A3(new_n291_), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n302_), .A2(new_n303_), .A3(new_n304_), .A4(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT71), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n307_), .B(KEYINPUT37), .C1(new_n292_), .C2(new_n295_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n297_), .A2(new_n306_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n243_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n267_), .A2(new_n213_), .A3(new_n210_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n214_), .A2(new_n264_), .A3(new_n280_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n312_), .A2(new_n313_), .A3(KEYINPUT12), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT12), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n267_), .A2(new_n315_), .A3(new_n213_), .A4(new_n210_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G230gat), .A2(G233gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n312_), .A2(new_n313_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n318_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(G176gat), .B(G204gat), .Z(new_n323_));
  XNOR2_X1  g122(.A(G120gat), .B(G148gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(KEYINPUT69), .B(KEYINPUT5), .Z(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n319_), .A2(new_n322_), .A3(new_n327_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n319_), .A2(new_n322_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n327_), .B(KEYINPUT70), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n328_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n331_), .B(KEYINPUT13), .Z(new_n332_));
  NAND2_X1  g131(.A1(new_n274_), .A2(new_n221_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G229gat), .A2(G233gat), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n221_), .A2(new_n272_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n333_), .A2(new_n334_), .A3(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n221_), .B(new_n272_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n338_), .A2(G229gat), .A3(G233gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(G169gat), .B(G197gat), .Z(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT78), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G113gat), .B(G141gat), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n342_), .B(new_n343_), .Z(new_n344_));
  OR2_X1    g143(.A1(new_n340_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n340_), .A2(new_n344_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n332_), .A2(new_n348_), .ZN(new_n349_));
  XOR2_X1   g148(.A(G155gat), .B(G162gat), .Z(new_n350_));
  INV_X1    g149(.A(G141gat), .ZN(new_n351_));
  INV_X1    g150(.A(G148gat), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(new_n352_), .A3(KEYINPUT3), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n354_), .B1(G141gat), .B2(G148gat), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G141gat), .A2(G148gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(KEYINPUT86), .A2(KEYINPUT2), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(KEYINPUT86), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n360_));
  OR2_X1    g159(.A1(KEYINPUT86), .A2(KEYINPUT2), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n359_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n350_), .B1(new_n356_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(G155gat), .ZN(new_n364_));
  INV_X1    g163(.A(G162gat), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT1), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT1), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n367_), .A2(G155gat), .A3(G162gat), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n366_), .B(new_n368_), .C1(G155gat), .C2(G162gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(G141gat), .B(G148gat), .Z(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n363_), .A2(new_n371_), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n372_), .A2(KEYINPUT29), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT28), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G22gat), .B(G50gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  OR2_X1    g175(.A1(new_n373_), .A2(KEYINPUT28), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n373_), .A2(KEYINPUT28), .ZN(new_n378_));
  INV_X1    g177(.A(new_n375_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n377_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n376_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(G197gat), .ZN(new_n382_));
  OR3_X1    g181(.A1(new_n382_), .A2(KEYINPUT89), .A3(G204gat), .ZN(new_n383_));
  AOI21_X1  g182(.A(KEYINPUT89), .B1(new_n382_), .B2(G204gat), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n382_), .A2(G204gat), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n383_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G211gat), .B(G218gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT90), .ZN(new_n388_));
  OR2_X1    g187(.A1(G211gat), .A2(G218gat), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT90), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G211gat), .A2(G218gat), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n389_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n388_), .A2(KEYINPUT21), .A3(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(G197gat), .B(G204gat), .Z(new_n394_));
  AOI22_X1  g193(.A1(new_n388_), .A2(new_n392_), .B1(new_n394_), .B2(KEYINPUT21), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT21), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n383_), .B(new_n396_), .C1(new_n385_), .C2(new_n384_), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n386_), .A2(new_n393_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n398_), .A2(KEYINPUT88), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n372_), .A2(KEYINPUT29), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G78gat), .B(G106gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT91), .ZN(new_n403_));
  INV_X1    g202(.A(G233gat), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT87), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n405_), .A2(G228gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(G228gat), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n404_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n403_), .B(new_n408_), .ZN(new_n409_));
  OR2_X1    g208(.A1(new_n401_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n401_), .A2(new_n409_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n381_), .A2(new_n412_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n376_), .A2(new_n410_), .A3(new_n380_), .A4(new_n411_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G169gat), .A2(G176gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT22), .B(G169gat), .ZN(new_n417_));
  INV_X1    g216(.A(G176gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT23), .ZN(new_n420_));
  AND3_X1   g219(.A1(KEYINPUT80), .A2(G183gat), .A3(G190gat), .ZN(new_n421_));
  AOI21_X1  g220(.A(KEYINPUT80), .B1(G183gat), .B2(G190gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n420_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G183gat), .A2(G190gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT23), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n423_), .A2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(G183gat), .A2(G190gat), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n416_), .B(new_n419_), .C1(new_n427_), .C2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT26), .B(G190gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(KEYINPUT25), .B(G183gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(G169gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n418_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n434_), .A2(KEYINPUT24), .A3(new_n416_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n432_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT92), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT92), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n432_), .A2(new_n438_), .A3(new_n435_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT24), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n440_), .A2(new_n433_), .A3(new_n418_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT23), .B1(new_n421_), .B2(new_n422_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT81), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n444_), .B1(new_n424_), .B2(KEYINPUT23), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n444_), .B(KEYINPUT23), .C1(new_n421_), .C2(new_n422_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n442_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT93), .ZN(new_n449_));
  OAI211_X1 g248(.A(new_n437_), .B(new_n439_), .C1(new_n448_), .C2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT80), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n424_), .A2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(KEYINPUT80), .A2(G183gat), .A3(G190gat), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n420_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n445_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n447_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n441_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n457_), .A2(KEYINPUT93), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n398_), .B(new_n429_), .C1(new_n450_), .C2(new_n458_), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n435_), .A2(new_n441_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT26), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(KEYINPUT79), .A3(G190gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(KEYINPUT79), .A2(G190gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT26), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n431_), .A2(new_n462_), .A3(new_n464_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n460_), .A2(new_n423_), .A3(new_n426_), .A4(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n428_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n419_), .A2(new_n416_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n466_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n395_), .A2(new_n397_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n386_), .A2(KEYINPUT21), .A3(new_n388_), .A4(new_n392_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(KEYINPUT98), .B(KEYINPUT20), .Z(new_n474_));
  NAND3_X1  g273(.A1(new_n459_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G226gat), .A2(G233gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT19), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n429_), .B1(new_n450_), .B2(new_n458_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(new_n472_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n477_), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT20), .B1(new_n469_), .B2(new_n472_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n480_), .A2(new_n481_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n478_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G8gat), .B(G36gat), .ZN(new_n486_));
  INV_X1    g285(.A(G92gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT18), .B(G64gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT32), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n485_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G225gat), .A2(G233gat), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  OR2_X1    g294(.A1(G127gat), .A2(G134gat), .ZN(new_n496_));
  INV_X1    g295(.A(G120gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(G113gat), .ZN(new_n498_));
  INV_X1    g297(.A(G113gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(G120gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G127gat), .A2(G134gat), .ZN(new_n501_));
  AND4_X1   g300(.A1(new_n496_), .A2(new_n498_), .A3(new_n500_), .A4(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  AOI22_X1  g302(.A1(new_n498_), .A2(new_n500_), .B1(new_n496_), .B2(new_n501_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  AOI22_X1  g304(.A1(new_n363_), .A2(new_n371_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT94), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n502_), .A2(new_n504_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n508_), .A2(new_n363_), .A3(new_n371_), .ZN(new_n509_));
  AOI22_X1  g308(.A1(new_n506_), .A2(new_n507_), .B1(new_n509_), .B2(KEYINPUT4), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n353_), .A2(new_n355_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(KEYINPUT86), .A2(KEYINPUT2), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n512_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n511_), .A2(new_n513_), .A3(new_n360_), .ZN(new_n514_));
  AOI22_X1  g313(.A1(new_n514_), .A2(new_n350_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT4), .ZN(new_n516_));
  NOR4_X1   g315(.A1(new_n515_), .A2(KEYINPUT94), .A3(new_n508_), .A4(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n495_), .B1(new_n510_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n508_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n372_), .A2(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n520_), .A2(new_n506_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(new_n494_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n518_), .A2(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(G1gat), .B(G29gat), .Z(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(G85gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT0), .B(G57gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n523_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n518_), .A2(new_n522_), .A3(new_n527_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n457_), .A2(KEYINPUT93), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n448_), .A2(new_n449_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n532_), .A2(new_n533_), .A3(new_n437_), .A4(new_n439_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n398_), .B1(new_n534_), .B2(new_n429_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n477_), .B1(new_n535_), .B2(new_n482_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n481_), .A2(KEYINPUT20), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n459_), .A2(new_n473_), .A3(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(new_n538_), .A3(new_n491_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n493_), .A2(new_n531_), .A3(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n527_), .B1(new_n521_), .B2(new_n495_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT96), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n509_), .A2(KEYINPUT4), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n372_), .A2(new_n519_), .A3(new_n507_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n372_), .A2(new_n519_), .A3(new_n507_), .A4(KEYINPUT4), .ZN(new_n546_));
  AOI211_X1 g345(.A(new_n542_), .B(new_n495_), .C1(new_n545_), .C2(new_n546_), .ZN(new_n547_));
  NOR3_X1   g346(.A1(new_n515_), .A2(KEYINPUT94), .A3(new_n508_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n516_), .B1(new_n515_), .B2(new_n508_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n546_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT96), .B1(new_n550_), .B2(new_n494_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n541_), .B1(new_n547_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT97), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(KEYINPUT95), .A2(KEYINPUT33), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n530_), .A2(new_n556_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n518_), .A2(new_n522_), .A3(new_n527_), .A4(new_n555_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  OAI211_X1 g358(.A(KEYINPUT97), .B(new_n541_), .C1(new_n547_), .C2(new_n551_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n554_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n490_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n481_), .B1(new_n480_), .B2(new_n483_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n538_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n562_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n482_), .B1(new_n472_), .B2(new_n479_), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n490_), .B(new_n538_), .C1(new_n566_), .C2(new_n481_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n415_), .B(new_n540_), .C1(new_n561_), .C2(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n508_), .B(KEYINPUT31), .Z(new_n570_));
  INV_X1    g369(.A(new_n428_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n468_), .B1(new_n456_), .B2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n465_), .A2(new_n441_), .A3(new_n435_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n573_), .A2(new_n427_), .ZN(new_n574_));
  OAI21_X1  g373(.A(KEYINPUT30), .B1(new_n572_), .B2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G15gat), .B(G43gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G71gat), .B(G99gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT30), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n466_), .B(new_n579_), .C1(new_n467_), .C2(new_n468_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n575_), .A2(new_n578_), .A3(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n578_), .B1(new_n575_), .B2(new_n580_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT82), .B(KEYINPUT83), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G227gat), .A2(G233gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NOR3_X1   g385(.A1(new_n581_), .A2(new_n582_), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n575_), .A2(new_n580_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n578_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n575_), .A2(new_n578_), .A3(new_n580_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n585_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(KEYINPUT84), .B1(new_n587_), .B2(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n586_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n590_), .A2(new_n585_), .A3(new_n591_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT84), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n594_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n570_), .B1(new_n593_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n570_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n587_), .A2(new_n592_), .A3(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(KEYINPUT85), .B1(new_n598_), .B2(new_n600_), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n594_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n596_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n599_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT85), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n569_), .A2(new_n601_), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n567_), .A2(KEYINPUT27), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n490_), .B1(new_n478_), .B2(new_n484_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(KEYINPUT27), .B1(new_n565_), .B2(new_n567_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n531_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n415_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(KEYINPUT99), .B1(new_n607_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n415_), .ZN(new_n616_));
  NOR3_X1   g415(.A1(new_n616_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n600_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n605_), .B1(new_n604_), .B2(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n598_), .A2(KEYINPUT85), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n617_), .B(new_n613_), .C1(new_n619_), .C2(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n619_), .A2(new_n620_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT99), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n485_), .A2(new_n562_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n624_), .A2(KEYINPUT27), .A3(new_n567_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT27), .ZN(new_n626_));
  INV_X1    g425(.A(new_n567_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n490_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n626_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n625_), .A2(new_n629_), .A3(new_n613_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(new_n616_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n622_), .A2(new_n623_), .A3(new_n631_), .A4(new_n569_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n615_), .A2(new_n621_), .A3(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n349_), .A2(new_n633_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n311_), .A2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n531_), .B(KEYINPUT100), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n635_), .A2(new_n216_), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT38), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n292_), .B1(new_n301_), .B2(new_n300_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(new_n303_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n243_), .A2(new_n642_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n643_), .A2(new_n634_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(G1gat), .B1(new_n645_), .B2(new_n613_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n637_), .A2(new_n638_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n639_), .A2(new_n646_), .A3(new_n647_), .ZN(G1324gat));
  INV_X1    g447(.A(new_n612_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n635_), .A2(new_n217_), .A3(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(G8gat), .B1(new_n645_), .B2(new_n612_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n651_), .A2(KEYINPUT39), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n651_), .A2(KEYINPUT39), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n650_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT40), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(G1325gat));
  OAI21_X1  g455(.A(G15gat), .B1(new_n645_), .B2(new_n622_), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n657_), .A2(KEYINPUT41), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(KEYINPUT41), .ZN(new_n659_));
  INV_X1    g458(.A(G15gat), .ZN(new_n660_));
  INV_X1    g459(.A(new_n622_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n635_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n658_), .A2(new_n659_), .A3(new_n662_), .ZN(G1326gat));
  INV_X1    g462(.A(G22gat), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n415_), .B(KEYINPUT101), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n635_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n665_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G22gat), .B1(new_n645_), .B2(new_n667_), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n668_), .A2(KEYINPUT103), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(KEYINPUT103), .ZN(new_n670_));
  XNOR2_X1  g469(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n669_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n666_), .B1(new_n672_), .B2(new_n673_), .ZN(G1327gat));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n675_));
  OAI21_X1  g474(.A(KEYINPUT43), .B1(new_n309_), .B2(new_n675_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n633_), .A2(new_n310_), .A3(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n633_), .B2(new_n310_), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n349_), .B(new_n243_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n633_), .A2(new_n310_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n676_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n633_), .A2(new_n310_), .A3(new_n676_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n680_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n686_), .A2(new_n349_), .A3(new_n243_), .A4(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n681_), .A2(new_n688_), .A3(new_n636_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G29gat), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n242_), .A2(new_n641_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n634_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(G29gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(new_n693_), .A3(new_n531_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n690_), .A2(new_n694_), .ZN(G1328gat));
  INV_X1    g494(.A(KEYINPUT46), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n696_), .A2(KEYINPUT108), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(KEYINPUT108), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT109), .Z(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n612_), .A2(G36gat), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n692_), .A2(new_n701_), .ZN(new_n702_));
  XOR2_X1   g501(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n692_), .A2(new_n701_), .A3(new_n703_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n681_), .A2(new_n688_), .A3(new_n649_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(G36gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n707_), .B1(new_n709_), .B2(KEYINPUT106), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n708_), .A2(new_n711_), .A3(G36gat), .ZN(new_n712_));
  AOI211_X1 g511(.A(new_n697_), .B(new_n700_), .C1(new_n710_), .C2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n709_), .A2(KEYINPUT106), .ZN(new_n714_));
  INV_X1    g513(.A(new_n707_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n714_), .A2(new_n712_), .A3(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n697_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n699_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n713_), .A2(new_n718_), .ZN(G1329gat));
  NAND4_X1  g518(.A1(new_n681_), .A2(new_n688_), .A3(G43gat), .A4(new_n661_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT110), .ZN(new_n721_));
  AOI21_X1  g520(.A(G43gat), .B1(new_n692_), .B2(new_n661_), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT111), .Z(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT47), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n721_), .A2(new_n723_), .A3(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1330gat));
  INV_X1    g527(.A(G50gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n681_), .A2(new_n688_), .A3(new_n616_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT112), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n729_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n732_), .B1(new_n731_), .B2(new_n730_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n692_), .A2(new_n729_), .A3(new_n665_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1331gat));
  AND3_X1   g534(.A1(new_n633_), .A2(new_n348_), .A3(new_n332_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n643_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(G57gat), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n737_), .A2(new_n738_), .A3(new_n613_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n636_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n311_), .A2(new_n736_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n741_), .B2(KEYINPUT113), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n742_), .B1(KEYINPUT113), .B2(new_n741_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n739_), .B1(new_n743_), .B2(new_n738_), .ZN(G1332gat));
  OAI21_X1  g543(.A(G64gat), .B1(new_n737_), .B2(new_n612_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT48), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n612_), .A2(G64gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n741_), .B2(new_n747_), .ZN(G1333gat));
  OAI21_X1  g547(.A(G71gat), .B1(new_n737_), .B2(new_n622_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT49), .ZN(new_n750_));
  OR2_X1    g549(.A1(new_n622_), .A2(G71gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n741_), .B2(new_n751_), .ZN(G1334gat));
  OAI21_X1  g551(.A(G78gat), .B1(new_n737_), .B2(new_n667_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT50), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n667_), .A2(G78gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n754_), .B1(new_n741_), .B2(new_n755_), .ZN(G1335gat));
  OR2_X1    g555(.A1(new_n686_), .A2(KEYINPUT115), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n686_), .A2(KEYINPUT115), .ZN(new_n758_));
  INV_X1    g557(.A(new_n332_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n242_), .A2(new_n759_), .A3(new_n347_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n757_), .A2(new_n758_), .A3(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n762_), .A2(G85gat), .A3(new_n531_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n736_), .A2(new_n691_), .ZN(new_n764_));
  AOI21_X1  g563(.A(G85gat), .B1(new_n764_), .B2(new_n636_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT114), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n763_), .A2(new_n766_), .ZN(G1336gat));
  AOI21_X1  g566(.A(G92gat), .B1(new_n764_), .B2(new_n649_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n612_), .A2(new_n487_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(new_n762_), .B2(new_n769_), .ZN(G1337gat));
  OAI21_X1  g569(.A(G99gat), .B1(new_n761_), .B2(new_n622_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n255_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n764_), .A2(new_n772_), .A3(new_n661_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g574(.A(G106gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n764_), .A2(new_n776_), .A3(new_n616_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n759_), .A2(new_n347_), .A3(new_n415_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n686_), .A2(new_n243_), .A3(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT116), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n776_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n781_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n782_), .B1(new_n781_), .B2(new_n783_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n777_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g586(.A1(new_n242_), .A2(new_n759_), .A3(new_n348_), .A4(new_n309_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n788_), .B(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n314_), .A2(new_n321_), .A3(new_n316_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n793_));
  AOI211_X1 g592(.A(KEYINPUT55), .B(new_n321_), .C1(new_n314_), .C2(new_n316_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n791_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n330_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT117), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT56), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n328_), .A2(new_n347_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n799_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(KEYINPUT117), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n800_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n338_), .A2(new_n334_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n333_), .A2(new_n336_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n344_), .B(new_n805_), .C1(new_n806_), .C2(new_n334_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n345_), .A2(new_n807_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n331_), .A2(new_n808_), .ZN(new_n809_));
  OAI211_X1 g608(.A(KEYINPUT57), .B(new_n641_), .C1(new_n804_), .C2(new_n809_), .ZN(new_n810_));
  XOR2_X1   g609(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n811_));
  AOI22_X1  g610(.A1(new_n800_), .A2(new_n803_), .B1(new_n331_), .B2(new_n808_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n812_), .B2(new_n642_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n810_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT121), .ZN(new_n816_));
  INV_X1    g615(.A(new_n791_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n319_), .A2(KEYINPUT55), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n317_), .A2(new_n792_), .A3(new_n318_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n817_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(KEYINPUT56), .B1(new_n820_), .B2(new_n330_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n795_), .A2(new_n799_), .A3(new_n796_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n808_), .A2(new_n328_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n821_), .A2(new_n822_), .A3(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT58), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT120), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n823_), .B1(new_n797_), .B2(KEYINPUT56), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT120), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n828_), .A2(new_n829_), .A3(KEYINPUT58), .A4(new_n822_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT58), .B1(new_n828_), .B2(new_n822_), .ZN(new_n831_));
  OAI21_X1  g630(.A(KEYINPUT119), .B1(new_n831_), .B2(new_n309_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n825_), .A2(new_n826_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n834_), .A3(new_n310_), .ZN(new_n835_));
  AOI221_X4 g634(.A(new_n816_), .B1(new_n827_), .B2(new_n830_), .C1(new_n832_), .C2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n832_), .A2(new_n835_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n827_), .A2(new_n830_), .ZN(new_n838_));
  AOI21_X1  g637(.A(KEYINPUT121), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n815_), .B1(new_n836_), .B2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n790_), .B1(new_n840_), .B2(new_n243_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n661_), .A2(new_n617_), .A3(new_n636_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(G113gat), .B1(new_n843_), .B2(new_n347_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n845_));
  INV_X1    g644(.A(new_n790_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n834_), .B1(new_n833_), .B2(new_n310_), .ZN(new_n847_));
  AOI211_X1 g646(.A(KEYINPUT119), .B(new_n309_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n838_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n816_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n837_), .A2(KEYINPUT121), .A3(new_n838_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n814_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n846_), .B1(new_n852_), .B2(new_n242_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n842_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n845_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n242_), .B1(new_n815_), .B2(new_n849_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n845_), .B(new_n854_), .C1(new_n856_), .C2(new_n790_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n855_), .A2(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n348_), .A2(new_n499_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n844_), .B1(new_n859_), .B2(new_n860_), .ZN(G1340gat));
  OAI21_X1  g660(.A(new_n497_), .B1(new_n759_), .B2(KEYINPUT60), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n843_), .B(new_n862_), .C1(KEYINPUT60), .C2(new_n497_), .ZN(new_n863_));
  AOI21_X1  g662(.A(KEYINPUT122), .B1(new_n859_), .B2(new_n332_), .ZN(new_n864_));
  OAI21_X1  g663(.A(KEYINPUT59), .B1(new_n841_), .B2(new_n842_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n865_), .A2(KEYINPUT122), .A3(new_n332_), .A4(new_n857_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(G120gat), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n863_), .B1(new_n864_), .B2(new_n867_), .ZN(G1341gat));
  AOI21_X1  g667(.A(G127gat), .B1(new_n843_), .B2(new_n242_), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n242_), .A2(G127gat), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n859_), .B2(new_n870_), .ZN(G1342gat));
  XNOR2_X1  g670(.A(KEYINPUT123), .B(G134gat), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n310_), .A2(new_n872_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n855_), .A2(new_n858_), .A3(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(G134gat), .B1(new_n843_), .B2(new_n642_), .ZN(new_n875_));
  OAI21_X1  g674(.A(KEYINPUT124), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n877_));
  INV_X1    g676(.A(G134gat), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n853_), .A2(new_n854_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n879_), .B2(new_n641_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n865_), .A2(new_n857_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n877_), .B(new_n880_), .C1(new_n881_), .C2(new_n873_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n876_), .A2(new_n882_), .ZN(G1343gat));
  NOR3_X1   g682(.A1(new_n841_), .A2(new_n415_), .A3(new_n661_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n649_), .A2(new_n740_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n884_), .A2(new_n347_), .A3(new_n885_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g686(.A1(new_n884_), .A2(new_n332_), .A3(new_n885_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g688(.A1(new_n884_), .A2(new_n242_), .A3(new_n885_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(KEYINPUT61), .B(G155gat), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1346gat));
  AND2_X1   g691(.A1(new_n884_), .A2(new_n885_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n309_), .A2(new_n365_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n884_), .A2(new_n642_), .A3(new_n885_), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n893_), .A2(new_n894_), .B1(new_n895_), .B2(new_n365_), .ZN(G1347gat));
  INV_X1    g695(.A(KEYINPUT62), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n856_), .A2(new_n790_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n622_), .A2(new_n612_), .A3(new_n636_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n667_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n898_), .A2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n347_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n897_), .B1(new_n902_), .B2(G169gat), .ZN(new_n903_));
  AOI211_X1 g702(.A(KEYINPUT62), .B(new_n433_), .C1(new_n901_), .C2(new_n347_), .ZN(new_n904_));
  OR3_X1    g703(.A1(new_n898_), .A2(KEYINPUT125), .A3(new_n900_), .ZN(new_n905_));
  OAI21_X1  g704(.A(KEYINPUT125), .B1(new_n898_), .B2(new_n900_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n347_), .A2(new_n417_), .ZN(new_n908_));
  OAI22_X1  g707(.A1(new_n903_), .A2(new_n904_), .B1(new_n907_), .B2(new_n908_), .ZN(G1348gat));
  NAND3_X1  g708(.A1(new_n905_), .A2(new_n906_), .A3(new_n332_), .ZN(new_n910_));
  AND3_X1   g709(.A1(new_n853_), .A2(new_n415_), .A3(new_n899_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n759_), .A2(new_n418_), .ZN(new_n912_));
  AOI22_X1  g711(.A1(new_n910_), .A2(new_n418_), .B1(new_n911_), .B2(new_n912_), .ZN(G1349gat));
  NOR3_X1   g712(.A1(new_n907_), .A2(new_n431_), .A3(new_n243_), .ZN(new_n914_));
  AOI21_X1  g713(.A(G183gat), .B1(new_n911_), .B2(new_n242_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1350gat));
  OAI21_X1  g715(.A(G190gat), .B1(new_n907_), .B2(new_n309_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n642_), .A2(new_n430_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n907_), .B2(new_n918_), .ZN(G1351gat));
  NOR2_X1   g718(.A1(new_n612_), .A2(new_n531_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n884_), .A2(new_n347_), .A3(new_n920_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g721(.A1(new_n884_), .A2(new_n332_), .A3(new_n920_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(G204gat), .ZN(G1353gat));
  NOR3_X1   g723(.A1(KEYINPUT126), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n925_));
  AOI211_X1 g724(.A(new_n925_), .B(new_n243_), .C1(KEYINPUT63), .C2(G211gat), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n884_), .A2(new_n920_), .A3(new_n926_), .ZN(new_n927_));
  OAI21_X1  g726(.A(KEYINPUT126), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n927_), .B(new_n929_), .ZN(G1354gat));
  AND2_X1   g729(.A1(new_n884_), .A2(new_n920_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(KEYINPUT127), .B(G218gat), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n309_), .A2(new_n932_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n884_), .A2(new_n642_), .A3(new_n920_), .ZN(new_n934_));
  AOI22_X1  g733(.A1(new_n931_), .A2(new_n933_), .B1(new_n934_), .B2(new_n932_), .ZN(G1355gat));
endmodule


