//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n856_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  INV_X1    g001(.A(G85gat), .ZN(new_n203_));
  INV_X1    g002(.A(G92gat), .ZN(new_n204_));
  NOR3_X1   g003(.A1(new_n203_), .A2(new_n204_), .A3(KEYINPUT9), .ZN(new_n205_));
  XOR2_X1   g004(.A(KEYINPUT10), .B(G99gat), .Z(new_n206_));
  INV_X1    g005(.A(G106gat), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n205_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(G85gat), .B(G92gat), .Z(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT9), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT6), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n208_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n214_));
  OR3_X1    g013(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n212_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT8), .ZN(new_n217_));
  AND3_X1   g016(.A1(new_n216_), .A2(new_n217_), .A3(new_n209_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n217_), .B1(new_n216_), .B2(new_n209_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n213_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G57gat), .B(G64gat), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n221_), .A2(KEYINPUT11), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(KEYINPUT11), .ZN(new_n223_));
  XOR2_X1   g022(.A(G71gat), .B(G78gat), .Z(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n223_), .A2(new_n224_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n220_), .A2(new_n228_), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n227_), .B(new_n213_), .C1(new_n218_), .C2(new_n219_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G230gat), .A2(G233gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT64), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n231_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n229_), .A2(KEYINPUT12), .A3(new_n230_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT12), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n220_), .A2(new_n238_), .A3(new_n228_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n236_), .B1(new_n240_), .B2(new_n233_), .ZN(new_n241_));
  AOI211_X1 g040(.A(KEYINPUT65), .B(new_n234_), .C1(new_n237_), .C2(new_n239_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n235_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G120gat), .B(G148gat), .ZN(new_n244_));
  INV_X1    g043(.A(G204gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT5), .B(G176gat), .ZN(new_n247_));
  XOR2_X1   g046(.A(new_n246_), .B(new_n247_), .Z(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n243_), .A2(new_n249_), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n235_), .B(new_n248_), .C1(new_n241_), .C2(new_n242_), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n250_), .A2(KEYINPUT66), .A3(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(KEYINPUT66), .B1(new_n250_), .B2(new_n251_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n202_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n250_), .A2(new_n251_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n250_), .A2(KEYINPUT66), .A3(new_n251_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(KEYINPUT13), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n254_), .A2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G1gat), .B(G8gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT70), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G15gat), .B(G22gat), .ZN(new_n263_));
  INV_X1    g062(.A(G1gat), .ZN(new_n264_));
  INV_X1    g063(.A(G8gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT14), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n263_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n262_), .A2(new_n267_), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n261_), .A2(KEYINPUT70), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n261_), .A2(KEYINPUT70), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n269_), .A2(new_n266_), .A3(new_n263_), .A4(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G29gat), .B(G36gat), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G43gat), .B(G50gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n275_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n273_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n272_), .B(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n280_), .A2(G229gat), .A3(G233gat), .ZN(new_n281_));
  OR2_X1    g080(.A1(new_n281_), .A2(KEYINPUT73), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(KEYINPUT73), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n272_), .A2(new_n279_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT15), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n279_), .B(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n284_), .B1(new_n272_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G229gat), .A2(G233gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n282_), .A2(new_n283_), .A3(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G113gat), .B(G141gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(G197gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT74), .B(G169gat), .ZN(new_n293_));
  XOR2_X1   g092(.A(new_n292_), .B(new_n293_), .Z(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n290_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n290_), .A2(new_n295_), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n260_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G155gat), .A2(G162gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT1), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT1), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n304_), .A2(G155gat), .A3(G162gat), .ZN(new_n305_));
  OR2_X1    g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n303_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(G141gat), .ZN(new_n308_));
  INV_X1    g107(.A(G148gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G141gat), .A2(G148gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n307_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT3), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT2), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n311_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n318_));
  AND4_X1   g117(.A1(new_n313_), .A2(new_n315_), .A3(new_n317_), .A4(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT84), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n306_), .A2(new_n320_), .A3(new_n302_), .ZN(new_n321_));
  AND2_X1   g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322_));
  NOR2_X1   g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT84), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n321_), .A2(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n312_), .B1(new_n319_), .B2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G127gat), .B(G134gat), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G113gat), .B(G120gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  XOR2_X1   g129(.A(G113gat), .B(G120gat), .Z(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(new_n327_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n326_), .A2(new_n333_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n315_), .A2(new_n317_), .A3(new_n313_), .A4(new_n318_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(new_n324_), .A3(new_n321_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n336_), .A2(new_n330_), .A3(new_n332_), .A4(new_n312_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n334_), .A2(KEYINPUT4), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT92), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n336_), .A2(new_n312_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT4), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n339_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n338_), .A2(new_n342_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n334_), .A2(new_n339_), .A3(KEYINPUT4), .A4(new_n337_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G225gat), .A2(G233gat), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n334_), .A2(new_n346_), .A3(new_n337_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G1gat), .B(G29gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(G85gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT0), .B(G57gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n348_), .A2(new_n350_), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT94), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n349_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT95), .B1(new_n358_), .B2(new_n355_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT95), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n346_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n360_), .B(new_n354_), .C1(new_n361_), .C2(new_n349_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT94), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n358_), .A2(new_n363_), .A3(new_n355_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n357_), .A2(new_n359_), .A3(new_n362_), .A4(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT96), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n363_), .B1(new_n358_), .B2(new_n355_), .ZN(new_n368_));
  NOR4_X1   g167(.A1(new_n361_), .A2(KEYINPUT94), .A3(new_n349_), .A4(new_n354_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n370_), .A2(KEYINPUT96), .A3(new_n359_), .A4(new_n362_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n367_), .A2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G8gat), .B(G36gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(G92gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT18), .B(G64gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G197gat), .B(G204gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G211gat), .B(G218gat), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT21), .ZN(new_n379_));
  OR3_X1    g178(.A1(new_n377_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n245_), .A2(G197gat), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n245_), .A2(G197gat), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT21), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n377_), .A2(new_n379_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(new_n384_), .A3(new_n378_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n380_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G169gat), .A2(G176gat), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT78), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G183gat), .A2(G190gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT23), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT23), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n393_), .A2(G183gat), .A3(G190gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n395_), .B1(G183gat), .B2(G190gat), .ZN(new_n396_));
  INV_X1    g195(.A(G176gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n397_), .B1(new_n398_), .B2(KEYINPUT81), .ZN(new_n399_));
  INV_X1    g198(.A(G169gat), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT80), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT22), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT81), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n399_), .B1(new_n400_), .B2(new_n403_), .ZN(new_n404_));
  OAI211_X1 g203(.A(KEYINPUT81), .B(G169gat), .C1(new_n401_), .C2(new_n402_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n404_), .A2(KEYINPUT82), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(KEYINPUT82), .B1(new_n404_), .B2(new_n405_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n390_), .B(new_n396_), .C1(new_n407_), .C2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT24), .ZN(new_n410_));
  NOR2_X1   g209(.A1(G169gat), .A2(G176gat), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT77), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(KEYINPUT77), .B1(G169gat), .B2(G176gat), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n410_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n390_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n413_), .A2(new_n410_), .A3(new_n414_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT75), .ZN(new_n419_));
  INV_X1    g218(.A(G190gat), .ZN(new_n420_));
  OR3_X1    g219(.A1(new_n419_), .A2(new_n420_), .A3(KEYINPUT26), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT25), .B(G183gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT26), .B1(new_n419_), .B2(new_n420_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n421_), .A2(KEYINPUT76), .A3(new_n422_), .A4(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT76), .ZN(new_n426_));
  AOI22_X1  g225(.A1(new_n394_), .A2(KEYINPUT79), .B1(KEYINPUT23), .B2(new_n391_), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n394_), .A2(KEYINPUT79), .ZN(new_n428_));
  AOI22_X1  g227(.A1(new_n425_), .A2(new_n426_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n418_), .A2(new_n424_), .A3(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n387_), .B1(new_n409_), .B2(new_n430_), .ZN(new_n431_));
  AND2_X1   g230(.A1(new_n415_), .A2(new_n388_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n411_), .A2(new_n410_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n422_), .ZN(new_n434_));
  XOR2_X1   g233(.A(KEYINPUT26), .B(G190gat), .Z(new_n435_));
  OAI211_X1 g234(.A(new_n395_), .B(new_n433_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(G183gat), .A2(G190gat), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n437_), .B1(new_n428_), .B2(new_n427_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT22), .B(G169gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n397_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(new_n390_), .ZN(new_n441_));
  OAI22_X1  g240(.A1(new_n432_), .A2(new_n436_), .B1(new_n438_), .B2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT20), .B1(new_n442_), .B2(new_n386_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G226gat), .A2(G233gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT19), .ZN(new_n445_));
  NOR3_X1   g244(.A1(new_n431_), .A2(new_n443_), .A3(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(KEYINPUT91), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n409_), .A2(new_n430_), .A3(new_n387_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT20), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n449_), .B1(new_n442_), .B2(new_n386_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n447_), .B1(new_n448_), .B2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n376_), .B1(new_n446_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n448_), .A2(new_n450_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n447_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n430_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n396_), .A2(new_n390_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n408_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n457_), .B1(new_n458_), .B2(new_n406_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n386_), .B1(new_n456_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n443_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n445_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n460_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n376_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n455_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n452_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT27), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(G233gat), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n469_), .A2(KEYINPUT87), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(KEYINPUT87), .ZN(new_n471_));
  OAI21_X1  g270(.A(G228gat), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT88), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n386_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT29), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n476_), .B1(new_n336_), .B2(new_n312_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n473_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n326_), .A2(KEYINPUT29), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n479_), .A2(new_n474_), .A3(new_n472_), .A4(new_n386_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G78gat), .B(G106gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT89), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n478_), .A2(new_n480_), .A3(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n485_), .B1(new_n326_), .B2(KEYINPUT29), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G22gat), .B(G50gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n485_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n336_), .A2(new_n476_), .A3(new_n312_), .A4(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n486_), .A2(new_n487_), .A3(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n487_), .B1(new_n486_), .B2(new_n489_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n484_), .A2(new_n490_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n481_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n494_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n483_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n484_), .B1(new_n497_), .B2(KEYINPUT90), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT90), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n478_), .A2(new_n480_), .A3(new_n499_), .A4(new_n483_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(KEYINPUT86), .B1(new_n492_), .B2(new_n490_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n490_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT86), .ZN(new_n504_));
  NOR3_X1   g303(.A1(new_n503_), .A2(new_n504_), .A3(new_n491_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n496_), .B1(new_n501_), .B2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n376_), .B(KEYINPUT97), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n453_), .A2(new_n454_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n462_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n508_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n511_), .A2(new_n465_), .A3(KEYINPUT27), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n468_), .A2(new_n507_), .A3(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT98), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G227gat), .A2(G233gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT31), .ZN(new_n517_));
  XOR2_X1   g316(.A(KEYINPUT30), .B(G15gat), .Z(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G71gat), .B(G99gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT83), .B(G43gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(new_n333_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n456_), .A2(new_n459_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n468_), .A2(new_n507_), .A3(new_n512_), .A4(KEYINPUT98), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n372_), .A2(new_n515_), .A3(new_n526_), .A4(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n468_), .A2(new_n512_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n507_), .B1(new_n372_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n525_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n524_), .B(new_n532_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n464_), .A2(KEYINPUT32), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n534_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n535_));
  OR3_X1    g334(.A1(new_n446_), .A2(new_n451_), .A3(new_n534_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n365_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  NOR3_X1   g336(.A1(new_n361_), .A2(new_n349_), .A3(new_n354_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT33), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n347_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n540_), .A2(KEYINPUT93), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n334_), .A2(new_n337_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n355_), .B1(new_n542_), .B2(new_n347_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n543_), .B1(new_n540_), .B2(KEYINPUT93), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n452_), .B(new_n465_), .C1(new_n541_), .C2(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n507_), .B1(new_n539_), .B2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n533_), .B1(new_n537_), .B2(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n528_), .B1(new_n531_), .B2(new_n547_), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n301_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G231gat), .A2(G233gat), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n268_), .A2(new_n271_), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n550_), .B1(new_n268_), .B2(new_n271_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n227_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n553_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n555_), .A2(new_n228_), .A3(new_n551_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT72), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n554_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G183gat), .B(G211gat), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n559_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n554_), .A2(new_n556_), .A3(new_n557_), .A4(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT71), .B(KEYINPUT16), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G127gat), .B(G155gat), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n564_), .B(new_n565_), .Z(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n566_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n560_), .A2(new_n562_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(KEYINPUT17), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT17), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n554_), .A2(new_n556_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n567_), .A2(new_n572_), .A3(new_n573_), .A4(new_n569_), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n571_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT69), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n576_), .A2(KEYINPUT37), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(KEYINPUT37), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G232gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT34), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n580_), .A2(KEYINPUT35), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n581_), .B1(new_n220_), .B2(new_n286_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n582_), .B1(new_n279_), .B2(new_n220_), .ZN(new_n583_));
  AOI21_X1  g382(.A(KEYINPUT68), .B1(new_n220_), .B2(new_n286_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n580_), .A2(KEYINPUT35), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT67), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n583_), .A2(new_n587_), .ZN(new_n588_));
  OAI221_X1 g387(.A(new_n582_), .B1(new_n279_), .B2(new_n220_), .C1(new_n584_), .C2(new_n586_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G190gat), .B(G218gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G134gat), .B(G162gat), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n590_), .B(new_n591_), .Z(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n593_), .A2(KEYINPUT36), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n588_), .A2(new_n589_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n592_), .B(KEYINPUT36), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n598_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n577_), .B(new_n578_), .C1(new_n596_), .C2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n599_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n601_), .A2(new_n576_), .A3(KEYINPUT37), .A4(new_n595_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n575_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n549_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n372_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n606_), .A2(new_n264_), .A3(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT38), .ZN(new_n609_));
  AOI21_X1  g408(.A(KEYINPUT99), .B1(new_n260_), .B2(new_n299_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT99), .ZN(new_n612_));
  AOI211_X1 g411(.A(new_n612_), .B(new_n298_), .C1(new_n254_), .C2(new_n259_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n601_), .A2(new_n595_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT100), .Z(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n548_), .A2(new_n617_), .A3(new_n575_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n611_), .A2(new_n614_), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT101), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n611_), .A2(new_n614_), .A3(KEYINPUT101), .A4(new_n618_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n623_), .A2(new_n607_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n609_), .B1(new_n264_), .B2(new_n624_), .ZN(G1324gat));
  NAND3_X1  g424(.A1(new_n606_), .A2(new_n265_), .A3(new_n529_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n611_), .A2(new_n614_), .A3(new_n529_), .A4(new_n618_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n627_), .A2(KEYINPUT102), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT39), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n265_), .B1(new_n627_), .B2(KEYINPUT102), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n628_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n629_), .B1(new_n628_), .B2(new_n630_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n626_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT40), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(G1325gat));
  NAND2_X1  g434(.A1(new_n623_), .A2(new_n526_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(G15gat), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n637_), .A2(KEYINPUT41), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(KEYINPUT41), .ZN(new_n639_));
  INV_X1    g438(.A(G15gat), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n606_), .A2(new_n640_), .A3(new_n526_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n638_), .A2(new_n639_), .A3(new_n641_), .ZN(G1326gat));
  INV_X1    g441(.A(G22gat), .ZN(new_n643_));
  INV_X1    g442(.A(new_n507_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n606_), .A2(new_n643_), .A3(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n621_), .A2(new_n644_), .A3(new_n622_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT42), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n646_), .A2(new_n647_), .A3(G22gat), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n647_), .B1(new_n646_), .B2(G22gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n645_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(G1327gat));
  NOR2_X1   g451(.A1(new_n575_), .A2(new_n615_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n549_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(G29gat), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n655_), .A3(new_n607_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n610_), .A2(new_n613_), .A3(new_n575_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n603_), .A2(KEYINPUT43), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n548_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(KEYINPUT105), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT105), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n548_), .A2(new_n661_), .A3(new_n658_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT104), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n603_), .B1(new_n548_), .B2(new_n665_), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n528_), .B(KEYINPUT104), .C1(new_n531_), .C2(new_n547_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n664_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n657_), .B1(new_n663_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  OAI211_X1 g470(.A(new_n657_), .B(KEYINPUT44), .C1(new_n668_), .C2(new_n663_), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n671_), .A2(new_n607_), .A3(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n656_), .B1(new_n673_), .B2(new_n655_), .ZN(G1328gat));
  XNOR2_X1  g473(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n671_), .A2(new_n529_), .A3(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(G36gat), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n529_), .B(KEYINPUT106), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n679_), .A2(G36gat), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n301_), .A2(new_n548_), .A3(new_n653_), .A4(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT45), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n677_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT107), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n675_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n682_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n676_), .B2(G36gat), .ZN(new_n687_));
  INV_X1    g486(.A(new_n675_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n687_), .A2(KEYINPUT107), .A3(new_n688_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n685_), .A2(new_n689_), .ZN(G1329gat));
  NAND4_X1  g489(.A1(new_n671_), .A2(G43gat), .A3(new_n526_), .A4(new_n672_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n654_), .A2(new_n526_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(KEYINPUT109), .B(G43gat), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n691_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g494(.A(G50gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n654_), .A2(new_n696_), .A3(new_n644_), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n671_), .A2(new_n644_), .A3(new_n672_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n697_), .B1(new_n698_), .B2(new_n696_), .ZN(G1331gat));
  NAND2_X1  g498(.A1(new_n548_), .A2(new_n298_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT110), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n254_), .A2(new_n259_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n701_), .A2(new_n702_), .A3(new_n605_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT111), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT112), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT111), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n703_), .B(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT112), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n705_), .A2(new_n709_), .A3(new_n607_), .ZN(new_n710_));
  INV_X1    g509(.A(G57gat), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n618_), .A2(new_n298_), .A3(new_n702_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n372_), .A2(new_n711_), .ZN(new_n713_));
  AOI22_X1  g512(.A1(new_n710_), .A2(new_n711_), .B1(new_n712_), .B2(new_n713_), .ZN(G1332gat));
  INV_X1    g513(.A(G64gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n712_), .B2(new_n678_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT48), .Z(new_n717_));
  NAND2_X1  g516(.A1(new_n678_), .A2(new_n715_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT113), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n717_), .B1(new_n707_), .B2(new_n719_), .ZN(G1333gat));
  INV_X1    g519(.A(G71gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n721_), .B1(new_n712_), .B2(new_n526_), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT49), .Z(new_n723_));
  NAND2_X1  g522(.A1(new_n526_), .A2(new_n721_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n723_), .B1(new_n707_), .B2(new_n724_), .ZN(G1334gat));
  INV_X1    g524(.A(G78gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n726_), .B1(new_n712_), .B2(new_n644_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT50), .Z(new_n728_));
  NAND2_X1  g527(.A1(new_n644_), .A2(new_n726_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n707_), .B2(new_n729_), .ZN(G1335gat));
  NAND3_X1  g529(.A1(new_n701_), .A2(new_n702_), .A3(new_n653_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(G85gat), .B1(new_n732_), .B2(new_n607_), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n663_), .A2(new_n668_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n575_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n702_), .A2(new_n298_), .A3(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT114), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n734_), .A2(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n372_), .A2(new_n203_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n733_), .B1(new_n738_), .B2(new_n739_), .ZN(G1336gat));
  AOI21_X1  g539(.A(G92gat), .B1(new_n732_), .B2(new_n529_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n679_), .A2(new_n204_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n738_), .B2(new_n742_), .ZN(G1337gat));
  INV_X1    g542(.A(G99gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(new_n738_), .B2(new_n526_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT51), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n746_), .A2(KEYINPUT115), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n732_), .A2(new_n206_), .A3(new_n526_), .ZN(new_n748_));
  OR3_X1    g547(.A1(new_n745_), .A2(new_n747_), .A3(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n747_), .B1(new_n745_), .B2(new_n748_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1338gat));
  NAND3_X1  g550(.A1(new_n732_), .A2(new_n207_), .A3(new_n644_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n734_), .A2(new_n644_), .A3(new_n737_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n753_), .A2(new_n754_), .A3(G106gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n753_), .B2(G106gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n752_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT53), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT53), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n752_), .B(new_n759_), .C1(new_n755_), .C2(new_n756_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1339gat));
  NOR2_X1   g560(.A1(new_n604_), .A2(new_n299_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT54), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n762_), .A2(new_n260_), .A3(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n762_), .B2(new_n260_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT55), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n767_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n240_), .A2(KEYINPUT116), .A3(new_n234_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n234_), .A2(KEYINPUT116), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n237_), .A2(new_n239_), .A3(new_n770_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n769_), .B(new_n771_), .C1(KEYINPUT55), .C2(new_n234_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n248_), .B1(new_n768_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT56), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n251_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  AOI211_X1 g574(.A(KEYINPUT56), .B(new_n248_), .C1(new_n768_), .C2(new_n772_), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n775_), .A2(new_n298_), .A3(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n280_), .A2(new_n288_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n287_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n295_), .B(new_n778_), .C1(new_n779_), .C2(new_n288_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n296_), .A2(new_n780_), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n252_), .A2(new_n253_), .A3(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n615_), .B1(new_n777_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT57), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n775_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n781_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n776_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n786_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT58), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n603_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n786_), .A2(KEYINPUT58), .A3(new_n787_), .A4(new_n788_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n791_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  OAI211_X1 g593(.A(KEYINPUT57), .B(new_n615_), .C1(new_n777_), .C2(new_n782_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n785_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n766_), .B1(new_n796_), .B2(new_n735_), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n515_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n798_), .A2(new_n607_), .ZN(new_n799_));
  OR2_X1    g598(.A1(new_n799_), .A2(KEYINPUT117), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(KEYINPUT117), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n797_), .A2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(G113gat), .B1(new_n803_), .B2(new_n299_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n802_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT59), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n796_), .A2(new_n735_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n766_), .B1(new_n808_), .B2(KEYINPUT118), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT118), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n796_), .A2(new_n810_), .A3(new_n735_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n807_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n766_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n808_), .A2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n806_), .B1(new_n814_), .B2(new_n805_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n812_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT119), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n817_), .A2(G113gat), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n299_), .A2(KEYINPUT119), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n818_), .B1(new_n819_), .B2(G113gat), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n804_), .B1(new_n816_), .B2(new_n820_), .ZN(G1340gat));
  INV_X1    g620(.A(G120gat), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n822_), .B1(new_n260_), .B2(KEYINPUT60), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n803_), .B(new_n823_), .C1(KEYINPUT60), .C2(new_n822_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(KEYINPUT120), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n812_), .A2(new_n815_), .A3(new_n260_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(new_n822_), .ZN(G1341gat));
  AOI21_X1  g626(.A(G127gat), .B1(new_n803_), .B2(new_n575_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n575_), .A2(G127gat), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n816_), .B2(new_n829_), .ZN(G1342gat));
  INV_X1    g629(.A(KEYINPUT122), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n797_), .A2(new_n617_), .A3(new_n802_), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT121), .B1(new_n832_), .B2(G134gat), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT121), .ZN(new_n834_));
  INV_X1    g633(.A(G134gat), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n814_), .A2(new_n805_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n834_), .B(new_n835_), .C1(new_n836_), .C2(new_n617_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n833_), .A2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n603_), .A2(new_n835_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n812_), .A2(new_n815_), .A3(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n831_), .B1(new_n838_), .B2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n809_), .A2(new_n811_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n807_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n815_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n846_), .A3(new_n839_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n847_), .A2(KEYINPUT122), .A3(new_n837_), .A4(new_n833_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n842_), .A2(new_n848_), .ZN(G1343gat));
  NOR3_X1   g648(.A1(new_n797_), .A2(new_n507_), .A3(new_n526_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n678_), .A2(new_n372_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n299_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n702_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT123), .B(G148gat), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1345gat));
  NOR2_X1   g656(.A1(new_n526_), .A2(new_n507_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n814_), .A2(new_n575_), .A3(new_n858_), .A4(new_n851_), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n859_), .A2(KEYINPUT124), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(KEYINPUT124), .ZN(new_n861_));
  XNOR2_X1  g660(.A(KEYINPUT61), .B(G155gat), .ZN(new_n862_));
  AND3_X1   g661(.A1(new_n860_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n862_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n863_), .A2(new_n864_), .ZN(G1346gat));
  AOI21_X1  g664(.A(G162gat), .B1(new_n852_), .B2(new_n616_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n792_), .A2(G162gat), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n852_), .B2(new_n867_), .ZN(G1347gat));
  XOR2_X1   g667(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n679_), .A2(new_n607_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n533_), .A2(new_n644_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n843_), .A2(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n298_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n870_), .B1(new_n876_), .B2(new_n400_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n439_), .ZN(new_n878_));
  OAI211_X1 g677(.A(G169gat), .B(new_n869_), .C1(new_n875_), .C2(new_n298_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n877_), .A2(new_n878_), .A3(new_n879_), .ZN(G1348gat));
  INV_X1    g679(.A(new_n875_), .ZN(new_n881_));
  AOI21_X1  g680(.A(G176gat), .B1(new_n881_), .B2(new_n702_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n873_), .A2(new_n397_), .A3(new_n260_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n814_), .B2(new_n883_), .ZN(G1349gat));
  NOR2_X1   g683(.A1(new_n873_), .A2(new_n735_), .ZN(new_n885_));
  AOI21_X1  g684(.A(G183gat), .B1(new_n766_), .B2(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n735_), .A2(new_n422_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n886_), .B1(new_n881_), .B2(new_n887_), .ZN(G1350gat));
  OAI21_X1  g687(.A(G190gat), .B1(new_n875_), .B2(new_n603_), .ZN(new_n889_));
  OR2_X1    g688(.A1(new_n617_), .A2(new_n435_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n875_), .B2(new_n890_), .ZN(G1351gat));
  AND2_X1   g690(.A1(new_n850_), .A2(new_n871_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n299_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n702_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g695(.A(new_n735_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n892_), .A2(new_n897_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(KEYINPUT126), .B(KEYINPUT127), .ZN(new_n899_));
  NOR2_X1   g698(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n899_), .B(new_n900_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n898_), .B(new_n901_), .ZN(G1354gat));
  AOI21_X1  g701(.A(G218gat), .B1(new_n892_), .B2(new_n616_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n792_), .A2(G218gat), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n903_), .B1(new_n892_), .B2(new_n904_), .ZN(G1355gat));
endmodule


