//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n579_, new_n580_, new_n581_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n618_, new_n619_, new_n620_, new_n622_,
    new_n623_, new_n624_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n772_, new_n774_, new_n775_, new_n777_, new_n778_, new_n779_,
    new_n781_, new_n783_, new_n784_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n832_, new_n833_,
    new_n834_, new_n836_, new_n837_, new_n838_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n863_;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(new_n202_), .B1(new_n203_), .B2(KEYINPUT23), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(KEYINPUT81), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  MUX2_X1   g006(.A(new_n204_), .B(new_n202_), .S(new_n207_), .Z(new_n208_));
  OAI21_X1  g007(.A(new_n208_), .B1(G183gat), .B2(G190gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT80), .ZN(new_n211_));
  XOR2_X1   g010(.A(KEYINPUT22), .B(G169gat), .Z(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G176gat), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n211_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  NOR3_X1   g014(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n205_), .A2(new_n206_), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n218_), .A2(KEYINPUT82), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n203_), .A2(KEYINPUT23), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n220_), .B1(new_n218_), .B2(KEYINPUT82), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n217_), .B1(new_n219_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT83), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT25), .B(G183gat), .ZN(new_n225_));
  INV_X1    g024(.A(G190gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT26), .B1(new_n226_), .B2(KEYINPUT79), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  NOR3_X1   g027(.A1(new_n226_), .A2(KEYINPUT79), .A3(KEYINPUT26), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n230_));
  OAI22_X1  g029(.A1(new_n228_), .A2(new_n229_), .B1(new_n211_), .B2(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n231_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n232_));
  AOI22_X1  g031(.A1(new_n209_), .A2(new_n215_), .B1(new_n224_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G227gat), .A2(G233gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(G15gat), .B(G43gat), .Z(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G127gat), .B(G134gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G113gat), .B(G120gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n238_), .A2(new_n239_), .ZN(new_n241_));
  MUX2_X1   g040(.A(new_n240_), .B(new_n241_), .S(KEYINPUT86), .Z(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT31), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G71gat), .B(G99gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT85), .B(KEYINPUT30), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n243_), .B(new_n246_), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n237_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n237_), .A2(new_n247_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G197gat), .B(G204gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G211gat), .B(G218gat), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT21), .ZN(new_n253_));
  OR3_X1    g052(.A1(new_n251_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n251_), .A2(new_n253_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n252_), .B1(new_n251_), .B2(new_n253_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n254_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  XOR2_X1   g056(.A(G155gat), .B(G162gat), .Z(new_n258_));
  OR2_X1    g057(.A1(G141gat), .A2(G148gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT2), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G141gat), .A2(G148gat), .ZN(new_n261_));
  AOI22_X1  g060(.A1(new_n259_), .A2(KEYINPUT3), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n262_), .B1(KEYINPUT3), .B2(new_n259_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT87), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n258_), .B1(new_n263_), .B2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT88), .ZN(new_n267_));
  NOR2_X1   g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G155gat), .A2(G162gat), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n268_), .B1(KEYINPUT1), .B2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n270_), .B1(KEYINPUT1), .B2(new_n269_), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n271_), .A2(new_n259_), .A3(new_n261_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n267_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT29), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n257_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G22gat), .B(G50gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT28), .ZN(new_n277_));
  XOR2_X1   g076(.A(G78gat), .B(G106gat), .Z(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n275_), .B(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n273_), .A2(new_n274_), .ZN(new_n281_));
  AND2_X1   g080(.A1(KEYINPUT89), .A2(G233gat), .ZN(new_n282_));
  NOR2_X1   g081(.A1(KEYINPUT89), .A2(G233gat), .ZN(new_n283_));
  OAI21_X1  g082(.A(G228gat), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n284_), .B(KEYINPUT90), .Z(new_n285_));
  XNOR2_X1  g084(.A(new_n281_), .B(new_n285_), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n280_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n280_), .A2(new_n286_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n250_), .A2(new_n289_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n273_), .A2(new_n240_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n291_), .A2(KEYINPUT92), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n273_), .A2(new_n242_), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n292_), .B1(new_n294_), .B2(KEYINPUT92), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G225gat), .A2(G233gat), .ZN(new_n296_));
  AOI21_X1  g095(.A(KEYINPUT93), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n296_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT4), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n299_), .B1(new_n273_), .B2(new_n242_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n300_), .B1(new_n295_), .B2(new_n299_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n297_), .B1(new_n298_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(KEYINPUT94), .B(KEYINPUT0), .Z(new_n304_));
  XNOR2_X1  g103(.A(G1gat), .B(G29gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G57gat), .B(G85gat), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n306_), .B(new_n307_), .Z(new_n308_));
  INV_X1    g107(.A(KEYINPUT93), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n301_), .A2(new_n309_), .A3(new_n298_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n303_), .A2(new_n308_), .A3(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n311_), .A2(KEYINPUT95), .A3(KEYINPUT33), .ZN(new_n312_));
  INV_X1    g111(.A(new_n310_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n313_), .A2(new_n302_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(KEYINPUT95), .A2(KEYINPUT33), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(KEYINPUT95), .A2(KEYINPUT33), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n314_), .A2(new_n308_), .A3(new_n316_), .A4(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n312_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT91), .ZN(new_n320_));
  INV_X1    g119(.A(new_n257_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n233_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT26), .B(G190gat), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n216_), .B1(new_n225_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n210_), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n208_), .B(new_n324_), .C1(new_n325_), .C2(new_n230_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n219_), .A2(new_n221_), .ZN(new_n327_));
  INV_X1    g126(.A(G183gat), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n327_), .B1(new_n328_), .B2(new_n226_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n215_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n326_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT20), .B1(new_n331_), .B2(new_n257_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n322_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G226gat), .A2(G233gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT19), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n333_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n233_), .A2(new_n321_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT20), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n339_), .B1(new_n331_), .B2(new_n257_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(new_n335_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n320_), .B1(new_n337_), .B2(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(KEYINPUT91), .B1(new_n333_), .B2(new_n336_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G8gat), .B(G36gat), .ZN(new_n346_));
  INV_X1    g145(.A(G92gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT18), .B(G64gat), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n348_), .B(new_n349_), .Z(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n345_), .B(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n301_), .A2(new_n296_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n308_), .B1(new_n295_), .B2(new_n298_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n352_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n319_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT96), .ZN(new_n357_));
  INV_X1    g156(.A(new_n308_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n358_), .B1(new_n313_), .B2(new_n302_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n311_), .A2(new_n357_), .A3(new_n359_), .ZN(new_n360_));
  OAI211_X1 g159(.A(KEYINPUT96), .B(new_n358_), .C1(new_n313_), .C2(new_n302_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n351_), .A2(KEYINPUT32), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n345_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n338_), .A2(new_n340_), .A3(new_n336_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n364_), .B1(new_n333_), .B2(new_n336_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(KEYINPUT32), .A3(new_n351_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n360_), .A2(new_n361_), .A3(new_n363_), .A4(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n290_), .B1(new_n356_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n360_), .A2(new_n361_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n250_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n289_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n289_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n250_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT27), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n345_), .A2(new_n351_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n375_), .B1(new_n365_), .B2(new_n350_), .ZN(new_n377_));
  AOI22_X1  g176(.A1(new_n352_), .A2(new_n375_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n369_), .A2(new_n374_), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n368_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT12), .ZN(new_n382_));
  OR2_X1    g181(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n383_));
  INV_X1    g182(.A(G85gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n347_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G85gat), .A2(G92gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n383_), .A2(new_n385_), .A3(new_n386_), .A4(new_n387_), .ZN(new_n388_));
  AND3_X1   g187(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n389_));
  AOI21_X1  g188(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT64), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G99gat), .A2(G106gat), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT6), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT64), .ZN(new_n395_));
  NAND3_X1  g194(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n391_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT7), .ZN(new_n399_));
  INV_X1    g198(.A(G99gat), .ZN(new_n400_));
  INV_X1    g199(.A(G106gat), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n388_), .B1(new_n398_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT8), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n402_), .A2(new_n394_), .A3(new_n396_), .A4(new_n403_), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n385_), .A2(new_n386_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT66), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n406_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n407_), .A2(KEYINPUT66), .A3(new_n408_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n405_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n385_), .A2(KEYINPUT9), .A3(new_n386_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT10), .B(G99gat), .ZN(new_n415_));
  OAI221_X1 g214(.A(new_n414_), .B1(KEYINPUT9), .B2(new_n386_), .C1(new_n415_), .C2(G106gat), .ZN(new_n416_));
  INV_X1    g215(.A(new_n398_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n382_), .B1(new_n413_), .B2(new_n418_), .ZN(new_n419_));
  XOR2_X1   g218(.A(G71gat), .B(G78gat), .Z(new_n420_));
  AND2_X1   g219(.A1(G57gat), .A2(G64gat), .ZN(new_n421_));
  NOR2_X1   g220(.A1(G57gat), .A2(G64gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT11), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(G57gat), .ZN(new_n424_));
  INV_X1    g223(.A(G64gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT11), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G57gat), .A2(G64gat), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n426_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n420_), .A2(new_n423_), .A3(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G71gat), .B(G78gat), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n431_), .B(KEYINPUT11), .C1(new_n422_), .C2(new_n421_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n430_), .A2(new_n432_), .A3(new_n434_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n413_), .A2(new_n438_), .A3(new_n418_), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n430_), .A2(new_n432_), .A3(new_n434_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n434_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n409_), .A2(new_n410_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n443_), .A2(KEYINPUT8), .A3(new_n412_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n405_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n418_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n442_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n419_), .B1(new_n439_), .B2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT70), .B(KEYINPUT12), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n418_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n450_), .B1(new_n451_), .B2(new_n442_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT71), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G230gat), .A2(G233gat), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT71), .ZN(new_n455_));
  OAI211_X1 g254(.A(new_n455_), .B(new_n450_), .C1(new_n451_), .C2(new_n442_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n449_), .A2(new_n453_), .A3(new_n454_), .A4(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n451_), .A2(new_n442_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n438_), .B1(new_n413_), .B2(new_n418_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n454_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT69), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT69), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n460_), .A2(new_n464_), .A3(new_n461_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n457_), .A2(new_n463_), .A3(new_n465_), .ZN(new_n466_));
  XOR2_X1   g265(.A(G120gat), .B(G148gat), .Z(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(G204gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT5), .B(G176gat), .ZN(new_n469_));
  XOR2_X1   g268(.A(new_n468_), .B(new_n469_), .Z(new_n470_));
  NOR2_X1   g269(.A1(new_n470_), .A2(KEYINPUT72), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n466_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n463_), .A2(new_n465_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n457_), .ZN(new_n474_));
  NOR3_X1   g273(.A1(new_n473_), .A2(new_n474_), .A3(new_n471_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n472_), .A2(new_n475_), .ZN(new_n476_));
  OR2_X1    g275(.A1(new_n476_), .A2(KEYINPUT13), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(KEYINPUT13), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G229gat), .A2(G233gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G1gat), .B(G8gat), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT73), .B(G15gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(G22gat), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT14), .ZN(new_n485_));
  XNOR2_X1  g284(.A(KEYINPUT74), .B(G1gat), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n485_), .B1(new_n486_), .B2(G8gat), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n482_), .B1(new_n484_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(G22gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n483_), .B(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n487_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n481_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n488_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(G43gat), .B(G50gat), .Z(new_n495_));
  XNOR2_X1  g294(.A(G29gat), .B(G36gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n494_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G43gat), .B(G50gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n496_), .B(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n493_), .A2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n480_), .B1(new_n498_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT77), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n500_), .A2(KEYINPUT15), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n500_), .A2(KEYINPUT15), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n492_), .B(new_n488_), .C1(new_n504_), .C2(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n503_), .B1(new_n506_), .B2(new_n501_), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n504_), .A2(new_n505_), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT77), .B1(new_n508_), .B2(new_n494_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n480_), .B(KEYINPUT78), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n502_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(G169gat), .B(G197gat), .Z(new_n514_));
  XNOR2_X1  g313(.A(G113gat), .B(G141gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n513_), .B(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n479_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G231gat), .A2(G233gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n438_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(new_n493_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT76), .ZN(new_n523_));
  XOR2_X1   g322(.A(G183gat), .B(G211gat), .Z(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G127gat), .B(G155gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n525_), .B(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT17), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n522_), .A2(new_n530_), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(KEYINPUT17), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n446_), .A2(new_n447_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n508_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G232gat), .A2(G233gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT34), .ZN(new_n538_));
  OAI221_X1 g337(.A(new_n536_), .B1(KEYINPUT35), .B2(new_n538_), .C1(new_n497_), .C2(new_n535_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(KEYINPUT35), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n539_), .B(new_n540_), .Z(new_n541_));
  XNOR2_X1  g340(.A(G190gat), .B(G218gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G134gat), .B(G162gat), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n542_), .B(new_n543_), .Z(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT36), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n541_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n539_), .B(new_n540_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT36), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n547_), .A2(new_n548_), .A3(new_n544_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n546_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT37), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n534_), .A2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n381_), .A2(new_n519_), .A3(new_n553_), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n369_), .A2(new_n486_), .ZN(new_n555_));
  OR3_X1    g354(.A1(new_n554_), .A2(KEYINPUT97), .A3(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT97), .B1(new_n554_), .B2(new_n555_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n558_), .A2(KEYINPUT38), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n550_), .B(KEYINPUT98), .Z(new_n560_));
  NOR2_X1   g359(.A1(new_n534_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n381_), .A2(new_n519_), .A3(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(G1gat), .B1(new_n562_), .B2(new_n369_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n558_), .A2(KEYINPUT38), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n559_), .A2(new_n563_), .A3(new_n564_), .ZN(G1324gat));
  NOR3_X1   g364(.A1(new_n554_), .A2(G8gat), .A3(new_n378_), .ZN(new_n566_));
  OAI21_X1  g365(.A(G8gat), .B1(new_n562_), .B2(new_n378_), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n567_), .A2(KEYINPUT39), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(KEYINPUT39), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n566_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n570_), .B(new_n572_), .ZN(G1325gat));
  OAI21_X1  g372(.A(G15gat), .B1(new_n562_), .B2(new_n250_), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n574_), .A2(KEYINPUT41), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(KEYINPUT41), .ZN(new_n576_));
  OR3_X1    g375(.A1(new_n554_), .A2(G15gat), .A3(new_n250_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .ZN(G1326gat));
  OAI21_X1  g377(.A(G22gat), .B1(new_n562_), .B2(new_n289_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT42), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n372_), .A2(new_n489_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n580_), .B1(new_n554_), .B2(new_n581_), .ZN(G1327gat));
  INV_X1    g381(.A(new_n534_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n583_), .A2(new_n550_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n381_), .A2(KEYINPUT100), .A3(new_n519_), .A4(new_n584_), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n519_), .B(new_n584_), .C1(new_n368_), .C2(new_n380_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT100), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n585_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n369_), .ZN(new_n591_));
  AOI21_X1  g390(.A(G29gat), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(G29gat), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n534_), .A2(new_n519_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n552_), .B1(new_n368_), .B2(new_n380_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(KEYINPUT43), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT43), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n597_), .B(new_n552_), .C1(new_n368_), .C2(new_n380_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n594_), .B1(new_n596_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT44), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n593_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n599_), .A2(KEYINPUT44), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n592_), .B1(new_n602_), .B2(new_n604_), .ZN(G1328gat));
  INV_X1    g404(.A(new_n378_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n606_), .B1(new_n599_), .B2(KEYINPUT44), .ZN(new_n607_));
  OAI21_X1  g406(.A(G36gat), .B1(new_n603_), .B2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n378_), .A2(G36gat), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n585_), .A2(new_n588_), .A3(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(KEYINPUT101), .B(KEYINPUT45), .Z(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT102), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n610_), .B(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(KEYINPUT103), .B(KEYINPUT46), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n608_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n614_), .B1(new_n608_), .B2(new_n613_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(G1329gat));
  OAI211_X1 g416(.A(G43gat), .B(new_n370_), .C1(new_n599_), .C2(KEYINPUT44), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n589_), .A2(new_n250_), .ZN(new_n619_));
  OAI22_X1  g418(.A1(new_n618_), .A2(new_n603_), .B1(new_n619_), .B2(G43gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g420(.A(G50gat), .B1(new_n590_), .B2(new_n372_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n372_), .A2(G50gat), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n623_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n622_), .B1(new_n624_), .B2(new_n604_), .ZN(G1331gat));
  INV_X1    g424(.A(new_n479_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n626_), .A2(new_n517_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n381_), .A2(new_n561_), .A3(new_n627_), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n628_), .A2(new_n424_), .A3(new_n369_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n381_), .A2(new_n627_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(new_n553_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(new_n591_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n629_), .B1(new_n633_), .B2(new_n424_), .ZN(G1332gat));
  OAI21_X1  g433(.A(G64gat), .B1(new_n628_), .B2(new_n378_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT48), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n632_), .A2(new_n425_), .A3(new_n606_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(G1333gat));
  OAI21_X1  g437(.A(G71gat), .B1(new_n628_), .B2(new_n250_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT105), .ZN(new_n640_));
  XNOR2_X1  g439(.A(KEYINPUT104), .B(KEYINPUT49), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n642_), .ZN(new_n644_));
  OR3_X1    g443(.A1(new_n631_), .A2(G71gat), .A3(new_n250_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n643_), .A2(new_n644_), .A3(new_n645_), .ZN(G1334gat));
  OAI21_X1  g445(.A(G78gat), .B1(new_n628_), .B2(new_n289_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT50), .ZN(new_n648_));
  OR3_X1    g447(.A1(new_n631_), .A2(G78gat), .A3(new_n289_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(KEYINPUT106), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT106), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n648_), .A2(new_n652_), .A3(new_n649_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(G1335gat));
  NAND2_X1  g453(.A1(new_n630_), .A2(new_n584_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(G85gat), .B1(new_n656_), .B2(new_n591_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n627_), .A2(new_n534_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT107), .Z(new_n659_));
  AOI21_X1  g458(.A(new_n659_), .B1(new_n596_), .B2(new_n598_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n369_), .A2(new_n384_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n657_), .B1(new_n660_), .B2(new_n661_), .ZN(G1336gat));
  AOI21_X1  g461(.A(G92gat), .B1(new_n656_), .B2(new_n606_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n378_), .A2(new_n347_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n660_), .B2(new_n664_), .ZN(G1337gat));
  OR3_X1    g464(.A1(new_n655_), .A2(new_n415_), .A3(new_n250_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n660_), .A2(new_n370_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n666_), .B1(new_n400_), .B2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(KEYINPUT51), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT51), .ZN(new_n670_));
  OAI211_X1 g469(.A(new_n666_), .B(new_n670_), .C1(new_n400_), .C2(new_n667_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(G1338gat));
  NAND3_X1  g471(.A1(new_n656_), .A2(new_n401_), .A3(new_n372_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT52), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n660_), .A2(new_n372_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n675_), .B2(G106gat), .ZN(new_n676_));
  AOI211_X1 g475(.A(KEYINPUT52), .B(new_n401_), .C1(new_n660_), .C2(new_n372_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n673_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT53), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT53), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n680_), .B(new_n673_), .C1(new_n676_), .C2(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(G1339gat));
  NAND4_X1  g481(.A1(new_n532_), .A2(new_n518_), .A3(new_n533_), .A4(new_n551_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n683_), .A2(new_n479_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT108), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n684_), .A2(new_n685_), .A3(KEYINPUT54), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n685_), .A2(KEYINPUT54), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(KEYINPUT54), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n687_), .B(new_n688_), .C1(new_n683_), .C2(new_n479_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n686_), .A2(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(KEYINPUT112), .A2(KEYINPUT58), .ZN(new_n691_));
  AOI22_X1  g490(.A1(new_n458_), .A2(new_n459_), .B1(new_n535_), .B2(new_n382_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n456_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n455_), .B1(new_n459_), .B2(new_n450_), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n692_), .A2(new_n693_), .A3(new_n694_), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n695_), .A2(KEYINPUT109), .A3(KEYINPUT55), .A4(new_n454_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT109), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT55), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n697_), .B1(new_n457_), .B2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n449_), .A2(new_n456_), .A3(new_n453_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n461_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n457_), .A2(new_n698_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n696_), .A2(new_n699_), .A3(new_n701_), .A4(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n470_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT56), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n703_), .A2(KEYINPUT56), .A3(new_n704_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n510_), .A2(new_n511_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n498_), .A2(new_n501_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n516_), .B1(new_n711_), .B2(new_n512_), .ZN(new_n712_));
  AOI22_X1  g511(.A1(new_n513_), .A2(new_n516_), .B1(new_n710_), .B2(new_n712_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n457_), .A2(new_n463_), .A3(new_n470_), .A4(new_n465_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT111), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n713_), .A2(KEYINPUT111), .A3(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n691_), .B1(new_n709_), .B2(new_n719_), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n703_), .A2(KEYINPUT56), .A3(new_n704_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT56), .B1(new_n703_), .B2(new_n704_), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n719_), .B(new_n691_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n552_), .B1(new_n720_), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT113), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n546_), .A2(KEYINPUT110), .A3(new_n549_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n517_), .A2(new_n714_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n713_), .B1(new_n472_), .B2(new_n475_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT110), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n729_), .B2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT57), .ZN(new_n733_));
  INV_X1    g532(.A(new_n728_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n734_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n731_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT57), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n737_), .A2(new_n738_), .A3(new_n727_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n733_), .A2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n719_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n691_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n551_), .B1(new_n743_), .B2(new_n723_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT113), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n726_), .A2(new_n740_), .A3(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT114), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n583_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n726_), .A2(new_n740_), .A3(new_n746_), .A4(KEYINPUT114), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n690_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n606_), .A2(new_n369_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n752_), .A2(new_n370_), .A3(new_n289_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n751_), .A2(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(G113gat), .B1(new_n754_), .B2(new_n517_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n583_), .B1(new_n740_), .B2(new_n725_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n690_), .A2(new_n756_), .ZN(new_n757_));
  OR3_X1    g556(.A1(new_n757_), .A2(KEYINPUT59), .A3(new_n753_), .ZN(new_n758_));
  OAI21_X1  g557(.A(KEYINPUT59), .B1(new_n751_), .B2(new_n753_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n517_), .A2(G113gat), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT115), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n755_), .B1(new_n761_), .B2(new_n763_), .ZN(G1340gat));
  OAI21_X1  g563(.A(G120gat), .B1(new_n760_), .B2(new_n626_), .ZN(new_n765_));
  INV_X1    g564(.A(G120gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n766_), .B1(new_n626_), .B2(KEYINPUT60), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n754_), .B(new_n767_), .C1(KEYINPUT60), .C2(new_n766_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n765_), .A2(new_n768_), .ZN(G1341gat));
  NAND2_X1  g568(.A1(new_n583_), .A2(G127gat), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n751_), .A2(new_n534_), .A3(new_n753_), .ZN(new_n771_));
  OAI22_X1  g570(.A1(new_n760_), .A2(new_n770_), .B1(G127gat), .B2(new_n771_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT116), .ZN(G1342gat));
  AOI21_X1  g572(.A(G134gat), .B1(new_n754_), .B2(new_n560_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n552_), .A2(G134gat), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n761_), .B2(new_n775_), .ZN(G1343gat));
  NOR2_X1   g575(.A1(new_n751_), .A2(new_n373_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n777_), .A2(new_n752_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n517_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n479_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g581(.A1(new_n778_), .A2(new_n583_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(KEYINPUT61), .B(G155gat), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n783_), .B(new_n784_), .ZN(G1346gat));
  NAND2_X1  g584(.A1(new_n778_), .A2(new_n560_), .ZN(new_n786_));
  INV_X1    g585(.A(G162gat), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n788_), .A2(KEYINPUT117), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n778_), .A2(G162gat), .A3(new_n552_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n790_), .B1(new_n788_), .B2(KEYINPUT117), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n789_), .A2(new_n791_), .ZN(G1347gat));
  NOR2_X1   g591(.A1(new_n591_), .A2(new_n378_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n370_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n289_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n796_), .A2(new_n757_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n517_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n798_), .A2(G169gat), .ZN(new_n799_));
  OR2_X1    g598(.A1(new_n799_), .A2(KEYINPUT62), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(KEYINPUT62), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n800_), .B(new_n801_), .C1(new_n212_), .C2(new_n798_), .ZN(G1348gat));
  INV_X1    g601(.A(KEYINPUT119), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n803_), .B1(new_n751_), .B2(new_n372_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n738_), .B1(new_n737_), .B2(new_n727_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n727_), .ZN(new_n806_));
  AOI211_X1 g605(.A(KEYINPUT57), .B(new_n806_), .C1(new_n735_), .C2(new_n736_), .ZN(new_n807_));
  OAI22_X1  g606(.A1(new_n805_), .A2(new_n807_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n725_), .A2(KEYINPUT113), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n748_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(new_n534_), .A3(new_n750_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n690_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n813_), .A2(KEYINPUT119), .A3(new_n289_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n626_), .A2(new_n214_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n804_), .A2(new_n814_), .A3(new_n795_), .A4(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT120), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n372_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n794_), .B1(new_n818_), .B2(KEYINPUT119), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT120), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n819_), .A2(new_n820_), .A3(new_n804_), .A4(new_n815_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n817_), .A2(new_n821_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n796_), .A2(new_n757_), .A3(new_n626_), .ZN(new_n823_));
  OR3_X1    g622(.A1(new_n823_), .A2(KEYINPUT118), .A3(G176gat), .ZN(new_n824_));
  OAI21_X1  g623(.A(KEYINPUT118), .B1(new_n823_), .B2(G176gat), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n822_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT121), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT121), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n822_), .A2(new_n829_), .A3(new_n826_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(G1349gat));
  INV_X1    g630(.A(new_n797_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n832_), .A2(new_n225_), .A3(new_n534_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n819_), .A2(new_n583_), .A3(new_n804_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n834_), .B2(new_n328_), .ZN(G1350gat));
  OAI21_X1  g634(.A(G190gat), .B1(new_n832_), .B2(new_n551_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n560_), .A2(new_n323_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(KEYINPUT122), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n836_), .B1(new_n832_), .B2(new_n838_), .ZN(G1351gat));
  NAND2_X1  g638(.A1(new_n777_), .A2(new_n793_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n517_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g642(.A1(new_n840_), .A2(new_n626_), .ZN(new_n844_));
  XOR2_X1   g643(.A(KEYINPUT123), .B(G204gat), .Z(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(G1353gat));
  AOI21_X1  g645(.A(new_n534_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n777_), .A2(KEYINPUT125), .A3(new_n793_), .A4(new_n847_), .ZN(new_n848_));
  OR2_X1    g647(.A1(new_n848_), .A2(KEYINPUT126), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(KEYINPUT126), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT125), .ZN(new_n852_));
  INV_X1    g651(.A(new_n847_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n840_), .B2(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT124), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n851_), .A2(new_n857_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n849_), .A2(new_n854_), .A3(new_n856_), .A4(new_n850_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(G1354gat));
  AOI21_X1  g659(.A(G218gat), .B1(new_n841_), .B2(new_n560_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n552_), .A2(G218gat), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT127), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n861_), .B1(new_n841_), .B2(new_n863_), .ZN(G1355gat));
endmodule


