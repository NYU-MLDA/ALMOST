//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1 1 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n793_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n829_, new_n830_, new_n831_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_, new_n938_, new_n939_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n954_,
    new_n955_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n965_, new_n966_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_,
    new_n997_, new_n998_, new_n1000_, new_n1001_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1016_, new_n1017_;
  NOR2_X1   g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT7), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n205_));
  AND2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT6), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT69), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT8), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT69), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n206_), .A2(new_n212_), .A3(new_n208_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G85gat), .B(G92gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n210_), .A2(new_n211_), .A3(new_n213_), .A4(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n209_), .A2(new_n215_), .ZN(new_n217_));
  AOI21_X1  g016(.A(KEYINPUT70), .B1(new_n217_), .B2(KEYINPUT8), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n214_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT70), .ZN(new_n220_));
  NOR3_X1   g019(.A1(new_n219_), .A2(new_n220_), .A3(new_n211_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n216_), .B1(new_n218_), .B2(new_n221_), .ZN(new_n222_));
  OR2_X1    g021(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n223_), .A2(KEYINPUT65), .A3(new_n224_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(G106gat), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT66), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(KEYINPUT67), .B(G92gat), .Z(new_n232_));
  AOI21_X1  g031(.A(KEYINPUT9), .B1(new_n232_), .B2(G85gat), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT68), .B1(G85gat), .B2(G92gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n208_), .B1(new_n233_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n238_));
  AOI211_X1 g037(.A(new_n238_), .B(G106gat), .C1(new_n227_), .C2(new_n228_), .ZN(new_n239_));
  OR3_X1    g038(.A1(new_n231_), .A2(new_n237_), .A3(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G57gat), .B(G64gat), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n241_), .A2(KEYINPUT11), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(KEYINPUT11), .ZN(new_n243_));
  XOR2_X1   g042(.A(G71gat), .B(G78gat), .Z(new_n244_));
  NAND3_X1  g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n243_), .A2(new_n244_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n222_), .A2(new_n240_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT71), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n222_), .A2(new_n240_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n247_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n222_), .A2(new_n240_), .A3(KEYINPUT71), .A4(new_n247_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n250_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G230gat), .A2(G233gat), .ZN(new_n256_));
  XOR2_X1   g055(.A(new_n256_), .B(KEYINPUT64), .Z(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n255_), .A2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n220_), .B1(new_n219_), .B2(new_n211_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n217_), .A2(KEYINPUT70), .A3(KEYINPUT8), .ZN(new_n261_));
  AND3_X1   g060(.A1(new_n213_), .A2(new_n211_), .A3(new_n215_), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n260_), .A2(new_n261_), .B1(new_n262_), .B2(new_n210_), .ZN(new_n263_));
  NOR3_X1   g062(.A1(new_n231_), .A2(new_n237_), .A3(new_n239_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT12), .ZN(new_n266_));
  OAI22_X1  g065(.A1(new_n265_), .A2(new_n247_), .B1(KEYINPUT72), .B2(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n258_), .B1(new_n265_), .B2(new_n247_), .ZN(new_n268_));
  XOR2_X1   g067(.A(KEYINPUT72), .B(KEYINPUT12), .Z(new_n269_));
  OAI211_X1 g068(.A(new_n252_), .B(new_n269_), .C1(new_n263_), .C2(new_n264_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n267_), .A2(new_n268_), .A3(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G120gat), .B(G148gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT5), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G176gat), .B(G204gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n273_), .B(new_n274_), .Z(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n259_), .A2(new_n271_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT73), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n259_), .A2(new_n271_), .A3(KEYINPUT73), .A4(new_n276_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n259_), .A2(new_n271_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(new_n275_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT13), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n281_), .A2(KEYINPUT13), .A3(new_n283_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT74), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT74), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n288_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G190gat), .B(G218gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G134gat), .B(G162gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n296_), .B(KEYINPUT36), .Z(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G29gat), .B(G36gat), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G43gat), .B(G50gat), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n299_), .A2(new_n301_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT75), .B(KEYINPUT15), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n303_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n305_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n251_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n303_), .A2(new_n304_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n265_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G232gat), .A2(G233gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT34), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT35), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n308_), .A2(new_n310_), .A3(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n313_), .A2(new_n314_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n317_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n308_), .A2(new_n310_), .A3(new_n319_), .A4(new_n315_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n298_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n296_), .A2(KEYINPUT36), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n318_), .A2(new_n322_), .A3(new_n320_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT76), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT76), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n318_), .A2(new_n325_), .A3(new_n322_), .A4(new_n320_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n321_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT37), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n327_), .A2(KEYINPUT37), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G15gat), .B(G22gat), .ZN(new_n331_));
  INV_X1    g130(.A(G1gat), .ZN(new_n332_));
  INV_X1    g131(.A(G8gat), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT14), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n331_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G1gat), .B(G8gat), .ZN(new_n336_));
  OR2_X1    g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n336_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G231gat), .A2(G233gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(new_n247_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G127gat), .B(G155gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT16), .ZN(new_n344_));
  XOR2_X1   g143(.A(G183gat), .B(G211gat), .Z(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT17), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n346_), .A2(new_n347_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n342_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n342_), .A2(new_n349_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n351_), .B1(new_n352_), .B2(KEYINPUT77), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n353_), .B1(KEYINPUT77), .B2(new_n351_), .ZN(new_n354_));
  NOR3_X1   g153(.A1(new_n329_), .A2(new_n330_), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n293_), .A2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT78), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT101), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT1), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT88), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT88), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n359_), .A2(new_n362_), .A3(KEYINPUT1), .ZN(new_n363_));
  OR2_X1    g162(.A1(G155gat), .A2(G162gat), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT1), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(G155gat), .A3(G162gat), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n361_), .A2(new_n363_), .A3(new_n364_), .A4(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(G141gat), .B(G148gat), .Z(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n364_), .A2(new_n359_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G141gat), .A2(G148gat), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT89), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT2), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n371_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT3), .ZN(new_n375_));
  INV_X1    g174(.A(G141gat), .ZN(new_n376_));
  INV_X1    g175(.A(G148gat), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n374_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n373_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n370_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n369_), .A2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n383_), .A2(KEYINPUT29), .ZN(new_n384_));
  XOR2_X1   g183(.A(G22gat), .B(G50gat), .Z(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n388_));
  INV_X1    g187(.A(new_n381_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n389_), .A2(new_n374_), .A3(new_n379_), .A4(new_n378_), .ZN(new_n390_));
  AOI22_X1  g189(.A1(new_n390_), .A2(new_n370_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT29), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n385_), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n387_), .A2(new_n388_), .A3(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n388_), .B1(new_n387_), .B2(new_n394_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G78gat), .B(G106gat), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n392_), .B1(new_n369_), .B2(new_n382_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT21), .ZN(new_n401_));
  INV_X1    g200(.A(G204gat), .ZN(new_n402_));
  INV_X1    g201(.A(G197gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT91), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT91), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(G197gat), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n402_), .B1(new_n404_), .B2(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(G197gat), .A2(G204gat), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n401_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(G218gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(G211gat), .ZN(new_n411_));
  INV_X1    g210(.A(G211gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(G218gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n404_), .A2(new_n406_), .A3(new_n402_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n401_), .B1(G197gat), .B2(G204gat), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n414_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n407_), .A2(new_n408_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n401_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n419_));
  AOI22_X1  g218(.A1(new_n409_), .A2(new_n417_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(G228gat), .ZN(new_n421_));
  INV_X1    g220(.A(G233gat), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NOR3_X1   g222(.A1(new_n400_), .A2(new_n420_), .A3(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n383_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n409_), .A2(new_n417_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n418_), .A2(new_n419_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n427_), .A2(KEYINPUT93), .A3(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(KEYINPUT93), .B1(new_n427_), .B2(new_n428_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n426_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  AOI211_X1 g230(.A(new_n399_), .B(new_n424_), .C1(new_n431_), .C2(new_n423_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n398_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n427_), .A2(new_n428_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT93), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n420_), .A2(KEYINPUT93), .ZN(new_n437_));
  AOI22_X1  g236(.A1(new_n436_), .A2(new_n437_), .B1(new_n383_), .B2(new_n425_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n423_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n434_), .A2(new_n439_), .ZN(new_n440_));
  OAI22_X1  g239(.A1(new_n438_), .A2(new_n439_), .B1(new_n400_), .B2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n441_), .A2(KEYINPUT96), .A3(new_n399_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n399_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT96), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n433_), .A2(new_n442_), .A3(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n424_), .B1(new_n431_), .B2(new_n423_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n399_), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT94), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n448_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n447_), .A2(KEYINPUT94), .A3(new_n448_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT95), .B1(new_n453_), .B2(new_n398_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT95), .ZN(new_n455_));
  AOI211_X1 g254(.A(new_n455_), .B(new_n397_), .C1(new_n451_), .C2(new_n452_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n446_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G1gat), .B(G29gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G57gat), .B(G85gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G225gat), .A2(G233gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G127gat), .B(G134gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G113gat), .B(G120gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT87), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n464_), .A2(new_n465_), .A3(KEYINPUT87), .ZN(new_n469_));
  XOR2_X1   g268(.A(G127gat), .B(G134gat), .Z(new_n470_));
  XOR2_X1   g269(.A(G113gat), .B(G120gat), .Z(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n468_), .A2(new_n469_), .A3(new_n472_), .ZN(new_n473_));
  NOR3_X1   g272(.A1(new_n391_), .A2(new_n473_), .A3(KEYINPUT4), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n466_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n369_), .A2(new_n475_), .A3(new_n382_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n476_), .B(KEYINPUT4), .C1(new_n391_), .C2(new_n473_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n474_), .B1(new_n477_), .B2(KEYINPUT98), .ZN(new_n478_));
  AND2_X1   g277(.A1(new_n472_), .A2(new_n469_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n383_), .A2(new_n468_), .A3(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT98), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n480_), .A2(new_n481_), .A3(KEYINPUT4), .A4(new_n476_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n463_), .B1(new_n478_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n463_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n484_), .B1(new_n480_), .B2(new_n476_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n462_), .B1(new_n483_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n477_), .A2(KEYINPUT98), .ZN(new_n487_));
  INV_X1    g286(.A(new_n474_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(new_n482_), .A3(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(new_n484_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n462_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n485_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n486_), .A2(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(G8gat), .B(G36gat), .Z(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT18), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G64gat), .B(G92gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n498_), .A2(KEYINPUT32), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT100), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G226gat), .A2(G233gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT19), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G183gat), .A2(G190gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT23), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT23), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n505_), .A2(G183gat), .A3(G190gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n507_), .B1(G183gat), .B2(G190gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G169gat), .A2(G176gat), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT22), .B(G169gat), .ZN(new_n511_));
  INV_X1    g310(.A(G176gat), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n510_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n508_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(G169gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n512_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n516_), .A2(KEYINPUT24), .A3(new_n509_), .ZN(new_n517_));
  OR3_X1    g316(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n507_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT26), .B(G190gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT25), .B(G183gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n514_), .B1(new_n519_), .B2(new_n523_), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n429_), .A2(new_n430_), .A3(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT86), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT85), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT22), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(G169gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n515_), .A2(KEYINPUT22), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n527_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n527_), .B1(new_n515_), .B2(KEYINPUT22), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n512_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n526_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(G176gat), .B1(new_n529_), .B2(new_n527_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n535_), .B(KEYINPUT86), .C1(new_n527_), .C2(new_n511_), .ZN(new_n536_));
  OR2_X1    g335(.A1(KEYINPUT83), .A2(G183gat), .ZN(new_n537_));
  INV_X1    g336(.A(G190gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(KEYINPUT83), .A2(G183gat), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n537_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n510_), .B1(new_n540_), .B2(new_n507_), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n534_), .A2(new_n536_), .A3(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n537_), .A2(new_n539_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT25), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n544_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT84), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n548_), .B1(new_n538_), .B2(KEYINPUT26), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(KEYINPUT26), .B(G190gat), .Z(new_n551_));
  AOI21_X1  g350(.A(new_n550_), .B1(new_n551_), .B2(KEYINPUT84), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n519_), .B1(new_n547_), .B2(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n434_), .B1(new_n542_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT20), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n500_), .B(new_n502_), .C1(new_n525_), .C2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n534_), .A2(new_n536_), .A3(new_n541_), .ZN(new_n557_));
  AND3_X1   g356(.A1(new_n507_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n537_), .A2(new_n539_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n543_), .B1(new_n559_), .B2(KEYINPUT25), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n549_), .B1(new_n520_), .B2(new_n548_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n558_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n420_), .A2(new_n557_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n558_), .A2(new_n522_), .B1(new_n508_), .B2(new_n513_), .ZN(new_n565_));
  OAI21_X1  g364(.A(KEYINPUT20), .B1(new_n565_), .B2(new_n420_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n502_), .B(KEYINPUT97), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n564_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n556_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n502_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n436_), .A2(new_n437_), .A3(new_n565_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT20), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n562_), .A2(new_n557_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n573_), .B1(new_n574_), .B2(new_n434_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n571_), .B1(new_n572_), .B2(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n576_), .A2(new_n500_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n499_), .B1(new_n570_), .B2(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n567_), .B1(new_n564_), .B2(new_n566_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n502_), .B1(new_n565_), .B2(new_n420_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n575_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n582_), .A2(new_n499_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n494_), .A2(new_n578_), .A3(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT33), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n485_), .B1(new_n489_), .B2(new_n484_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n585_), .B1(new_n586_), .B2(new_n491_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n498_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n571_), .B1(new_n434_), .B2(new_n524_), .ZN(new_n589_));
  AOI22_X1  g388(.A1(new_n562_), .A2(new_n557_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n590_));
  NOR3_X1   g389(.A1(new_n589_), .A2(new_n590_), .A3(new_n573_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n567_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n573_), .B1(new_n434_), .B2(new_n524_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n592_), .B1(new_n593_), .B2(new_n563_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n588_), .B1(new_n591_), .B2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n579_), .A2(new_n498_), .A3(new_n581_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  OAI211_X1 g397(.A(KEYINPUT33), .B(new_n462_), .C1(new_n483_), .C2(new_n485_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n478_), .A2(new_n463_), .A3(new_n482_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n480_), .A2(new_n476_), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n600_), .B(new_n491_), .C1(new_n463_), .C2(new_n601_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n587_), .A2(new_n598_), .A3(new_n599_), .A4(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n584_), .A2(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n358_), .B1(new_n457_), .B2(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n432_), .B1(new_n443_), .B2(KEYINPUT94), .ZN(new_n606_));
  INV_X1    g405(.A(new_n452_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n398_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(new_n455_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n453_), .A2(KEYINPUT95), .A3(new_n398_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n584_), .A2(new_n603_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n611_), .A2(KEYINPUT101), .A3(new_n446_), .A4(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT102), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n586_), .A2(new_n491_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n483_), .A2(new_n462_), .A3(new_n485_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n614_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n486_), .A2(new_n493_), .A3(KEYINPUT102), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(KEYINPUT27), .B1(new_n595_), .B2(new_n596_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n576_), .A2(new_n500_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n568_), .B1(new_n576_), .B2(new_n500_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n498_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n596_), .A2(KEYINPUT27), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n621_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n619_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n457_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n605_), .A2(new_n613_), .A3(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G227gat), .A2(G233gat), .ZN(new_n630_));
  INV_X1    g429(.A(G15gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT30), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n574_), .B(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(new_n473_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G71gat), .B(G99gat), .ZN(new_n636_));
  INV_X1    g435(.A(G43gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT31), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n635_), .B(new_n639_), .Z(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n617_), .A2(new_n618_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n588_), .B1(new_n570_), .B2(new_n577_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n625_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT103), .B1(new_n645_), .B2(new_n621_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT103), .ZN(new_n647_));
  AOI211_X1 g446(.A(new_n647_), .B(new_n620_), .C1(new_n643_), .C2(new_n644_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n642_), .B1(new_n646_), .B2(new_n648_), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n640_), .B(new_n446_), .C1(new_n454_), .C2(new_n456_), .ZN(new_n650_));
  OAI21_X1  g449(.A(KEYINPUT104), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n626_), .A2(new_n647_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n645_), .A2(KEYINPUT103), .A3(new_n621_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n619_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n446_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n655_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT104), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n654_), .A2(new_n656_), .A3(new_n657_), .A4(new_n640_), .ZN(new_n658_));
  AOI22_X1  g457(.A1(new_n629_), .A2(new_n641_), .B1(new_n651_), .B2(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n339_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n309_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(G229gat), .A2(G233gat), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(KEYINPUT79), .B1(new_n662_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT79), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n660_), .A2(new_n666_), .A3(new_n663_), .A4(new_n661_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n339_), .A2(new_n304_), .A3(new_n303_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(new_n661_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(new_n664_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(G113gat), .B(G141gat), .ZN(new_n671_));
  XNOR2_X1  g470(.A(G169gat), .B(G197gat), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n671_), .B(new_n672_), .Z(new_n673_));
  NAND4_X1  g472(.A1(new_n665_), .A2(new_n667_), .A3(new_n670_), .A4(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT80), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n670_), .A2(new_n667_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n677_), .A2(KEYINPUT80), .A3(new_n665_), .A4(new_n673_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n665_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n673_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n679_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT81), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n679_), .A2(KEYINPUT81), .A3(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT82), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n659_), .A2(new_n688_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT105), .Z(new_n690_));
  NAND2_X1  g489(.A1(new_n357_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n692_), .A2(new_n332_), .A3(new_n619_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT38), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n694_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n293_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n687_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n697_), .A2(new_n698_), .A3(new_n354_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n659_), .A2(new_n327_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G1gat), .B1(new_n701_), .B2(new_n642_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n695_), .A2(new_n696_), .A3(new_n702_), .ZN(G1324gat));
  NOR2_X1   g502(.A1(new_n646_), .A2(new_n648_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(G8gat), .B1(new_n701_), .B2(new_n705_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n706_), .A2(KEYINPUT39), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(KEYINPUT39), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n704_), .A2(new_n333_), .ZN(new_n709_));
  OAI22_X1  g508(.A1(new_n707_), .A2(new_n708_), .B1(new_n691_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT40), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  OAI221_X1 g511(.A(KEYINPUT40), .B1(new_n691_), .B2(new_n709_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1325gat));
  OAI21_X1  g513(.A(G15gat), .B1(new_n701_), .B2(new_n641_), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n715_), .A2(KEYINPUT41), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n692_), .A2(new_n631_), .A3(new_n640_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(KEYINPUT41), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n716_), .A2(new_n717_), .A3(new_n718_), .ZN(G1326gat));
  XNOR2_X1  g518(.A(new_n656_), .B(KEYINPUT106), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n699_), .A2(new_n700_), .A3(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(G22gat), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n723_), .A2(KEYINPUT42), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n723_), .A2(KEYINPUT42), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n720_), .A2(G22gat), .ZN(new_n726_));
  OAI22_X1  g525(.A1(new_n724_), .A2(new_n725_), .B1(new_n691_), .B2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT107), .ZN(G1327gat));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n329_), .A2(new_n330_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n629_), .A2(new_n641_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n651_), .A2(new_n658_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n730_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n734_));
  OAI21_X1  g533(.A(KEYINPUT108), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n736_), .B(KEYINPUT43), .C1(new_n659_), .C2(new_n730_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n327_), .A2(KEYINPUT37), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(new_n328_), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n612_), .B(new_n446_), .C1(new_n454_), .C2(new_n456_), .ZN(new_n740_));
  AOI22_X1  g539(.A1(new_n740_), .A2(new_n358_), .B1(new_n457_), .B2(new_n627_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n640_), .B1(new_n741_), .B2(new_n613_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n651_), .A2(new_n658_), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n734_), .B(new_n739_), .C1(new_n742_), .C2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT109), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n733_), .A2(new_n746_), .A3(new_n734_), .ZN(new_n747_));
  AOI22_X1  g546(.A1(new_n735_), .A2(new_n737_), .B1(new_n745_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n354_), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n697_), .A2(new_n698_), .A3(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n729_), .B1(new_n748_), .B2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n739_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n736_), .B1(new_n753_), .B2(KEYINPUT43), .ZN(new_n754_));
  INV_X1    g553(.A(new_n737_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n746_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n756_));
  NOR4_X1   g555(.A1(new_n659_), .A2(KEYINPUT109), .A3(new_n730_), .A4(KEYINPUT43), .ZN(new_n757_));
  OAI22_X1  g556(.A1(new_n754_), .A2(new_n755_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(KEYINPUT44), .A3(new_n750_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n752_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n619_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(G29gat), .ZN(new_n762_));
  INV_X1    g561(.A(new_n327_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n763_), .A2(new_n749_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n293_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n690_), .A2(new_n765_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n642_), .A2(G29gat), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n767_), .B(KEYINPUT110), .Z(new_n768_));
  OAI21_X1  g567(.A(new_n762_), .B1(new_n766_), .B2(new_n768_), .ZN(G1328gat));
  NOR2_X1   g568(.A1(new_n705_), .A2(G36gat), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n690_), .A2(new_n765_), .A3(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT45), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n752_), .A2(new_n704_), .A3(new_n759_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(G36gat), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT46), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n772_), .A2(new_n774_), .A3(KEYINPUT46), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(G1329gat));
  NOR2_X1   g578(.A1(new_n641_), .A2(new_n637_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n752_), .A2(new_n759_), .A3(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT111), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n752_), .A2(new_n759_), .A3(KEYINPUT111), .A4(new_n780_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n637_), .B1(new_n766_), .B2(new_n641_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n783_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT47), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT47), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n783_), .A2(new_n788_), .A3(new_n784_), .A4(new_n785_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(G1330gat));
  INV_X1    g589(.A(G50gat), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n656_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n690_), .A2(new_n721_), .A3(new_n765_), .ZN(new_n793_));
  AOI22_X1  g592(.A1(new_n760_), .A2(new_n792_), .B1(new_n791_), .B2(new_n793_), .ZN(G1331gat));
  NOR3_X1   g593(.A1(new_n293_), .A2(new_n659_), .A3(new_n687_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n355_), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n796_), .B(KEYINPUT112), .Z(new_n797_));
  INV_X1    g596(.A(G57gat), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(new_n798_), .A3(new_n619_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n697_), .A2(new_n688_), .A3(new_n749_), .A4(new_n700_), .ZN(new_n800_));
  OAI21_X1  g599(.A(G57gat), .B1(new_n800_), .B2(new_n642_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(G1332gat));
  INV_X1    g601(.A(G64gat), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n797_), .A2(new_n803_), .A3(new_n704_), .ZN(new_n804_));
  OAI21_X1  g603(.A(G64gat), .B1(new_n800_), .B2(new_n705_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(KEYINPUT48), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(G1333gat));
  INV_X1    g606(.A(G71gat), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n797_), .A2(new_n808_), .A3(new_n640_), .ZN(new_n809_));
  OAI21_X1  g608(.A(G71gat), .B1(new_n800_), .B2(new_n641_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(KEYINPUT49), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(G1334gat));
  INV_X1    g611(.A(G78gat), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n797_), .A2(new_n813_), .A3(new_n721_), .ZN(new_n814_));
  OAI21_X1  g613(.A(G78gat), .B1(new_n800_), .B2(new_n720_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(KEYINPUT50), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n816_), .ZN(G1335gat));
  NAND2_X1  g616(.A1(new_n795_), .A2(new_n764_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(G85gat), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n820_), .A3(new_n619_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n293_), .A2(new_n687_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n354_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n822_), .B1(new_n748_), .B2(new_n824_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n758_), .A2(KEYINPUT113), .A3(new_n354_), .A4(new_n823_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n642_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n821_), .B1(new_n827_), .B2(new_n820_), .ZN(G1336gat));
  AOI21_X1  g627(.A(G92gat), .B1(new_n819_), .B2(new_n704_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n825_), .A2(new_n826_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n704_), .A2(new_n232_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n829_), .B1(new_n830_), .B2(new_n831_), .ZN(G1337gat));
  AND4_X1   g631(.A1(new_n640_), .A2(new_n795_), .A3(new_n229_), .A4(new_n764_), .ZN(new_n833_));
  XOR2_X1   g632(.A(new_n833_), .B(KEYINPUT114), .Z(new_n834_));
  INV_X1    g633(.A(G99gat), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n641_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n834_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT51), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT51), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n834_), .B(new_n839_), .C1(new_n835_), .C2(new_n836_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(G1338gat));
  XNOR2_X1  g640(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n748_), .A2(new_n656_), .A3(new_n824_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT52), .B1(new_n843_), .B2(new_n230_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n758_), .A2(new_n457_), .A3(new_n354_), .A4(new_n823_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n846_), .A3(G106gat), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n844_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n457_), .A2(new_n230_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n818_), .A2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n842_), .B1(new_n848_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n842_), .ZN(new_n853_));
  AOI211_X1 g652(.A(new_n850_), .B(new_n853_), .C1(new_n844_), .C2(new_n847_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n852_), .A2(new_n854_), .ZN(G1339gat));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n250_), .A2(new_n254_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n247_), .B1(new_n222_), .B2(new_n240_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n266_), .A2(KEYINPUT72), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n270_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n258_), .B1(new_n857_), .B2(new_n860_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n267_), .A2(new_n268_), .A3(KEYINPUT55), .A4(new_n270_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT55), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n248_), .A2(new_n257_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n860_), .B2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n861_), .A2(new_n862_), .A3(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n275_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT56), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n866_), .A2(KEYINPUT56), .A3(new_n275_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  AOI22_X1  g670(.A1(new_n685_), .A2(new_n686_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n673_), .B1(new_n669_), .B2(new_n663_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(new_n663_), .B2(new_n662_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n679_), .A2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT116), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n679_), .A2(new_n877_), .A3(new_n874_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n871_), .A2(new_n872_), .B1(new_n284_), .B2(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n856_), .B1(new_n880_), .B2(new_n327_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n871_), .A2(new_n872_), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n284_), .A2(new_n879_), .ZN(new_n883_));
  OAI211_X1 g682(.A(KEYINPUT57), .B(new_n763_), .C1(new_n882_), .C2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n879_), .A2(new_n281_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(KEYINPUT117), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT117), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n879_), .A2(new_n281_), .A3(new_n887_), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n886_), .A2(KEYINPUT58), .A3(new_n888_), .A4(new_n871_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n739_), .ZN(new_n890_));
  AOI22_X1  g689(.A1(new_n878_), .A2(new_n876_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n891_));
  AOI22_X1  g690(.A1(new_n891_), .A2(new_n887_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n892_));
  AOI21_X1  g691(.A(KEYINPUT58), .B1(new_n892_), .B2(new_n886_), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n881_), .B(new_n884_), .C1(new_n890_), .C2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT118), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT58), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n888_), .A2(new_n871_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n891_), .A2(new_n887_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n897_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n900_), .A2(new_n739_), .A3(new_n889_), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n901_), .A2(KEYINPUT118), .A3(new_n881_), .A4(new_n884_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n896_), .A2(new_n354_), .A3(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT54), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n355_), .A2(new_n904_), .A3(new_n289_), .A4(new_n688_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n688_), .A2(new_n287_), .A3(new_n286_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n738_), .A2(new_n749_), .A3(new_n328_), .ZN(new_n907_));
  OAI21_X1  g706(.A(KEYINPUT54), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n905_), .A2(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n903_), .A2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT119), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n903_), .A2(KEYINPUT119), .A3(new_n909_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n704_), .A2(new_n642_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(new_n650_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n912_), .A2(new_n913_), .A3(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(G113gat), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n918_), .A2(new_n919_), .A3(new_n687_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n894_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n909_), .B1(new_n921_), .B2(new_n749_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n923_));
  AND3_X1   g722(.A1(new_n922_), .A2(new_n916_), .A3(new_n923_), .ZN(new_n924_));
  AOI211_X1 g723(.A(new_n688_), .B(new_n924_), .C1(new_n917_), .C2(KEYINPUT59), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n920_), .B1(new_n925_), .B2(new_n919_), .ZN(G1340gat));
  AOI211_X1 g725(.A(new_n293_), .B(new_n924_), .C1(new_n917_), .C2(KEYINPUT59), .ZN(new_n927_));
  INV_X1    g726(.A(G120gat), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n928_), .B1(new_n293_), .B2(KEYINPUT60), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n929_), .B1(KEYINPUT60), .B2(new_n928_), .ZN(new_n930_));
  OAI22_X1  g729(.A1(new_n927_), .A2(new_n928_), .B1(new_n917_), .B2(new_n930_), .ZN(G1341gat));
  INV_X1    g730(.A(G127gat), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n918_), .A2(new_n932_), .A3(new_n749_), .ZN(new_n933_));
  AOI211_X1 g732(.A(new_n354_), .B(new_n924_), .C1(new_n917_), .C2(KEYINPUT59), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n933_), .B1(new_n934_), .B2(new_n932_), .ZN(G1342gat));
  AOI21_X1  g734(.A(G134gat), .B1(new_n918_), .B2(new_n327_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n924_), .B1(new_n917_), .B2(KEYINPUT59), .ZN(new_n937_));
  XOR2_X1   g736(.A(KEYINPUT121), .B(G134gat), .Z(new_n938_));
  NOR2_X1   g737(.A1(new_n730_), .A2(new_n938_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n936_), .B1(new_n937_), .B2(new_n939_), .ZN(G1343gat));
  INV_X1    g739(.A(new_n909_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n749_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n942_));
  AOI211_X1 g741(.A(new_n911_), .B(new_n941_), .C1(new_n942_), .C2(new_n902_), .ZN(new_n943_));
  AOI21_X1  g742(.A(KEYINPUT119), .B1(new_n903_), .B2(new_n909_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n943_), .A2(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n457_), .A2(new_n641_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n915_), .A2(new_n946_), .ZN(new_n947_));
  XOR2_X1   g746(.A(new_n947_), .B(KEYINPUT122), .Z(new_n948_));
  NAND2_X1  g747(.A1(new_n945_), .A2(new_n948_), .ZN(new_n949_));
  INV_X1    g748(.A(new_n949_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n950_), .A2(new_n376_), .A3(new_n687_), .ZN(new_n951_));
  OAI21_X1  g750(.A(G141gat), .B1(new_n949_), .B2(new_n698_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n951_), .A2(new_n952_), .ZN(G1344gat));
  NAND3_X1  g752(.A1(new_n950_), .A2(new_n377_), .A3(new_n697_), .ZN(new_n954_));
  OAI21_X1  g753(.A(G148gat), .B1(new_n949_), .B2(new_n293_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n954_), .A2(new_n955_), .ZN(G1345gat));
  NAND4_X1  g755(.A1(new_n912_), .A2(new_n749_), .A3(new_n913_), .A4(new_n948_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n957_), .A2(KEYINPUT123), .ZN(new_n958_));
  INV_X1    g757(.A(KEYINPUT123), .ZN(new_n959_));
  NAND4_X1  g758(.A1(new_n945_), .A2(new_n959_), .A3(new_n749_), .A4(new_n948_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(KEYINPUT61), .B(G155gat), .ZN(new_n961_));
  AND3_X1   g760(.A1(new_n958_), .A2(new_n960_), .A3(new_n961_), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n961_), .B1(new_n958_), .B2(new_n960_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n962_), .A2(new_n963_), .ZN(G1346gat));
  OR3_X1    g763(.A1(new_n949_), .A2(G162gat), .A3(new_n763_), .ZN(new_n965_));
  OAI21_X1  g764(.A(G162gat), .B1(new_n949_), .B2(new_n730_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n965_), .A2(new_n966_), .ZN(G1347gat));
  NAND2_X1  g766(.A1(new_n704_), .A2(new_n642_), .ZN(new_n968_));
  NOR2_X1   g767(.A1(new_n968_), .A2(new_n641_), .ZN(new_n969_));
  INV_X1    g768(.A(new_n969_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(new_n721_), .A2(new_n970_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n922_), .A2(new_n971_), .ZN(new_n972_));
  INV_X1    g771(.A(new_n972_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n973_), .A2(new_n687_), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n974_), .A2(G169gat), .ZN(new_n975_));
  INV_X1    g774(.A(KEYINPUT124), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n975_), .A2(new_n976_), .ZN(new_n977_));
  NAND3_X1  g776(.A1(new_n974_), .A2(KEYINPUT124), .A3(G169gat), .ZN(new_n978_));
  NAND3_X1  g777(.A1(new_n977_), .A2(KEYINPUT62), .A3(new_n978_), .ZN(new_n979_));
  INV_X1    g778(.A(KEYINPUT62), .ZN(new_n980_));
  NAND3_X1  g779(.A1(new_n975_), .A2(new_n976_), .A3(new_n980_), .ZN(new_n981_));
  NAND3_X1  g780(.A1(new_n973_), .A2(new_n511_), .A3(new_n687_), .ZN(new_n982_));
  NAND3_X1  g781(.A1(new_n979_), .A2(new_n981_), .A3(new_n982_), .ZN(G1348gat));
  AOI21_X1  g782(.A(G176gat), .B1(new_n973_), .B2(new_n697_), .ZN(new_n984_));
  NAND3_X1  g783(.A1(new_n912_), .A2(new_n656_), .A3(new_n913_), .ZN(new_n985_));
  INV_X1    g784(.A(KEYINPUT125), .ZN(new_n986_));
  XNOR2_X1  g785(.A(new_n985_), .B(new_n986_), .ZN(new_n987_));
  NOR3_X1   g786(.A1(new_n293_), .A2(new_n512_), .A3(new_n970_), .ZN(new_n988_));
  AOI21_X1  g787(.A(new_n984_), .B1(new_n987_), .B2(new_n988_), .ZN(G1349gat));
  OR3_X1    g788(.A1(new_n972_), .A2(new_n521_), .A3(new_n354_), .ZN(new_n990_));
  XNOR2_X1  g789(.A(new_n990_), .B(KEYINPUT126), .ZN(new_n991_));
  NOR2_X1   g790(.A1(new_n970_), .A2(new_n354_), .ZN(new_n992_));
  AOI21_X1  g791(.A(KEYINPUT125), .B1(new_n945_), .B2(new_n656_), .ZN(new_n993_));
  NOR4_X1   g792(.A1(new_n943_), .A2(new_n944_), .A3(new_n986_), .A4(new_n457_), .ZN(new_n994_));
  OAI21_X1  g793(.A(new_n992_), .B1(new_n993_), .B2(new_n994_), .ZN(new_n995_));
  AOI21_X1  g794(.A(new_n991_), .B1(new_n995_), .B2(new_n545_), .ZN(G1350gat));
  OAI21_X1  g795(.A(G190gat), .B1(new_n972_), .B2(new_n730_), .ZN(new_n997_));
  NAND2_X1  g796(.A1(new_n327_), .A2(new_n520_), .ZN(new_n998_));
  OAI21_X1  g797(.A(new_n997_), .B1(new_n972_), .B2(new_n998_), .ZN(G1351gat));
  NOR2_X1   g798(.A1(new_n968_), .A2(new_n946_), .ZN(new_n1000_));
  NAND3_X1  g799(.A1(new_n945_), .A2(new_n687_), .A3(new_n1000_), .ZN(new_n1001_));
  XNOR2_X1  g800(.A(new_n1001_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g801(.A1(new_n912_), .A2(new_n913_), .ZN(new_n1003_));
  INV_X1    g802(.A(new_n1000_), .ZN(new_n1004_));
  NOR2_X1   g803(.A1(new_n1003_), .A2(new_n1004_), .ZN(new_n1005_));
  NAND2_X1  g804(.A1(new_n1005_), .A2(new_n697_), .ZN(new_n1006_));
  OAI21_X1  g805(.A(new_n1006_), .B1(KEYINPUT127), .B2(G204gat), .ZN(new_n1007_));
  XNOR2_X1  g806(.A(KEYINPUT127), .B(G204gat), .ZN(new_n1008_));
  NAND3_X1  g807(.A1(new_n1005_), .A2(new_n697_), .A3(new_n1008_), .ZN(new_n1009_));
  NAND2_X1  g808(.A1(new_n1007_), .A2(new_n1009_), .ZN(G1353gat));
  NAND2_X1  g809(.A1(new_n1005_), .A2(new_n749_), .ZN(new_n1011_));
  OAI21_X1  g810(.A(new_n1011_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n1012_));
  XNOR2_X1  g811(.A(KEYINPUT63), .B(G211gat), .ZN(new_n1013_));
  NAND3_X1  g812(.A1(new_n1005_), .A2(new_n749_), .A3(new_n1013_), .ZN(new_n1014_));
  NAND2_X1  g813(.A1(new_n1012_), .A2(new_n1014_), .ZN(G1354gat));
  NAND3_X1  g814(.A1(new_n1005_), .A2(new_n410_), .A3(new_n327_), .ZN(new_n1016_));
  NOR3_X1   g815(.A1(new_n1003_), .A2(new_n730_), .A3(new_n1004_), .ZN(new_n1017_));
  OAI21_X1  g816(.A(new_n1016_), .B1(new_n410_), .B2(new_n1017_), .ZN(G1355gat));
endmodule


