//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G113gat), .B(G120gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(G71gat), .B(G99gat), .Z(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(G43gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT30), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n207_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G227gat), .A2(G233gat), .ZN(new_n211_));
  INV_X1    g010(.A(G15gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n210_), .B(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT25), .B(G183gat), .ZN(new_n215_));
  INV_X1    g014(.A(G190gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT26), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT82), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n216_), .A2(KEYINPUT26), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n216_), .A2(KEYINPUT82), .A3(KEYINPUT26), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n215_), .A2(new_n219_), .A3(new_n220_), .A4(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223_));
  INV_X1    g022(.A(G169gat), .ZN(new_n224_));
  INV_X1    g023(.A(G176gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT23), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT23), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(G183gat), .A3(G190gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n224_), .A2(new_n225_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(KEYINPUT24), .A3(new_n233_), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n222_), .A2(new_n226_), .A3(new_n231_), .A4(new_n234_), .ZN(new_n235_));
  OR2_X1    g034(.A1(KEYINPUT86), .A2(G176gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(KEYINPUT86), .A2(G176gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT85), .ZN(new_n238_));
  OAI21_X1  g037(.A(G169gat), .B1(new_n238_), .B2(KEYINPUT22), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT22), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n240_), .A2(KEYINPUT85), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n236_), .B(new_n237_), .C1(new_n239_), .C2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT83), .B(G169gat), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT84), .B1(new_n243_), .B2(new_n240_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT84), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT83), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n246_), .A2(G169gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n224_), .A2(KEYINPUT83), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n245_), .B(KEYINPUT22), .C1(new_n247_), .C2(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n242_), .B1(new_n244_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT87), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n228_), .A2(new_n230_), .A3(new_n251_), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n229_), .A2(KEYINPUT87), .A3(G183gat), .A4(G190gat), .ZN(new_n253_));
  OR2_X1    g052(.A1(G183gat), .A2(G190gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n233_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n235_), .B1(new_n250_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(KEYINPUT88), .B1(new_n214_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT31), .ZN(new_n260_));
  INV_X1    g059(.A(new_n213_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n210_), .B(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(new_n257_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n259_), .A2(new_n260_), .A3(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n260_), .B1(new_n259_), .B2(new_n263_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n204_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n266_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n204_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(new_n269_), .A3(new_n264_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G225gat), .A2(G233gat), .ZN(new_n271_));
  XOR2_X1   g070(.A(new_n271_), .B(KEYINPUT98), .Z(new_n272_));
  XNOR2_X1  g071(.A(G155gat), .B(G162gat), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(G141gat), .A2(G148gat), .ZN(new_n275_));
  NOR2_X1   g074(.A1(KEYINPUT89), .A2(KEYINPUT3), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G141gat), .A2(G148gat), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT90), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT2), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n278_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  OAI22_X1  g080(.A1(KEYINPUT89), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n277_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n280_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n274_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(G141gat), .B(G148gat), .Z(new_n286_));
  NAND3_X1  g085(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n286_), .B(new_n287_), .C1(KEYINPUT1), .C2(new_n273_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n285_), .A2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n269_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(KEYINPUT91), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT91), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n285_), .A2(new_n293_), .A3(new_n288_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n292_), .A2(new_n294_), .A3(new_n269_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n291_), .A2(KEYINPUT4), .A3(new_n295_), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n285_), .A2(new_n293_), .A3(new_n288_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n293_), .B1(new_n285_), .B2(new_n288_), .ZN(new_n298_));
  NOR3_X1   g097(.A1(new_n297_), .A2(new_n298_), .A3(new_n204_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT4), .ZN(new_n300_));
  AOI21_X1  g099(.A(KEYINPUT99), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n292_), .A2(new_n300_), .A3(new_n294_), .A4(new_n269_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT99), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n272_), .B(new_n296_), .C1(new_n301_), .C2(new_n304_), .ZN(new_n305_));
  NOR3_X1   g104(.A1(new_n299_), .A2(new_n290_), .A3(new_n272_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G1gat), .B(G29gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G57gat), .B(G85gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT100), .B(KEYINPUT0), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n308_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n313_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n305_), .A2(new_n307_), .A3(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n267_), .A2(new_n270_), .A3(new_n318_), .ZN(new_n319_));
  XOR2_X1   g118(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n320_));
  NOR2_X1   g119(.A1(new_n297_), .A2(new_n298_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n320_), .B1(new_n321_), .B2(KEYINPUT29), .ZN(new_n322_));
  XOR2_X1   g121(.A(G22gat), .B(G50gat), .Z(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n292_), .A2(new_n294_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT29), .ZN(new_n326_));
  INV_X1    g125(.A(new_n320_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n325_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n322_), .A2(new_n324_), .A3(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n324_), .B1(new_n322_), .B2(new_n328_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  XOR2_X1   g130(.A(G78gat), .B(G106gat), .Z(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  XOR2_X1   g132(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n334_));
  AOI21_X1  g133(.A(new_n334_), .B1(new_n285_), .B2(new_n288_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT94), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  OR2_X1    g136(.A1(G197gat), .A2(G204gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G197gat), .A2(G204gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n338_), .A2(KEYINPUT21), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT21), .ZN(new_n341_));
  AND2_X1   g140(.A1(G197gat), .A2(G204gat), .ZN(new_n342_));
  NOR2_X1   g141(.A1(G197gat), .A2(G204gat), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n341_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G211gat), .B(G218gat), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n340_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(G218gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(G211gat), .ZN(new_n348_));
  INV_X1    g147(.A(G211gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(G218gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n351_), .A2(KEYINPUT21), .A3(new_n338_), .A4(new_n339_), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n346_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n354_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n355_));
  OAI211_X1 g154(.A(G228gat), .B(G233gat), .C1(new_n337_), .C2(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n353_), .B1(G228gat), .B2(G233gat), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n357_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n333_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n356_), .A2(new_n333_), .A3(new_n358_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n331_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n361_), .ZN(new_n363_));
  OAI22_X1  g162(.A1(new_n363_), .A2(new_n359_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G226gat), .A2(G233gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT19), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n353_), .B(new_n235_), .C1(new_n250_), .C2(new_n256_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT20), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n252_), .A2(new_n226_), .A3(new_n253_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT95), .ZN(new_n372_));
  INV_X1    g171(.A(new_n234_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n220_), .A2(new_n217_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n373_), .B1(new_n374_), .B2(new_n215_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT95), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n252_), .A2(new_n376_), .A3(new_n226_), .A4(new_n253_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n372_), .A2(new_n375_), .A3(new_n377_), .ZN(new_n378_));
  AOI22_X1  g177(.A1(new_n231_), .A2(new_n254_), .B1(G169gat), .B2(G176gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT22), .B(G169gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT96), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n236_), .A2(new_n237_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n379_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n353_), .B1(new_n378_), .B2(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n368_), .B1(new_n370_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n257_), .A2(new_n354_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n378_), .A2(new_n383_), .A3(new_n353_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n368_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n386_), .A2(new_n387_), .A3(KEYINPUT20), .A4(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n385_), .A2(new_n389_), .ZN(new_n390_));
  XOR2_X1   g189(.A(G8gat), .B(G36gat), .Z(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT18), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G64gat), .B(G92gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n390_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT97), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n385_), .A2(new_n394_), .A3(new_n389_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n396_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n385_), .A2(KEYINPUT97), .A3(new_n389_), .A4(new_n394_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT27), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n386_), .A2(new_n387_), .A3(KEYINPUT20), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(new_n368_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n378_), .A2(new_n383_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n354_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n406_), .A2(KEYINPUT20), .A3(new_n388_), .A4(new_n369_), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n404_), .A2(new_n407_), .ZN(new_n408_));
  OAI211_X1 g207(.A(KEYINPUT27), .B(new_n398_), .C1(new_n408_), .C2(new_n394_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n402_), .A2(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n366_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n319_), .A2(new_n411_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n362_), .A2(new_n314_), .A3(new_n364_), .A4(new_n316_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT101), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n385_), .A2(new_n415_), .A3(new_n389_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n394_), .A2(KEYINPUT32), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n404_), .A2(new_n407_), .A3(KEYINPUT32), .A4(new_n394_), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n385_), .A2(KEYINPUT101), .A3(new_n389_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n418_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n272_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n290_), .B1(new_n321_), .B2(new_n269_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n422_), .B1(new_n423_), .B2(KEYINPUT4), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n299_), .A2(KEYINPUT99), .A3(new_n300_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n302_), .A2(new_n303_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  AOI211_X1 g226(.A(new_n306_), .B(new_n313_), .C1(new_n424_), .C2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n315_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n421_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT102), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n291_), .A2(new_n295_), .A3(new_n272_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n313_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n272_), .B1(new_n423_), .B2(KEYINPUT4), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n433_), .B1(new_n434_), .B2(new_n427_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT33), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n435_), .B1(new_n316_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n399_), .A2(new_n400_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n305_), .A2(KEYINPUT33), .A3(new_n307_), .A4(new_n315_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT102), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n421_), .B(new_n441_), .C1(new_n428_), .C2(new_n429_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n431_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n414_), .B1(new_n443_), .B2(new_n365_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n267_), .A2(new_n270_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n412_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G1gat), .B(G8gat), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT14), .ZN(new_n449_));
  XOR2_X1   g248(.A(KEYINPUT76), .B(G8gat), .Z(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT75), .B(G1gat), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n449_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  XOR2_X1   g251(.A(G15gat), .B(G22gat), .Z(new_n453_));
  NOR3_X1   g252(.A1(new_n452_), .A2(KEYINPUT77), .A3(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT77), .ZN(new_n455_));
  XOR2_X1   g254(.A(KEYINPUT75), .B(G1gat), .Z(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT76), .B(G8gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT14), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n453_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n455_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n448_), .B1(new_n454_), .B2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT77), .B1(new_n452_), .B2(new_n453_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n458_), .A2(new_n455_), .A3(new_n459_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(new_n463_), .A3(new_n447_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G29gat), .B(G36gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G43gat), .B(G50gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n461_), .A2(new_n464_), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT79), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT79), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n461_), .A2(new_n470_), .A3(new_n464_), .A4(new_n467_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n461_), .A2(new_n464_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n467_), .ZN(new_n473_));
  AOI22_X1  g272(.A1(new_n469_), .A2(new_n471_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G229gat), .A2(G233gat), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT80), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n469_), .A2(new_n471_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n475_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n467_), .B(KEYINPUT15), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n479_), .B1(new_n472_), .B2(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n477_), .B1(new_n478_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n478_), .A2(new_n477_), .A3(new_n481_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n476_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G113gat), .B(G141gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G169gat), .B(G197gat), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n486_), .B(new_n487_), .Z(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT81), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n485_), .A2(new_n491_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n476_), .A2(new_n483_), .A3(new_n490_), .A4(new_n484_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n446_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT103), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G230gat), .A2(G233gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT64), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G85gat), .B(G92gat), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT9), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(KEYINPUT10), .B(G99gat), .Z(new_n502_));
  INV_X1    g301(.A(G106gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G99gat), .A2(G106gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT6), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n500_), .A2(G85gat), .A3(G92gat), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n501_), .A2(new_n504_), .A3(new_n506_), .A4(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n499_), .B(KEYINPUT66), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT8), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT65), .ZN(new_n511_));
  OR4_X1    g310(.A1(new_n511_), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n512_));
  OAI22_X1  g311(.A1(new_n511_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n506_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n509_), .A2(new_n510_), .A3(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n510_), .B1(new_n509_), .B2(new_n514_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n508_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G57gat), .B(G64gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT11), .ZN(new_n519_));
  XOR2_X1   g318(.A(G71gat), .B(G78gat), .Z(new_n520_));
  OR2_X1    g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n518_), .A2(KEYINPUT11), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n519_), .A2(new_n520_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n521_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT67), .B1(new_n517_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n508_), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n506_), .A2(new_n513_), .A3(new_n512_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT66), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n499_), .B(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(KEYINPUT8), .B1(new_n528_), .B2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n509_), .A2(new_n510_), .A3(new_n514_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n527_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(new_n524_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n498_), .B1(new_n526_), .B2(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n535_), .B1(new_n534_), .B2(new_n526_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT68), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n517_), .A2(new_n525_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n498_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n537_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT12), .B1(new_n533_), .B2(new_n524_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT12), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n517_), .A2(new_n542_), .A3(new_n525_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n534_), .A2(KEYINPUT68), .A3(new_n498_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n540_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n536_), .A2(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(G120gat), .B(G148gat), .Z(new_n548_));
  XNOR2_X1  g347(.A(G176gat), .B(G204gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n550_), .B(new_n551_), .Z(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n547_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n536_), .A2(new_n546_), .A3(new_n552_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT13), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n554_), .B(new_n555_), .C1(KEYINPUT70), .C2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT37), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G190gat), .B(G218gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT73), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT74), .ZN(new_n566_));
  XOR2_X1   g365(.A(G134gat), .B(G162gat), .Z(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT36), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n568_), .A2(new_n569_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT71), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT15), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n467_), .B(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n573_), .B1(new_n533_), .B2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n517_), .A2(KEYINPUT71), .A3(new_n480_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT72), .ZN(new_n579_));
  AOI211_X1 g378(.A(new_n473_), .B(new_n527_), .C1(new_n531_), .C2(new_n532_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n578_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT34), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT35), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n579_), .A2(new_n582_), .A3(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n580_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n585_), .A2(new_n586_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT72), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n591_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n587_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n589_), .B(new_n590_), .C1(new_n592_), .C2(new_n593_), .ZN(new_n594_));
  AOI211_X1 g393(.A(new_n571_), .B(new_n572_), .C1(new_n588_), .C2(new_n594_), .ZN(new_n595_));
  AND4_X1   g394(.A1(new_n569_), .A2(new_n588_), .A3(new_n594_), .A4(new_n568_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n563_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n572_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n593_), .B1(new_n578_), .B2(KEYINPUT72), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n578_), .A2(new_n581_), .A3(new_n590_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NOR3_X1   g400(.A1(new_n592_), .A2(new_n589_), .A3(new_n593_), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n570_), .B(new_n598_), .C1(new_n601_), .C2(new_n602_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n588_), .A2(new_n594_), .A3(new_n569_), .A4(new_n568_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n603_), .A2(KEYINPUT37), .A3(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n597_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(G231gat), .A2(G233gat), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n524_), .B(new_n607_), .Z(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(new_n472_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G127gat), .B(G155gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G183gat), .B(G211gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT17), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n609_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n609_), .A2(KEYINPUT17), .A3(new_n614_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n606_), .A2(new_n619_), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n496_), .A2(new_n562_), .A3(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(new_n317_), .A3(new_n456_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT38), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n595_), .A2(new_n596_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n446_), .A2(new_n626_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n562_), .A2(KEYINPUT104), .A3(new_n494_), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT104), .B1(new_n562_), .B2(new_n494_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n628_), .A2(new_n629_), .A3(new_n619_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n627_), .A2(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G1gat), .B1(new_n631_), .B2(new_n318_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n622_), .A2(new_n623_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n624_), .A2(new_n632_), .A3(new_n633_), .ZN(G1324gat));
  INV_X1    g433(.A(KEYINPUT40), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n627_), .A2(new_n630_), .A3(new_n410_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT105), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(G8gat), .B1(new_n636_), .B2(new_n637_), .ZN(new_n639_));
  OR3_X1    g438(.A1(new_n638_), .A2(new_n639_), .A3(KEYINPUT106), .ZN(new_n640_));
  OAI21_X1  g439(.A(KEYINPUT106), .B1(new_n638_), .B2(new_n639_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n640_), .A2(KEYINPUT39), .A3(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n621_), .A2(new_n410_), .A3(new_n457_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n643_), .B1(KEYINPUT39), .B2(new_n641_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n635_), .B1(new_n642_), .B2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n640_), .A2(KEYINPUT39), .A3(new_n641_), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n641_), .A2(KEYINPUT39), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n646_), .A2(KEYINPUT40), .A3(new_n647_), .A4(new_n643_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n645_), .A2(new_n648_), .ZN(G1325gat));
  NAND3_X1  g448(.A1(new_n621_), .A2(new_n212_), .A3(new_n445_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n631_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(new_n445_), .ZN(new_n652_));
  AOI21_X1  g451(.A(KEYINPUT41), .B1(new_n652_), .B2(G15gat), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n652_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n650_), .B1(new_n653_), .B2(new_n654_), .ZN(G1326gat));
  INV_X1    g454(.A(G22gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n621_), .A2(new_n656_), .A3(new_n366_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G22gat), .B1(new_n631_), .B2(new_n365_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n658_), .A2(KEYINPUT42), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n658_), .A2(KEYINPUT42), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n657_), .B1(new_n659_), .B2(new_n660_), .ZN(G1327gat));
  INV_X1    g460(.A(new_n562_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n662_), .A2(new_n618_), .A3(new_n626_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n496_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(G29gat), .B1(new_n665_), .B2(new_n317_), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n603_), .A2(KEYINPUT37), .A3(new_n604_), .ZN(new_n667_));
  AOI21_X1  g466(.A(KEYINPUT37), .B1(new_n603_), .B2(new_n604_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT107), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n667_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT107), .B1(new_n597_), .B2(new_n605_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n446_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n606_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n674_), .A2(KEYINPUT43), .ZN(new_n675_));
  AOI22_X1  g474(.A1(new_n673_), .A2(KEYINPUT43), .B1(new_n446_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n628_), .A2(new_n629_), .A3(new_n618_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n677_), .A2(KEYINPUT44), .A3(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n678_), .ZN(new_n681_));
  OAI21_X1  g480(.A(KEYINPUT108), .B1(new_n676_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT108), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n446_), .A2(new_n675_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n446_), .B2(new_n672_), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n684_), .B(new_n678_), .C1(new_n685_), .C2(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n682_), .A2(new_n683_), .A3(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(KEYINPUT109), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n678_), .B1(new_n685_), .B2(new_n687_), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT44), .B1(new_n691_), .B2(KEYINPUT108), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT109), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(new_n693_), .A3(new_n688_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n680_), .B1(new_n690_), .B2(new_n694_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n317_), .A2(G29gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n666_), .B1(new_n695_), .B2(new_n696_), .ZN(G1328gat));
  INV_X1    g496(.A(new_n410_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n698_), .A2(G36gat), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  OR3_X1    g499(.A1(new_n664_), .A2(KEYINPUT45), .A3(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(KEYINPUT45), .B1(new_n664_), .B2(new_n700_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n679_), .A2(new_n410_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n704_), .B1(new_n690_), .B2(new_n694_), .ZN(new_n705_));
  INV_X1    g504(.A(G36gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n703_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT46), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  OAI211_X1 g508(.A(KEYINPUT46), .B(new_n703_), .C1(new_n705_), .C2(new_n706_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1329gat));
  AND2_X1   g510(.A1(new_n445_), .A2(G43gat), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n689_), .A2(KEYINPUT109), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n693_), .B1(new_n692_), .B2(new_n688_), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n679_), .B(new_n712_), .C1(new_n713_), .C2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n665_), .A2(new_n445_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(KEYINPUT110), .B(G43gat), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n715_), .A2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n715_), .A2(new_n718_), .A3(new_n720_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1330gat));
  AOI21_X1  g523(.A(G50gat), .B1(new_n665_), .B2(new_n366_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n366_), .A2(G50gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n695_), .B2(new_n726_), .ZN(G1331gat));
  INV_X1    g526(.A(new_n494_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n446_), .A2(new_n728_), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n729_), .A2(new_n662_), .A3(new_n620_), .ZN(new_n730_));
  INV_X1    g529(.A(G57gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n731_), .A3(new_n317_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n492_), .A2(new_n618_), .A3(new_n493_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n562_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n627_), .A2(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(G57gat), .B1(new_n735_), .B2(new_n318_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n732_), .A2(new_n736_), .ZN(G1332gat));
  OAI21_X1  g536(.A(G64gat), .B1(new_n735_), .B2(new_n698_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT48), .ZN(new_n739_));
  INV_X1    g538(.A(G64gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n730_), .A2(new_n740_), .A3(new_n410_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(G1333gat));
  INV_X1    g541(.A(G71gat), .ZN(new_n743_));
  INV_X1    g542(.A(new_n735_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n744_), .B2(new_n445_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT49), .Z(new_n746_));
  NAND3_X1  g545(.A1(new_n730_), .A2(new_n743_), .A3(new_n445_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1334gat));
  OAI21_X1  g547(.A(G78gat), .B1(new_n735_), .B2(new_n365_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT50), .ZN(new_n750_));
  INV_X1    g549(.A(G78gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n730_), .A2(new_n751_), .A3(new_n366_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1335gat));
  NOR3_X1   g552(.A1(new_n562_), .A2(new_n626_), .A3(new_n618_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n729_), .A2(new_n754_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT112), .Z(new_n756_));
  AOI21_X1  g555(.A(G85gat), .B1(new_n756_), .B2(new_n317_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT113), .ZN(new_n758_));
  NOR4_X1   g557(.A1(new_n676_), .A2(new_n494_), .A3(new_n562_), .A4(new_n618_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n759_), .A2(G85gat), .A3(new_n317_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n758_), .A2(new_n761_), .ZN(G1336gat));
  INV_X1    g561(.A(G92gat), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n756_), .A2(new_n763_), .A3(new_n410_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n759_), .A2(new_n410_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n764_), .B1(new_n766_), .B2(new_n763_), .ZN(G1337gat));
  NAND3_X1  g566(.A1(new_n756_), .A2(new_n445_), .A3(new_n502_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n759_), .A2(new_n445_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(G99gat), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g571(.A1(new_n756_), .A2(new_n503_), .A3(new_n366_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n759_), .A2(new_n366_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(G106gat), .ZN(new_n776_));
  AOI211_X1 g575(.A(KEYINPUT52), .B(new_n503_), .C1(new_n759_), .C2(new_n366_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n773_), .B(new_n779_), .C1(new_n776_), .C2(new_n777_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(G1339gat));
  INV_X1    g582(.A(KEYINPUT59), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n733_), .B(KEYINPUT115), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n562_), .A2(new_n605_), .A3(new_n597_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n785_), .A2(KEYINPUT54), .A3(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n662_), .A2(new_n606_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT115), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n733_), .B(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n788_), .B1(new_n789_), .B2(new_n791_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n787_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n546_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n544_), .A2(new_n534_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n797_), .A3(new_n539_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n540_), .A2(KEYINPUT55), .A3(new_n544_), .A4(new_n545_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n538_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT116), .B1(new_n800_), .B2(new_n498_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n795_), .A2(new_n798_), .A3(new_n799_), .A4(new_n801_), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n802_), .A2(KEYINPUT56), .A3(new_n553_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT56), .B1(new_n802_), .B2(new_n553_), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n494_), .B(new_n555_), .C1(new_n803_), .C2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n485_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n489_), .B1(new_n474_), .B2(new_n479_), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n807_), .A2(KEYINPUT117), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n475_), .B1(new_n472_), .B2(new_n480_), .ZN(new_n809_));
  AOI22_X1  g608(.A1(new_n807_), .A2(KEYINPUT117), .B1(new_n478_), .B2(new_n809_), .ZN(new_n810_));
  AOI22_X1  g609(.A1(new_n806_), .A2(new_n488_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n556_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n625_), .B1(new_n805_), .B2(new_n812_), .ZN(new_n813_));
  OR2_X1    g612(.A1(new_n813_), .A2(KEYINPUT57), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(KEYINPUT57), .ZN(new_n815_));
  INV_X1    g614(.A(new_n555_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n804_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n802_), .A2(KEYINPUT56), .A3(new_n553_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n816_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n819_), .A2(KEYINPUT58), .A3(new_n811_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n811_), .B(new_n555_), .C1(new_n804_), .C2(new_n803_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT58), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n820_), .A2(new_n823_), .A3(new_n606_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n814_), .A2(new_n815_), .A3(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n793_), .B1(new_n825_), .B2(new_n619_), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n445_), .A2(new_n317_), .A3(new_n411_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT118), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n784_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n606_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT58), .B1(new_n819_), .B2(new_n811_), .ZN(new_n831_));
  OAI22_X1  g630(.A1(new_n830_), .A2(new_n831_), .B1(new_n813_), .B2(KEYINPUT57), .ZN(new_n832_));
  INV_X1    g631(.A(new_n815_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n619_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  OR2_X1    g633(.A1(new_n787_), .A2(new_n792_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n828_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(KEYINPUT59), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n829_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(G113gat), .B1(new_n840_), .B2(new_n728_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n826_), .A2(new_n828_), .ZN(new_n842_));
  INV_X1    g641(.A(G113gat), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n843_), .A3(new_n494_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n841_), .A2(new_n844_), .ZN(G1340gat));
  INV_X1    g644(.A(KEYINPUT120), .ZN(new_n846_));
  INV_X1    g645(.A(G120gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n562_), .B2(KEYINPUT60), .ZN(new_n848_));
  OR2_X1    g647(.A1(new_n847_), .A2(KEYINPUT60), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n836_), .A2(new_n837_), .A3(new_n848_), .A4(new_n849_), .ZN(new_n850_));
  XOR2_X1   g649(.A(new_n850_), .B(KEYINPUT119), .Z(new_n851_));
  AOI21_X1  g650(.A(new_n847_), .B1(new_n839_), .B2(new_n662_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n846_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n852_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n850_), .B(KEYINPUT119), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n854_), .A2(KEYINPUT120), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n853_), .A2(new_n856_), .ZN(G1341gat));
  OAI21_X1  g656(.A(G127gat), .B1(new_n840_), .B2(new_n619_), .ZN(new_n858_));
  INV_X1    g657(.A(G127gat), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n842_), .A2(new_n859_), .A3(new_n618_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(G1342gat));
  OAI21_X1  g660(.A(G134gat), .B1(new_n840_), .B2(new_n674_), .ZN(new_n862_));
  INV_X1    g661(.A(G134gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n842_), .A2(new_n863_), .A3(new_n625_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(G1343gat));
  NOR4_X1   g664(.A1(new_n445_), .A2(new_n318_), .A3(new_n365_), .A4(new_n410_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n836_), .A2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n494_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n662_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n872_), .B1(new_n867_), .B2(new_n618_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n867_), .A2(new_n872_), .A3(new_n618_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT61), .B(G155gat), .ZN(new_n876_));
  AND3_X1   g675(.A1(new_n874_), .A2(new_n875_), .A3(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n876_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(G1346gat));
  AOI21_X1  g678(.A(G162gat), .B1(new_n867_), .B2(new_n625_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n672_), .A2(G162gat), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n867_), .B2(new_n881_), .ZN(G1347gat));
  INV_X1    g681(.A(KEYINPUT123), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT122), .B(KEYINPUT62), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n319_), .A2(new_n365_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n826_), .A2(new_n698_), .A3(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n728_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n883_), .B(new_n884_), .C1(new_n888_), .C2(new_n224_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n884_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n224_), .B1(new_n890_), .B2(KEYINPUT123), .ZN(new_n891_));
  OAI221_X1 g690(.A(new_n891_), .B1(KEYINPUT123), .B2(new_n890_), .C1(new_n887_), .C2(new_n728_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n888_), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n889_), .B(new_n892_), .C1(new_n381_), .C2(new_n893_), .ZN(G1348gat));
  INV_X1    g693(.A(KEYINPUT124), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n886_), .A2(new_n895_), .A3(G176gat), .A4(new_n662_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n885_), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n836_), .A2(new_n410_), .A3(new_n662_), .A4(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n382_), .ZN(new_n899_));
  AOI21_X1  g698(.A(KEYINPUT124), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n898_), .A2(new_n225_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n896_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT125), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n902_), .B(new_n903_), .ZN(G1349gat));
  NOR2_X1   g703(.A1(new_n887_), .A2(new_n619_), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n905_), .B(new_n215_), .C1(KEYINPUT126), .C2(G183gat), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT126), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(G183gat), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n906_), .B1(new_n905_), .B2(new_n908_), .ZN(G1350gat));
  OAI21_X1  g708(.A(G190gat), .B1(new_n887_), .B2(new_n674_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n886_), .A2(new_n374_), .A3(new_n625_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1351gat));
  NOR4_X1   g711(.A1(new_n826_), .A2(new_n413_), .A3(new_n698_), .A4(new_n445_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n494_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g714(.A1(new_n913_), .A2(new_n662_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g716(.A(KEYINPUT63), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n618_), .B1(new_n918_), .B2(new_n349_), .ZN(new_n919_));
  XOR2_X1   g718(.A(new_n919_), .B(KEYINPUT127), .Z(new_n920_));
  NAND2_X1  g719(.A1(new_n913_), .A2(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n918_), .A2(new_n349_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n921_), .B(new_n922_), .ZN(G1354gat));
  NAND3_X1  g722(.A1(new_n913_), .A2(new_n347_), .A3(new_n625_), .ZN(new_n924_));
  AND2_X1   g723(.A1(new_n913_), .A2(new_n606_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n925_), .B2(new_n347_), .ZN(G1355gat));
endmodule


