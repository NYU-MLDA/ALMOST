//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n748_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_;
  INV_X1    g000(.A(KEYINPUT100), .ZN(new_n202_));
  XOR2_X1   g001(.A(G22gat), .B(G50gat), .Z(new_n203_));
  OR2_X1    g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT1), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  OAI211_X1 g006(.A(new_n204_), .B(new_n205_), .C1(new_n206_), .C2(new_n207_), .ZN(new_n208_));
  AND2_X1   g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  NOR3_X1   g009(.A1(new_n209_), .A2(new_n210_), .A3(KEYINPUT1), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n208_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT81), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n205_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT2), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT2), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n205_), .A2(new_n214_), .A3(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n219_));
  OR3_X1    g018(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n216_), .A2(new_n218_), .A3(new_n219_), .A4(new_n220_), .ZN(new_n221_));
  OR2_X1    g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(KEYINPUT82), .A3(new_n207_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT82), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n224_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  AND3_X1   g025(.A1(new_n221_), .A2(KEYINPUT83), .A3(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(KEYINPUT83), .B1(new_n221_), .B2(new_n226_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n213_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n203_), .B1(new_n229_), .B2(KEYINPUT29), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n221_), .A2(new_n226_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT83), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n221_), .A2(KEYINPUT83), .A3(new_n226_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n212_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT29), .ZN(new_n236_));
  INV_X1    g035(.A(new_n203_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT84), .B(KEYINPUT28), .ZN(new_n239_));
  AND3_X1   g038(.A1(new_n230_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n239_), .B1(new_n230_), .B2(new_n238_), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT85), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n230_), .A2(new_n238_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n239_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT85), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n230_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(G211gat), .B(G218gat), .Z(new_n249_));
  NOR2_X1   g048(.A1(G197gat), .A2(G204gat), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G197gat), .A2(G204gat), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n249_), .A2(KEYINPUT21), .A3(new_n251_), .A4(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n251_), .A2(KEYINPUT21), .A3(new_n252_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT21), .ZN(new_n255_));
  AND2_X1   g054(.A1(G197gat), .A2(G204gat), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n255_), .B1(new_n256_), .B2(new_n250_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G211gat), .B(G218gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n254_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n253_), .A2(new_n259_), .A3(KEYINPUT86), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(KEYINPUT86), .B1(new_n253_), .B2(new_n259_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G228gat), .A2(G233gat), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n263_), .B(new_n264_), .C1(new_n235_), .C2(new_n236_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G78gat), .B(G106gat), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n253_), .A2(new_n259_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n267_), .B1(new_n229_), .B2(KEYINPUT29), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n265_), .B(new_n266_), .C1(new_n264_), .C2(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n265_), .B1(new_n264_), .B2(new_n268_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n266_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n242_), .A2(new_n248_), .A3(new_n269_), .A4(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n245_), .A2(new_n247_), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n272_), .A2(new_n269_), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n273_), .B(KEYINPUT87), .C1(new_n274_), .C2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT87), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n275_), .A2(new_n277_), .A3(new_n248_), .A4(new_n242_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT26), .B(G190gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT25), .B(G183gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT77), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n280_), .A2(new_n281_), .A3(KEYINPUT77), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT24), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT24), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n289_), .B1(new_n291_), .B2(new_n287_), .ZN(new_n292_));
  AND2_X1   g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT23), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT78), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT78), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT23), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n293_), .B1(new_n295_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G183gat), .A2(G190gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT79), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT79), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n302_), .A2(G183gat), .A3(G190gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n294_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n292_), .B1(new_n299_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n286_), .A2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n295_), .A2(new_n297_), .A3(new_n293_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n308_), .B1(new_n304_), .B2(new_n294_), .ZN(new_n309_));
  OR2_X1    g108(.A1(G183gat), .A2(G190gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(G169gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n307_), .B(new_n314_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n315_));
  INV_X1    g114(.A(G176gat), .ZN(new_n316_));
  INV_X1    g115(.A(G169gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT22), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT22), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(G169gat), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n318_), .A2(new_n320_), .A3(KEYINPUT89), .ZN(new_n321_));
  AOI21_X1  g120(.A(KEYINPUT89), .B1(new_n318_), .B2(new_n320_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n316_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(KEYINPUT23), .B1(new_n301_), .B2(new_n303_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n310_), .B1(new_n324_), .B2(new_n298_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n323_), .A2(new_n325_), .A3(new_n290_), .ZN(new_n326_));
  INV_X1    g125(.A(G183gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT25), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT25), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(G183gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT88), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT88), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n328_), .A2(new_n330_), .A3(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n332_), .A2(new_n280_), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n292_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(new_n336_), .A3(new_n309_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n326_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n253_), .A2(new_n259_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n315_), .A2(new_n340_), .A3(KEYINPUT20), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G226gat), .A2(G233gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT19), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n307_), .A2(new_n314_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n263_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n343_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n326_), .A2(new_n337_), .A3(new_n267_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n346_), .A2(KEYINPUT20), .A3(new_n347_), .A4(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G8gat), .B(G36gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT18), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G64gat), .B(G92gat), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n351_), .B(new_n352_), .Z(new_n353_));
  NAND3_X1  g152(.A1(new_n344_), .A2(new_n349_), .A3(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT27), .ZN(new_n355_));
  INV_X1    g154(.A(new_n353_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n315_), .A2(new_n340_), .A3(KEYINPUT20), .A4(new_n347_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT96), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT20), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n360_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n361_), .A2(KEYINPUT96), .A3(new_n347_), .A4(new_n315_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n359_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT95), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n364_), .B1(new_n348_), .B2(KEYINPUT20), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT86), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n339_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(new_n260_), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n286_), .A2(new_n306_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n365_), .A2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n348_), .A2(new_n364_), .A3(KEYINPUT20), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n347_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n356_), .B1(new_n363_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT99), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  AND3_X1   g175(.A1(new_n348_), .A2(new_n364_), .A3(KEYINPUT20), .ZN(new_n377_));
  NOR3_X1   g176(.A1(new_n377_), .A2(new_n365_), .A3(new_n370_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n359_), .B(new_n362_), .C1(new_n378_), .C2(new_n347_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(KEYINPUT99), .A3(new_n356_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n355_), .B1(new_n376_), .B2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G1gat), .B(G29gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(G85gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT0), .B(G57gat), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n383_), .B(new_n384_), .Z(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT4), .ZN(new_n387_));
  XOR2_X1   g186(.A(G127gat), .B(G134gat), .Z(new_n388_));
  XNOR2_X1  g187(.A(G113gat), .B(G120gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n229_), .A2(new_n387_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT90), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT90), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n229_), .A2(new_n393_), .A3(new_n387_), .A4(new_n390_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G225gat), .A2(G233gat), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n229_), .A2(new_n390_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n390_), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n399_), .B(new_n213_), .C1(new_n227_), .C2(new_n228_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n398_), .A2(new_n400_), .A3(KEYINPUT4), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n395_), .A2(KEYINPUT91), .A3(new_n397_), .A4(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n398_), .A2(new_n400_), .A3(new_n396_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT92), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n398_), .A2(new_n400_), .A3(KEYINPUT92), .A4(new_n396_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n402_), .A2(new_n407_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n401_), .A2(new_n397_), .ZN(new_n409_));
  AOI21_X1  g208(.A(KEYINPUT91), .B1(new_n409_), .B2(new_n395_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n386_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT91), .ZN(new_n412_));
  INV_X1    g211(.A(new_n395_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n401_), .A2(new_n397_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n412_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n415_), .A2(new_n385_), .A3(new_n402_), .A4(new_n407_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n411_), .A2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n347_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n348_), .A2(KEYINPUT20), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n347_), .B1(new_n361_), .B2(new_n315_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n356_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n422_), .A2(new_n354_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n423_), .A2(KEYINPUT27), .ZN(new_n424_));
  NOR4_X1   g223(.A1(new_n279_), .A2(new_n381_), .A3(new_n417_), .A4(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT98), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n411_), .A2(new_n416_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n353_), .A2(KEYINPUT32), .ZN(new_n428_));
  OAI211_X1 g227(.A(KEYINPUT97), .B(new_n428_), .C1(new_n363_), .C2(new_n373_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT97), .B1(new_n379_), .B2(new_n428_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n344_), .A2(new_n349_), .ZN(new_n432_));
  XOR2_X1   g231(.A(new_n428_), .B(KEYINPUT94), .Z(new_n433_));
  OAI22_X1  g232(.A1(new_n430_), .A2(new_n431_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n426_), .B1(new_n427_), .B2(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n433_), .A2(new_n432_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n428_), .B1(new_n363_), .B2(new_n373_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT97), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n436_), .B1(new_n439_), .B2(new_n429_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n440_), .A2(new_n417_), .A3(KEYINPUT98), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n395_), .A2(new_n396_), .A3(new_n401_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n398_), .A2(new_n400_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT93), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT93), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n398_), .A2(new_n400_), .A3(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n444_), .A2(new_n397_), .A3(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n442_), .A2(new_n386_), .A3(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n423_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT33), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n449_), .B1(new_n450_), .B2(new_n416_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n402_), .A2(new_n407_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n452_), .A2(KEYINPUT33), .A3(new_n385_), .A4(new_n415_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n435_), .A2(new_n441_), .A3(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n425_), .B1(new_n455_), .B2(new_n279_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n369_), .B(KEYINPUT30), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G227gat), .A2(G233gat), .ZN(new_n458_));
  INV_X1    g257(.A(G15gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(G71gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(G99gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n457_), .B(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(new_n390_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT80), .B(G43gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT31), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n464_), .B(new_n466_), .Z(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n202_), .B1(new_n456_), .B2(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n381_), .A2(new_n424_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n468_), .A2(new_n470_), .A3(new_n427_), .A4(new_n279_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n279_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n440_), .A2(new_n417_), .ZN(new_n473_));
  AOI22_X1  g272(.A1(new_n473_), .A2(new_n426_), .B1(new_n453_), .B2(new_n451_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n472_), .B1(new_n474_), .B2(new_n441_), .ZN(new_n475_));
  OAI211_X1 g274(.A(KEYINPUT100), .B(new_n467_), .C1(new_n475_), .C2(new_n425_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n469_), .A2(new_n471_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(G1gat), .ZN(new_n478_));
  INV_X1    g277(.A(G8gat), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT14), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n480_), .A2(KEYINPUT74), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(KEYINPUT74), .ZN(new_n482_));
  XOR2_X1   g281(.A(G15gat), .B(G22gat), .Z(new_n483_));
  NOR3_X1   g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(G1gat), .B(G8gat), .Z(new_n485_));
  OR2_X1    g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n485_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G29gat), .B(G36gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G43gat), .B(G50gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  XOR2_X1   g290(.A(new_n488_), .B(new_n491_), .Z(new_n492_));
  NAND3_X1  g291(.A1(new_n492_), .A2(G229gat), .A3(G233gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n491_), .B(KEYINPUT15), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n488_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G229gat), .A2(G233gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n486_), .A2(new_n487_), .A3(new_n491_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n493_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G113gat), .B(G141gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G169gat), .B(G197gat), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n500_), .B(new_n501_), .Z(new_n502_));
  XOR2_X1   g301(.A(new_n499_), .B(new_n502_), .Z(new_n503_));
  AND2_X1   g302(.A1(new_n477_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT6), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT65), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT65), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT6), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G99gat), .A2(G106gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n506_), .A2(new_n508_), .A3(G99gat), .A4(G106gat), .ZN(new_n512_));
  INV_X1    g311(.A(G99gat), .ZN(new_n513_));
  INV_X1    g312(.A(G106gat), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(new_n514_), .A3(KEYINPUT66), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT7), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT7), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n517_), .A2(new_n513_), .A3(new_n514_), .A4(KEYINPUT66), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n511_), .A2(new_n512_), .A3(new_n516_), .A4(new_n518_), .ZN(new_n519_));
  OR2_X1    g318(.A1(G85gat), .A2(G92gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G85gat), .A2(G92gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n519_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT8), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n525_), .B1(new_n522_), .B2(KEYINPUT67), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n519_), .A2(new_n523_), .A3(new_n526_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT9), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT64), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n521_), .A2(new_n531_), .A3(new_n530_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n531_), .B1(new_n521_), .B2(new_n530_), .ZN(new_n533_));
  OAI221_X1 g332(.A(new_n520_), .B1(new_n530_), .B2(new_n521_), .C1(new_n532_), .C2(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(KEYINPUT10), .B(G99gat), .Z(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n514_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n534_), .A2(new_n512_), .A3(new_n511_), .A4(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n528_), .A2(new_n529_), .A3(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT69), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT69), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n528_), .A2(new_n540_), .A3(new_n529_), .A4(new_n537_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n539_), .A2(new_n494_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT71), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n538_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G232gat), .A2(G233gat), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n546_), .B(KEYINPUT34), .Z(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT70), .B(KEYINPUT35), .ZN(new_n548_));
  AOI22_X1  g347(.A1(new_n545_), .A2(new_n491_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n539_), .A2(KEYINPUT71), .A3(new_n494_), .A4(new_n541_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n544_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n547_), .A2(new_n548_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  XOR2_X1   g352(.A(new_n552_), .B(KEYINPUT72), .Z(new_n554_));
  NAND3_X1  g353(.A1(new_n549_), .A2(new_n542_), .A3(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G190gat), .B(G218gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G134gat), .B(G162gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n559_), .A2(KEYINPUT36), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n556_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n553_), .A2(new_n555_), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n559_), .B(KEYINPUT36), .Z(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n561_), .A2(new_n564_), .A3(KEYINPUT37), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n556_), .A2(KEYINPUT73), .ZN(new_n566_));
  INV_X1    g365(.A(new_n563_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT73), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n567_), .B1(new_n562_), .B2(new_n568_), .ZN(new_n569_));
  AOI22_X1  g368(.A1(new_n566_), .A2(new_n569_), .B1(new_n556_), .B2(new_n560_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n565_), .B1(new_n570_), .B2(KEYINPUT37), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G230gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G57gat), .B(G64gat), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT11), .ZN(new_n574_));
  XOR2_X1   g373(.A(G71gat), .B(G78gat), .Z(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n574_), .A2(new_n575_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n573_), .A2(KEYINPUT11), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n577_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n538_), .A2(new_n581_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n528_), .A2(new_n580_), .A3(new_n529_), .A4(new_n537_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n572_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n584_), .A2(KEYINPUT68), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n539_), .A2(KEYINPUT12), .A3(new_n541_), .A4(new_n581_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(KEYINPUT12), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(new_n582_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n586_), .A2(new_n588_), .A3(new_n572_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n582_), .A2(new_n583_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n572_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n590_), .A2(KEYINPUT68), .A3(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n585_), .A2(new_n589_), .A3(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G120gat), .B(G148gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT5), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G176gat), .B(G204gat), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n595_), .B(new_n596_), .Z(new_n597_));
  XNOR2_X1  g396(.A(new_n593_), .B(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT13), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(G127gat), .B(G155gat), .Z(new_n601_));
  XNOR2_X1  g400(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G183gat), .B(G211gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT17), .ZN(new_n606_));
  NOR3_X1   g405(.A1(new_n605_), .A2(KEYINPUT75), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n488_), .B(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(new_n581_), .ZN(new_n610_));
  AOI211_X1 g409(.A(new_n607_), .B(new_n610_), .C1(new_n606_), .C2(new_n605_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n610_), .A2(new_n607_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n571_), .A2(new_n600_), .A3(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n504_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n616_), .A2(new_n478_), .A3(new_n417_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT38), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT101), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(new_n618_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT102), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n566_), .A2(new_n569_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(new_n561_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n477_), .A2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n598_), .B(KEYINPUT13), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(new_n503_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n627_), .A2(new_n614_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n625_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G1gat), .B1(new_n630_), .B2(new_n427_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n620_), .A2(new_n622_), .A3(new_n631_), .ZN(G1324gat));
  INV_X1    g431(.A(new_n470_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n616_), .A2(new_n479_), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT39), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n477_), .A2(new_n633_), .A3(new_n624_), .A4(new_n628_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT103), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n638_), .A2(G8gat), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n636_), .A2(new_n637_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n635_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  AND4_X1   g440(.A1(new_n635_), .A2(new_n638_), .A3(G8gat), .A4(new_n640_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n634_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT40), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  OAI211_X1 g444(.A(KEYINPUT40), .B(new_n634_), .C1(new_n641_), .C2(new_n642_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(G1325gat));
  NAND3_X1  g446(.A1(new_n616_), .A2(new_n459_), .A3(new_n468_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n629_), .A2(new_n468_), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n649_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n650_));
  AOI21_X1  g449(.A(KEYINPUT41), .B1(new_n649_), .B2(G15gat), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n648_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT104), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  OAI211_X1 g453(.A(KEYINPUT104), .B(new_n648_), .C1(new_n650_), .C2(new_n651_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1326gat));
  INV_X1    g455(.A(G22gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n657_), .B1(new_n629_), .B2(new_n472_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n658_), .B(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n472_), .A2(new_n657_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT106), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n616_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n660_), .A2(new_n663_), .ZN(G1327gat));
  NAND2_X1  g463(.A1(new_n614_), .A2(new_n570_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n665_), .A2(new_n600_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n504_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(G29gat), .B1(new_n668_), .B2(new_n417_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n627_), .A2(new_n613_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n476_), .A2(new_n471_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n425_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n440_), .A2(new_n417_), .A3(KEYINPUT98), .ZN(new_n674_));
  AOI21_X1  g473(.A(KEYINPUT98), .B1(new_n440_), .B2(new_n417_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n416_), .A2(new_n450_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n449_), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n676_), .A2(new_n453_), .A3(new_n677_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n674_), .A2(new_n675_), .A3(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n673_), .B1(new_n679_), .B2(new_n472_), .ZN(new_n680_));
  AOI21_X1  g479(.A(KEYINPUT100), .B1(new_n680_), .B2(new_n467_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n571_), .B1(new_n672_), .B2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT43), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT43), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n477_), .A2(new_n684_), .A3(new_n571_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n671_), .B1(new_n683_), .B2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(KEYINPUT107), .B1(new_n686_), .B2(KEYINPUT44), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n477_), .A2(new_n684_), .A3(new_n571_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n684_), .B1(new_n477_), .B2(new_n571_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n670_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT107), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n690_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n693_));
  AOI22_X1  g492(.A1(new_n687_), .A2(new_n693_), .B1(KEYINPUT44), .B2(new_n686_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n417_), .A2(G29gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n669_), .B1(new_n694_), .B2(new_n695_), .ZN(G1328gat));
  INV_X1    g495(.A(G36gat), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n633_), .A2(new_n697_), .ZN(new_n698_));
  OR3_X1    g497(.A1(new_n667_), .A2(KEYINPUT45), .A3(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(KEYINPUT45), .B1(new_n667_), .B2(new_n698_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  OAI211_X1 g500(.A(KEYINPUT44), .B(new_n670_), .C1(new_n688_), .C2(new_n689_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(new_n633_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n687_), .B2(new_n693_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n701_), .B1(new_n704_), .B2(new_n697_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT46), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  OAI211_X1 g506(.A(KEYINPUT46), .B(new_n701_), .C1(new_n704_), .C2(new_n697_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1329gat));
  INV_X1    g508(.A(G43gat), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n467_), .A2(new_n710_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n686_), .A2(KEYINPUT107), .A3(KEYINPUT44), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n691_), .B1(new_n690_), .B2(new_n692_), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n702_), .B(new_n711_), .C1(new_n712_), .C2(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n710_), .B1(new_n667_), .B2(new_n467_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n714_), .A2(new_n715_), .A3(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1330gat));
  AOI21_X1  g518(.A(G50gat), .B1(new_n668_), .B2(new_n472_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n472_), .A2(G50gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n694_), .B2(new_n721_), .ZN(G1331gat));
  INV_X1    g521(.A(new_n503_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n477_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n561_), .A2(KEYINPUT37), .A3(new_n564_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT37), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n624_), .B2(new_n727_), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n725_), .A2(new_n728_), .A3(new_n613_), .A4(new_n600_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n730_), .A2(KEYINPUT109), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(KEYINPUT109), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n731_), .A2(new_n417_), .A3(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(G57gat), .ZN(new_n734_));
  AND4_X1   g533(.A1(new_n723_), .A2(new_n625_), .A3(new_n613_), .A4(new_n600_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n427_), .A2(new_n734_), .ZN(new_n736_));
  AOI22_X1  g535(.A1(new_n733_), .A2(new_n734_), .B1(new_n735_), .B2(new_n736_), .ZN(G1332gat));
  INV_X1    g536(.A(G64gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n738_), .B1(new_n735_), .B2(new_n633_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT48), .Z(new_n740_));
  NAND3_X1  g539(.A1(new_n730_), .A2(new_n738_), .A3(new_n633_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1333gat));
  INV_X1    g541(.A(G71gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n735_), .B2(new_n468_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT49), .Z(new_n745_));
  NAND3_X1  g544(.A1(new_n730_), .A2(new_n743_), .A3(new_n468_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1334gat));
  INV_X1    g546(.A(G78gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n735_), .B2(new_n472_), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT50), .Z(new_n750_));
  NAND3_X1  g549(.A1(new_n730_), .A2(new_n748_), .A3(new_n472_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1335gat));
  NOR3_X1   g551(.A1(new_n724_), .A2(new_n626_), .A3(new_n665_), .ZN(new_n753_));
  INV_X1    g552(.A(G85gat), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n753_), .A2(new_n754_), .A3(new_n417_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n683_), .A2(new_n685_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n626_), .A2(new_n503_), .A3(new_n613_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT110), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n758_), .B(new_n759_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n760_), .A2(new_n417_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n755_), .B1(new_n761_), .B2(new_n754_), .ZN(G1336gat));
  AOI21_X1  g561(.A(G92gat), .B1(new_n753_), .B2(new_n633_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n633_), .A2(G92gat), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT111), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n763_), .B1(new_n760_), .B2(new_n765_), .ZN(G1337gat));
  NAND3_X1  g565(.A1(new_n753_), .A2(new_n468_), .A3(new_n535_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT112), .ZN(new_n768_));
  OAI21_X1  g567(.A(G99gat), .B1(new_n758_), .B2(new_n467_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT51), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n768_), .A2(new_n769_), .A3(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1338gat));
  NAND3_X1  g573(.A1(new_n753_), .A2(new_n514_), .A3(new_n472_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n472_), .B(new_n757_), .C1(new_n688_), .C2(new_n689_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n776_), .A2(new_n777_), .A3(G106gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n776_), .B2(G106gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g580(.A(new_n499_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n495_), .A2(new_n497_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n496_), .B1(new_n783_), .B2(KEYINPUT117), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n784_), .B1(KEYINPUT117), .B2(new_n783_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n502_), .B1(new_n492_), .B2(new_n496_), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n782_), .A2(new_n502_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n593_), .A2(new_n597_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n586_), .A2(new_n588_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n591_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n791_), .A2(KEYINPUT55), .A3(new_n589_), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n586_), .A2(new_n588_), .A3(new_n572_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n572_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n793_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n792_), .A2(new_n796_), .A3(KEYINPUT115), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT115), .B1(new_n792_), .B2(new_n796_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n597_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT56), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  OAI211_X1 g600(.A(KEYINPUT56), .B(new_n597_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n789_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n803_), .A2(KEYINPUT58), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n571_), .B1(new_n803_), .B2(KEYINPUT58), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n598_), .A2(new_n787_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n801_), .A2(new_n808_), .A3(new_n802_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n503_), .B(new_n788_), .C1(new_n802_), .C2(new_n808_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n807_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT57), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n624_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n807_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n503_), .A2(new_n788_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n597_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n793_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n790_), .A2(KEYINPUT55), .A3(new_n591_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n817_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n792_), .A2(new_n796_), .A3(KEYINPUT115), .ZN(new_n821_));
  AOI211_X1 g620(.A(new_n800_), .B(new_n816_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n815_), .B1(new_n822_), .B2(KEYINPUT116), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n801_), .A2(new_n808_), .A3(new_n802_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n814_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT57), .B1(new_n825_), .B2(new_n570_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n806_), .B1(new_n813_), .B2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT119), .B1(new_n827_), .B2(new_n613_), .ZN(new_n828_));
  OR2_X1    g627(.A1(new_n804_), .A2(new_n805_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n812_), .B1(new_n811_), .B2(new_n624_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n825_), .A2(KEYINPUT57), .A3(new_n570_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n829_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(new_n833_), .A3(new_n614_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n728_), .A2(new_n723_), .A3(new_n613_), .A4(new_n626_), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT114), .B1(new_n835_), .B2(KEYINPUT113), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT113), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n615_), .A2(new_n837_), .A3(new_n838_), .A4(new_n723_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n836_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n835_), .A2(KEYINPUT113), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n840_), .A2(new_n843_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n836_), .A2(new_n839_), .A3(new_n842_), .A4(new_n841_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n828_), .A2(new_n834_), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n470_), .A2(new_n279_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n467_), .A2(new_n848_), .A3(new_n427_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n850_), .A2(KEYINPUT59), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n847_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(G113gat), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n723_), .A2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT118), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n832_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n827_), .A2(KEYINPUT118), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n856_), .A2(new_n857_), .A3(new_n614_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n850_), .B1(new_n858_), .B2(new_n846_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n852_), .B(new_n854_), .C1(new_n859_), .C2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n614_), .B1(new_n827_), .B2(KEYINPUT118), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n832_), .A2(new_n855_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n846_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n849_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n853_), .B1(new_n865_), .B2(new_n723_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n861_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n861_), .A2(new_n866_), .A3(KEYINPUT120), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1340gat));
  XOR2_X1   g670(.A(KEYINPUT121), .B(G120gat), .Z(new_n872_));
  OR2_X1    g671(.A1(new_n872_), .A2(KEYINPUT60), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n626_), .B2(KEYINPUT60), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n864_), .A2(new_n849_), .A3(new_n873_), .A4(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT122), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n875_), .B(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n852_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n878_), .A2(new_n626_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n877_), .B1(new_n872_), .B2(new_n879_), .ZN(G1341gat));
  OAI21_X1  g679(.A(G127gat), .B1(new_n878_), .B2(new_n614_), .ZN(new_n881_));
  OR2_X1    g680(.A1(new_n614_), .A2(G127gat), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n865_), .B2(new_n882_), .ZN(G1342gat));
  OAI21_X1  g682(.A(G134gat), .B1(new_n878_), .B2(new_n728_), .ZN(new_n884_));
  OR2_X1    g683(.A1(new_n624_), .A2(G134gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n865_), .B2(new_n885_), .ZN(G1343gat));
  NOR3_X1   g685(.A1(new_n468_), .A2(new_n427_), .A3(new_n279_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n864_), .A2(new_n470_), .A3(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(new_n723_), .ZN(new_n889_));
  XOR2_X1   g688(.A(KEYINPUT123), .B(G141gat), .Z(new_n890_));
  XNOR2_X1  g689(.A(new_n889_), .B(new_n890_), .ZN(G1344gat));
  OR2_X1    g690(.A1(new_n888_), .A2(new_n626_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g692(.A1(new_n888_), .A2(new_n614_), .ZN(new_n894_));
  XOR2_X1   g693(.A(KEYINPUT61), .B(G155gat), .Z(new_n895_));
  XNOR2_X1  g694(.A(new_n894_), .B(new_n895_), .ZN(G1346gat));
  OAI21_X1  g695(.A(G162gat), .B1(new_n888_), .B2(new_n728_), .ZN(new_n897_));
  OR2_X1    g696(.A1(new_n624_), .A2(G162gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n888_), .B2(new_n898_), .ZN(G1347gat));
  NOR4_X1   g698(.A1(new_n467_), .A2(new_n472_), .A3(new_n470_), .A4(new_n417_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n847_), .A2(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n901_), .A2(new_n723_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n902_), .A2(KEYINPUT62), .A3(new_n317_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n847_), .A2(new_n900_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n503_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n904_), .B1(new_n906_), .B2(G169gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n902_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n903_), .B1(new_n907_), .B2(new_n908_), .ZN(G1348gat));
  NAND4_X1  g708(.A1(new_n864_), .A2(G176gat), .A3(new_n600_), .A4(new_n900_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(G176gat), .B1(new_n905_), .B2(new_n600_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n910_), .A2(new_n911_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n912_), .A2(new_n913_), .A3(new_n914_), .ZN(G1349gat));
  AND3_X1   g714(.A1(new_n864_), .A2(new_n613_), .A3(new_n900_), .ZN(new_n916_));
  OR2_X1    g715(.A1(new_n916_), .A2(KEYINPUT125), .ZN(new_n917_));
  AOI21_X1  g716(.A(G183gat), .B1(new_n916_), .B2(KEYINPUT125), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n614_), .B1(new_n332_), .B2(new_n334_), .ZN(new_n919_));
  AOI22_X1  g718(.A1(new_n917_), .A2(new_n918_), .B1(new_n905_), .B2(new_n919_), .ZN(G1350gat));
  NAND3_X1  g719(.A1(new_n905_), .A2(new_n280_), .A3(new_n570_), .ZN(new_n921_));
  OAI21_X1  g720(.A(G190gat), .B1(new_n901_), .B2(new_n728_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT126), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n921_), .A2(new_n922_), .A3(KEYINPUT126), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n925_), .A2(new_n926_), .ZN(G1351gat));
  NOR4_X1   g726(.A1(new_n468_), .A2(new_n470_), .A3(new_n417_), .A4(new_n279_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n864_), .A2(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(new_n503_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g731(.A1(new_n930_), .A2(new_n600_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g733(.A(new_n614_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n935_));
  INV_X1    g734(.A(new_n935_), .ZN(new_n936_));
  OAI21_X1  g735(.A(KEYINPUT127), .B1(new_n929_), .B2(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT127), .ZN(new_n939_));
  NAND4_X1  g738(.A1(new_n864_), .A2(new_n939_), .A3(new_n928_), .A4(new_n935_), .ZN(new_n940_));
  AND3_X1   g739(.A1(new_n937_), .A2(new_n938_), .A3(new_n940_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n938_), .B1(new_n937_), .B2(new_n940_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n941_), .A2(new_n942_), .ZN(G1354gat));
  OAI21_X1  g742(.A(G218gat), .B1(new_n929_), .B2(new_n728_), .ZN(new_n944_));
  OR2_X1    g743(.A1(new_n624_), .A2(G218gat), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n944_), .B1(new_n929_), .B2(new_n945_), .ZN(G1355gat));
endmodule


