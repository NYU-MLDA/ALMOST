//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 1 0 1 1 0 1 0 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 0 1 0 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n946_, new_n947_,
    new_n948_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n961_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n972_, new_n973_, new_n974_;
  XOR2_X1   g000(.A(G134gat), .B(G162gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G190gat), .B(G218gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT36), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n204_), .A2(new_n205_), .ZN(new_n207_));
  AND2_X1   g006(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n208_));
  NOR2_X1   g007(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n209_));
  OAI22_X1  g008(.A1(new_n208_), .A2(new_n209_), .B1(G99gat), .B2(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n211_));
  INV_X1    g010(.A(G99gat), .ZN(new_n212_));
  INV_X1    g011(.A(G106gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n210_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT6), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT6), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  AND3_X1   g018(.A1(new_n217_), .A2(new_n219_), .A3(KEYINPUT67), .ZN(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT67), .B1(new_n217_), .B2(new_n219_), .ZN(new_n221_));
  NOR3_X1   g020(.A1(new_n215_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  OR2_X1    g021(.A1(G85gat), .A2(G92gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G85gat), .A2(G92gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT8), .B1(new_n222_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n225_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT8), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n215_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n217_), .A2(new_n219_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n229_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(G85gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n234_), .A2(KEYINPUT9), .ZN(new_n235_));
  AND2_X1   g034(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n235_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n223_), .A2(KEYINPUT9), .A3(new_n224_), .ZN(new_n239_));
  OR2_X1    g038(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(new_n213_), .A3(new_n241_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n238_), .A2(new_n239_), .A3(new_n242_), .A4(new_n231_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT65), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n239_), .A2(new_n231_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n245_), .A2(new_n246_), .A3(new_n242_), .A4(new_n238_), .ZN(new_n247_));
  AOI22_X1  g046(.A1(new_n226_), .A2(new_n233_), .B1(new_n244_), .B2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G29gat), .B(G36gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G43gat), .B(G50gat), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n250_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n248_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n247_), .A2(new_n244_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n231_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n217_), .A2(new_n219_), .A3(KEYINPUT67), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n257_), .A2(new_n258_), .A3(new_n210_), .A4(new_n214_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n228_), .B1(new_n259_), .B2(new_n227_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n255_), .B1(new_n260_), .B2(new_n232_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT72), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT15), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n253_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n251_), .A2(KEYINPUT15), .A3(new_n252_), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n261_), .A2(new_n262_), .A3(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n262_), .B1(new_n261_), .B2(new_n266_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n254_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT73), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G232gat), .A2(G233gat), .ZN(new_n271_));
  XOR2_X1   g070(.A(new_n271_), .B(KEYINPUT34), .Z(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT71), .B(KEYINPUT35), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  AND3_X1   g073(.A1(new_n269_), .A2(new_n270_), .A3(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n270_), .B1(new_n269_), .B2(new_n274_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n272_), .A2(new_n273_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n278_), .B1(new_n274_), .B2(KEYINPUT74), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n279_), .B1(KEYINPUT74), .B2(new_n274_), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n254_), .B(new_n280_), .C1(new_n267_), .C2(new_n268_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT75), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n206_), .B(new_n207_), .C1(new_n277_), .C2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n276_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n269_), .A2(new_n270_), .A3(new_n274_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n281_), .B(KEYINPUT75), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n287_), .A2(new_n288_), .A3(new_n205_), .A4(new_n204_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT76), .B(KEYINPUT37), .ZN(new_n290_));
  AND3_X1   g089(.A1(new_n284_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(KEYINPUT76), .A2(KEYINPUT37), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n292_), .B1(new_n284_), .B2(new_n289_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(G64gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G57gat), .ZN(new_n296_));
  INV_X1    g095(.A(G57gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G64gat), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G71gat), .B(G78gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n299_), .A2(new_n300_), .A3(KEYINPUT11), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n299_), .A2(KEYINPUT11), .ZN(new_n302_));
  INV_X1    g101(.A(new_n300_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n296_), .A2(new_n298_), .A3(KEYINPUT11), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n301_), .B1(new_n302_), .B2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G15gat), .B(G22gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G1gat), .A2(G8gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT14), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(G1gat), .ZN(new_n311_));
  INV_X1    g110(.A(G8gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n308_), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n310_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n310_), .A2(new_n314_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G231gat), .A2(G233gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n317_), .A2(new_n318_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n306_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n321_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n306_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n319_), .A3(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G127gat), .B(G155gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT16), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G183gat), .B(G211gat), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n327_), .A2(new_n328_), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n322_), .A2(new_n325_), .A3(KEYINPUT17), .A4(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n306_), .A2(KEYINPUT68), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT68), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n334_), .B(new_n301_), .C1(new_n302_), .C2(new_n305_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n336_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n331_), .A2(KEYINPUT17), .ZN(new_n338_));
  OR3_X1    g137(.A1(new_n329_), .A2(new_n330_), .A3(KEYINPUT17), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  NOR3_X1   g139(.A1(new_n320_), .A2(new_n336_), .A3(new_n321_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n332_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT77), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n294_), .A2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G78gat), .B(G106gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT93), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT28), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G155gat), .A2(G162gat), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n350_), .A2(KEYINPUT1), .ZN(new_n351_));
  NOR2_X1   g150(.A1(G155gat), .A2(G162gat), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n350_), .B1(new_n352_), .B2(KEYINPUT1), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT86), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n351_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  OAI211_X1 g154(.A(KEYINPUT86), .B(new_n350_), .C1(new_n352_), .C2(KEYINPUT1), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G141gat), .A2(G148gat), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT85), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(KEYINPUT85), .A2(G141gat), .A3(G148gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(G141gat), .A2(G148gat), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n352_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT88), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(new_n366_), .A3(new_n350_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n350_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT88), .B1(new_n368_), .B2(new_n352_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT2), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n360_), .A2(new_n372_), .A3(new_n361_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(KEYINPUT87), .A2(KEYINPUT3), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n363_), .A2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n376_));
  OAI22_X1  g175(.A1(KEYINPUT87), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n373_), .A2(new_n375_), .A3(new_n376_), .A4(new_n377_), .ZN(new_n378_));
  AOI22_X1  g177(.A1(new_n357_), .A2(new_n364_), .B1(new_n371_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT29), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n349_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n357_), .A2(new_n364_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n371_), .A2(new_n378_), .ZN(new_n383_));
  AND4_X1   g182(.A1(new_n349_), .A2(new_n382_), .A3(new_n380_), .A4(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT89), .B1(new_n381_), .B2(new_n384_), .ZN(new_n385_));
  XOR2_X1   g184(.A(G22gat), .B(G50gat), .Z(new_n386_));
  NAND2_X1  g185(.A1(new_n382_), .A2(new_n383_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT28), .B1(new_n387_), .B2(KEYINPUT29), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT89), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n379_), .A2(new_n349_), .A3(new_n380_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n388_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n385_), .A2(new_n386_), .A3(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n386_), .B1(new_n385_), .B2(new_n391_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n348_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n385_), .A2(new_n391_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n386_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n348_), .A2(KEYINPUT94), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n385_), .A2(new_n391_), .A3(new_n386_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n379_), .A2(new_n380_), .ZN(new_n401_));
  OR2_X1    g200(.A1(G197gat), .A2(G204gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G197gat), .A2(G204gat), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(KEYINPUT21), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT91), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(G218gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(G211gat), .ZN(new_n408_));
  INV_X1    g207(.A(G211gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(G218gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT21), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n402_), .A2(new_n403_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n411_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(KEYINPUT92), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n412_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT92), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n402_), .A2(new_n417_), .A3(new_n403_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  AOI22_X1  g218(.A1(new_n406_), .A2(new_n414_), .B1(new_n415_), .B2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT90), .B1(new_n401_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n406_), .A2(new_n414_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n419_), .A2(new_n415_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT90), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n424_), .B(new_n425_), .C1(new_n380_), .C2(new_n379_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n421_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G228gat), .A2(G233gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n421_), .A2(G228gat), .A3(G233gat), .A4(new_n426_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n394_), .A2(new_n400_), .A3(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n431_), .B1(new_n394_), .B2(new_n400_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  XOR2_X1   g233(.A(G127gat), .B(G134gat), .Z(new_n435_));
  XOR2_X1   g234(.A(G113gat), .B(G120gat), .Z(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  OR2_X1    g237(.A1(new_n362_), .A2(new_n363_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n439_), .B1(new_n356_), .B2(new_n355_), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n375_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n370_), .B1(new_n373_), .B2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n438_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n382_), .A2(new_n383_), .A3(new_n437_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(KEYINPUT4), .A3(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT4), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n387_), .A2(new_n446_), .A3(new_n438_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G225gat), .A2(G233gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT96), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G1gat), .B(G29gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G57gat), .B(G85gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n450_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n451_), .A2(new_n456_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n456_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n450_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n461_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n460_), .B1(new_n462_), .B2(new_n457_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n459_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT23), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n465_), .A2(G183gat), .A3(G190gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(G183gat), .ZN(new_n468_));
  INV_X1    g267(.A(G190gat), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT23), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT81), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  OAI211_X1 g271(.A(KEYINPUT81), .B(KEYINPUT23), .C1(new_n468_), .C2(new_n469_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n467_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT25), .B(G183gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT26), .B(G190gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G169gat), .A2(G176gat), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT80), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(KEYINPUT80), .A2(G169gat), .A3(G176gat), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n480_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(G169gat), .A2(G176gat), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT24), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n478_), .A2(new_n485_), .A3(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n483_), .A2(new_n484_), .ZN(new_n490_));
  XOR2_X1   g289(.A(KEYINPUT82), .B(G176gat), .Z(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT22), .B(G169gat), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n490_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n470_), .A2(new_n466_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n494_), .B1(G183gat), .B2(G190gat), .ZN(new_n495_));
  AOI22_X1  g294(.A1(new_n475_), .A2(new_n489_), .B1(new_n493_), .B2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT30), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT84), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n493_), .A2(new_n495_), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n476_), .A2(new_n477_), .B1(new_n487_), .B2(new_n486_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n485_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n499_), .B1(new_n501_), .B2(new_n474_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT30), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT84), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n498_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G227gat), .A2(G233gat), .ZN(new_n507_));
  INV_X1    g306(.A(G15gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(G71gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(new_n212_), .ZN(new_n511_));
  XOR2_X1   g310(.A(KEYINPUT83), .B(G43gat), .Z(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n506_), .A2(new_n513_), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n511_), .B(new_n512_), .Z(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n505_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  XOR2_X1   g316(.A(new_n437_), .B(KEYINPUT31), .Z(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n514_), .A2(new_n516_), .A3(new_n518_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n464_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT20), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n523_), .B1(new_n496_), .B2(new_n420_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(G183gat), .A2(G190gat), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n493_), .B1(new_n474_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n480_), .A2(new_n481_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n478_), .A2(new_n494_), .A3(new_n488_), .A4(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT95), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT95), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n500_), .A2(new_n530_), .A3(new_n494_), .A4(new_n527_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n526_), .A2(new_n529_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n424_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n524_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G226gat), .A2(G233gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT19), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(G8gat), .B(G36gat), .Z(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT18), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G64gat), .B(G92gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n523_), .B1(new_n424_), .B2(new_n502_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n420_), .A2(new_n526_), .A3(new_n529_), .A4(new_n531_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n536_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n537_), .A2(new_n541_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n541_), .ZN(new_n547_));
  OAI211_X1 g346(.A(KEYINPUT20), .B(new_n544_), .C1(new_n496_), .C2(new_n420_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n532_), .A2(new_n424_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n544_), .B1(new_n524_), .B2(new_n533_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n547_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(KEYINPUT27), .B1(new_n546_), .B2(new_n552_), .ZN(new_n553_));
  AND3_X1   g352(.A1(new_n524_), .A2(new_n533_), .A3(new_n544_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n420_), .A2(new_n526_), .A3(new_n528_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n544_), .B1(new_n542_), .B2(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n547_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT99), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT99), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n559_), .B(new_n547_), .C1(new_n554_), .C2(new_n556_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n546_), .A2(KEYINPUT27), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n553_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n434_), .A2(new_n522_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n394_), .A2(new_n400_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n431_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n394_), .A2(new_n400_), .A3(new_n431_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n464_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n443_), .A2(new_n450_), .A3(new_n444_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n456_), .B(new_n570_), .C1(new_n448_), .C2(new_n450_), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n546_), .A2(new_n552_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT98), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT33), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n573_), .B1(new_n463_), .B2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n451_), .A2(new_n458_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n576_), .A2(KEYINPUT98), .A3(KEYINPUT33), .A4(new_n460_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n463_), .A2(new_n574_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n572_), .A2(new_n575_), .A3(new_n577_), .A4(new_n578_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n541_), .A2(KEYINPUT32), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n580_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n537_), .A2(new_n545_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n464_), .B(new_n581_), .C1(new_n580_), .C2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n583_), .ZN(new_n584_));
  AOI22_X1  g383(.A1(new_n569_), .A2(new_n563_), .B1(new_n434_), .B2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n520_), .A2(new_n521_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n564_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT13), .ZN(new_n588_));
  AND2_X1   g387(.A1(G230gat), .A2(G233gat), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT69), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n333_), .A2(new_n335_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n248_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n248_), .A2(new_n591_), .ZN(new_n593_));
  OAI21_X1  g392(.A(KEYINPUT69), .B1(new_n261_), .B2(new_n336_), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n589_), .B(new_n592_), .C1(new_n593_), .C2(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n589_), .B1(new_n248_), .B2(new_n591_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT12), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n261_), .A2(new_n597_), .A3(new_n336_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n597_), .B1(new_n261_), .B2(new_n324_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n596_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G120gat), .B(G148gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT5), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G176gat), .B(G204gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n595_), .A2(new_n600_), .A3(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n595_), .A2(new_n600_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n604_), .B(KEYINPUT70), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n588_), .B(new_n605_), .C1(new_n606_), .C2(new_n607_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n595_), .A2(new_n600_), .A3(new_n604_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n607_), .B1(new_n595_), .B2(new_n600_), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT13), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n608_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n317_), .A2(new_n252_), .A3(new_n251_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n253_), .A2(new_n316_), .A3(new_n315_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G229gat), .A2(G233gat), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n264_), .A2(new_n317_), .A3(new_n265_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(new_n615_), .A3(new_n617_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G113gat), .B(G141gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G169gat), .B(G197gat), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n623_), .B(new_n624_), .Z(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n622_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT78), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n619_), .A2(new_n621_), .A3(new_n625_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n627_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n622_), .A2(KEYINPUT78), .A3(new_n626_), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n630_), .A2(KEYINPUT79), .A3(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(KEYINPUT79), .B1(new_n630_), .B2(new_n631_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n613_), .A2(new_n634_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n345_), .A2(new_n587_), .A3(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n636_), .A2(new_n311_), .A3(new_n464_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n637_), .B(KEYINPUT38), .Z(new_n638_));
  NAND2_X1  g437(.A1(new_n284_), .A2(new_n289_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n630_), .A2(new_n631_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n612_), .A2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT100), .ZN(new_n643_));
  INV_X1    g442(.A(new_n344_), .ZN(new_n644_));
  AND4_X1   g443(.A1(new_n587_), .A2(new_n639_), .A3(new_n643_), .A4(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT101), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n311_), .B1(new_n646_), .B2(new_n464_), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n638_), .A2(new_n647_), .ZN(G1324gat));
  INV_X1    g447(.A(new_n563_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n312_), .B1(new_n645_), .B2(new_n649_), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n650_), .B(KEYINPUT39), .Z(new_n651_));
  NAND3_X1  g450(.A1(new_n636_), .A2(new_n312_), .A3(new_n649_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT40), .Z(G1325gat));
  AOI21_X1  g453(.A(new_n508_), .B1(new_n646_), .B2(new_n586_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT102), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n656_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT41), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n657_), .A2(KEYINPUT41), .A3(new_n658_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n636_), .A2(new_n508_), .A3(new_n586_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n661_), .A2(new_n662_), .A3(new_n663_), .ZN(G1326gat));
  INV_X1    g463(.A(G22gat), .ZN(new_n665_));
  INV_X1    g464(.A(new_n434_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n646_), .B2(new_n666_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT42), .Z(new_n668_));
  NOR2_X1   g467(.A1(new_n434_), .A2(G22gat), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT103), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n636_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n668_), .A2(new_n671_), .ZN(G1327gat));
  NOR2_X1   g471(.A1(new_n639_), .A2(new_n644_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n434_), .A2(new_n584_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n464_), .ZN(new_n675_));
  OAI211_X1 g474(.A(new_n563_), .B(new_n675_), .C1(new_n432_), .C2(new_n433_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n586_), .B1(new_n674_), .B2(new_n676_), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n434_), .A2(new_n522_), .A3(new_n563_), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n635_), .B(new_n673_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n587_), .A2(KEYINPUT105), .A3(new_n635_), .A4(new_n673_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G29gat), .B1(new_n684_), .B2(new_n464_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n643_), .A2(new_n344_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n674_), .A2(new_n676_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n586_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n678_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n284_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n284_), .A2(new_n289_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(new_n692_), .B2(new_n292_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n690_), .A2(new_n693_), .A3(KEYINPUT43), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n695_), .B1(new_n587_), .B2(new_n294_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n687_), .B1(new_n694_), .B2(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT44), .B1(new_n697_), .B2(KEYINPUT104), .ZN(new_n698_));
  OAI21_X1  g497(.A(KEYINPUT43), .B1(new_n690_), .B2(new_n693_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n587_), .A2(new_n294_), .A3(new_n695_), .ZN(new_n700_));
  AOI211_X1 g499(.A(KEYINPUT104), .B(new_n686_), .C1(new_n699_), .C2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n686_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n703_));
  AOI22_X1  g502(.A1(new_n698_), .A2(new_n702_), .B1(KEYINPUT44), .B2(new_n703_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n464_), .A2(G29gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n685_), .B1(new_n704_), .B2(new_n705_), .ZN(G1328gat));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT46), .ZN(new_n708_));
  INV_X1    g507(.A(G36gat), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n681_), .A2(new_n682_), .A3(new_n709_), .A4(new_n649_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT45), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n710_), .B(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n563_), .B1(new_n703_), .B2(KEYINPUT44), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT104), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n714_), .B1(new_n703_), .B2(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n713_), .B1(new_n716_), .B2(new_n701_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n712_), .B1(new_n717_), .B2(G36gat), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n707_), .B(new_n708_), .C1(new_n718_), .C2(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n710_), .B(KEYINPUT45), .ZN(new_n721_));
  OAI211_X1 g520(.A(KEYINPUT44), .B(new_n687_), .C1(new_n694_), .C2(new_n696_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(new_n649_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n723_), .B1(new_n698_), .B2(new_n702_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n721_), .B1(new_n724_), .B2(new_n709_), .ZN(new_n725_));
  AOI21_X1  g524(.A(KEYINPUT107), .B1(new_n725_), .B2(KEYINPUT106), .ZN(new_n726_));
  OAI21_X1  g525(.A(KEYINPUT46), .B1(new_n718_), .B2(new_n707_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n720_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(G1329gat));
  NAND3_X1  g528(.A1(new_n704_), .A2(G43gat), .A3(new_n586_), .ZN(new_n730_));
  INV_X1    g529(.A(G43gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n731_), .B1(new_n683_), .B2(new_n689_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g533(.A(G50gat), .B1(new_n684_), .B2(new_n666_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n666_), .A2(G50gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n704_), .B2(new_n736_), .ZN(G1331gat));
  NOR2_X1   g536(.A1(new_n612_), .A2(new_n641_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n345_), .A2(new_n587_), .A3(new_n738_), .ZN(new_n739_));
  AOI211_X1 g538(.A(G57gat), .B(new_n675_), .C1(new_n739_), .C2(KEYINPUT108), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n740_), .B1(KEYINPUT108), .B2(new_n739_), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n344_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n587_), .A2(new_n639_), .A3(new_n613_), .A4(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(G57gat), .B1(new_n743_), .B2(new_n675_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n741_), .A2(new_n744_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT109), .ZN(G1332gat));
  OAI21_X1  g545(.A(G64gat), .B1(new_n743_), .B2(new_n563_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n747_), .B(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n649_), .A2(new_n295_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n749_), .B1(new_n739_), .B2(new_n750_), .ZN(G1333gat));
  OAI21_X1  g550(.A(G71gat), .B1(new_n743_), .B2(new_n689_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT49), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n689_), .A2(G71gat), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n753_), .B1(new_n739_), .B2(new_n754_), .ZN(G1334gat));
  OAI21_X1  g554(.A(G78gat), .B1(new_n743_), .B2(new_n434_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT50), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n434_), .A2(G78gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n739_), .B2(new_n758_), .ZN(G1335gat));
  NAND3_X1  g558(.A1(new_n587_), .A2(new_n673_), .A3(new_n738_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(new_n234_), .A3(new_n464_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n738_), .A2(new_n344_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n763_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n764_), .A2(new_n464_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n762_), .B1(new_n765_), .B2(new_n234_), .ZN(G1336gat));
  AOI21_X1  g565(.A(G92gat), .B1(new_n761_), .B2(new_n649_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n236_), .A2(new_n237_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n563_), .A2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n767_), .B1(new_n764_), .B2(new_n769_), .ZN(G1337gat));
  NAND3_X1  g569(.A1(new_n586_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772_));
  OAI22_X1  g571(.A1(new_n760_), .A2(new_n771_), .B1(KEYINPUT111), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n764_), .A2(new_n586_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n773_), .B1(new_n774_), .B2(G99gat), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n772_), .A2(KEYINPUT111), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n775_), .B(new_n776_), .Z(G1338gat));
  AOI21_X1  g576(.A(new_n213_), .B1(new_n764_), .B2(new_n666_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT52), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n760_), .A2(G106gat), .A3(new_n434_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  XOR2_X1   g580(.A(new_n781_), .B(KEYINPUT53), .Z(G1339gat));
  NOR4_X1   g581(.A1(new_n666_), .A2(new_n689_), .A3(new_n649_), .A4(new_n675_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n784_), .A2(KEYINPUT59), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT118), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT56), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n600_), .A2(KEYINPUT55), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n261_), .A2(new_n597_), .A3(new_n336_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n226_), .A2(new_n233_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n306_), .B1(new_n790_), .B2(new_n255_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n789_), .B1(new_n791_), .B2(new_n597_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(new_n793_), .A3(new_n596_), .ZN(new_n794_));
  OAI22_X1  g593(.A1(new_n598_), .A2(new_n599_), .B1(new_n261_), .B2(new_n336_), .ZN(new_n795_));
  AOI22_X1  g594(.A1(new_n788_), .A2(new_n794_), .B1(new_n589_), .B2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n787_), .B1(new_n796_), .B2(new_n607_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n607_), .A2(new_n787_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT114), .B1(new_n796_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n795_), .A2(new_n589_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n600_), .A2(KEYINPUT55), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n793_), .B1(new_n792_), .B2(new_n596_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n801_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(new_n805_), .A3(new_n798_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n797_), .A2(new_n800_), .A3(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n640_), .A2(new_n609_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n616_), .A2(new_n617_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n620_), .A2(new_n615_), .A3(new_n618_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n810_), .A2(new_n626_), .A3(new_n811_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n812_), .A2(new_n629_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  OAI211_X1 g615(.A(KEYINPUT115), .B(new_n813_), .C1(new_n609_), .C2(new_n610_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n692_), .B1(new_n809_), .B2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n786_), .B1(new_n820_), .B2(KEYINPUT57), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n818_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT57), .ZN(new_n823_));
  NOR4_X1   g622(.A1(new_n822_), .A2(new_n692_), .A3(KEYINPUT118), .A4(new_n823_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n821_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT58), .ZN(new_n827_));
  INV_X1    g626(.A(new_n607_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT56), .B1(new_n804_), .B2(new_n828_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n796_), .A2(new_n799_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n605_), .A2(new_n813_), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n826_), .B(new_n827_), .C1(new_n831_), .C2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n830_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n832_), .B1(new_n834_), .B2(new_n797_), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT58), .B1(new_n835_), .B2(KEYINPUT117), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n294_), .A2(new_n833_), .A3(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT116), .B1(new_n822_), .B2(new_n692_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n823_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n822_), .A2(KEYINPUT116), .A3(new_n692_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n837_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n825_), .B1(new_n841_), .B2(KEYINPUT119), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n843_), .B(new_n837_), .C1(new_n839_), .C2(new_n840_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n644_), .B1(new_n842_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT112), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n846_), .B1(new_n742_), .B2(new_n612_), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n742_), .A2(new_n846_), .A3(new_n612_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n693_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT113), .B1(new_n849_), .B2(KEYINPUT54), .ZN(new_n850_));
  OR2_X1    g649(.A1(new_n848_), .A2(new_n847_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT113), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n851_), .A2(new_n852_), .A3(new_n853_), .A4(new_n693_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n849_), .A2(KEYINPUT54), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n850_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n785_), .B1(new_n845_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n344_), .B1(new_n841_), .B2(new_n825_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n784_), .B1(new_n860_), .B2(new_n856_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n858_), .B1(new_n859_), .B2(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(G113gat), .B1(new_n862_), .B2(new_n634_), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n294_), .A2(new_n833_), .A3(new_n836_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n809_), .A2(new_n819_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n639_), .ZN(new_n866_));
  AOI21_X1  g665(.A(KEYINPUT57), .B1(new_n866_), .B2(KEYINPUT116), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT116), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n820_), .A2(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n864_), .B1(new_n867_), .B2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n824_), .ZN(new_n871_));
  OAI21_X1  g670(.A(KEYINPUT118), .B1(new_n866_), .B2(new_n823_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n644_), .B1(new_n870_), .B2(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n783_), .B1(new_n874_), .B2(new_n857_), .ZN(new_n875_));
  OR2_X1    g674(.A1(new_n640_), .A2(G113gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n863_), .B1(new_n875_), .B2(new_n876_), .ZN(G1340gat));
  INV_X1    g676(.A(G120gat), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n612_), .B1(new_n875_), .B2(KEYINPUT59), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n878_), .B1(new_n879_), .B2(new_n858_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n860_), .A2(new_n856_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n878_), .A2(KEYINPUT60), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n612_), .A2(KEYINPUT60), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n883_), .B1(new_n884_), .B2(new_n878_), .ZN(new_n885_));
  AND4_X1   g684(.A1(new_n881_), .A2(new_n882_), .A3(new_n783_), .A4(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n881_), .B1(new_n861_), .B2(new_n885_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(KEYINPUT121), .B1(new_n880_), .B2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n785_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n841_), .A2(KEYINPUT119), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n891_), .A2(new_n873_), .A3(new_n844_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n344_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n890_), .B1(new_n893_), .B2(new_n856_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n613_), .B1(new_n861_), .B2(new_n859_), .ZN(new_n895_));
  OAI21_X1  g694(.A(G120gat), .B1(new_n894_), .B2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n897_));
  INV_X1    g696(.A(new_n885_), .ZN(new_n898_));
  OAI21_X1  g697(.A(KEYINPUT120), .B1(new_n875_), .B2(new_n898_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n861_), .A2(new_n881_), .A3(new_n885_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n896_), .A2(new_n897_), .A3(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n889_), .A2(new_n902_), .ZN(G1341gat));
  OAI21_X1  g702(.A(G127gat), .B1(new_n862_), .B2(new_n344_), .ZN(new_n904_));
  OR2_X1    g703(.A1(new_n344_), .A2(G127gat), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n875_), .B2(new_n905_), .ZN(G1342gat));
  OAI21_X1  g705(.A(G134gat), .B1(new_n862_), .B2(new_n693_), .ZN(new_n907_));
  OR2_X1    g706(.A1(new_n639_), .A2(G134gat), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n875_), .B2(new_n908_), .ZN(G1343gat));
  NAND3_X1  g708(.A1(new_n666_), .A2(new_n464_), .A3(new_n563_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n882_), .A2(new_n689_), .A3(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(new_n640_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(KEYINPUT122), .B(G141gat), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n913_), .B(new_n914_), .ZN(G1344gat));
  NOR2_X1   g714(.A1(new_n912_), .A2(new_n612_), .ZN(new_n916_));
  XOR2_X1   g715(.A(new_n916_), .B(G148gat), .Z(G1345gat));
  NAND4_X1  g716(.A1(new_n882_), .A2(new_n689_), .A3(new_n644_), .A4(new_n911_), .ZN(new_n918_));
  OR2_X1    g717(.A1(new_n918_), .A2(KEYINPUT123), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(KEYINPUT123), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(KEYINPUT61), .B(G155gat), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n923_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n919_), .A2(new_n920_), .A3(new_n922_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(G1346gat));
  OAI21_X1  g725(.A(G162gat), .B1(new_n912_), .B2(new_n693_), .ZN(new_n927_));
  OR2_X1    g726(.A1(new_n639_), .A2(G162gat), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n927_), .B1(new_n912_), .B2(new_n928_), .ZN(G1347gat));
  NAND2_X1  g728(.A1(new_n649_), .A2(new_n522_), .ZN(new_n930_));
  AOI211_X1 g729(.A(new_n666_), .B(new_n930_), .C1(new_n893_), .C2(new_n856_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n931_), .A2(new_n492_), .A3(new_n641_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n930_), .A2(new_n666_), .ZN(new_n933_));
  OAI211_X1 g732(.A(new_n641_), .B(new_n933_), .C1(new_n845_), .C2(new_n857_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(G169gat), .ZN(new_n935_));
  XNOR2_X1  g734(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(new_n936_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n934_), .A2(G169gat), .A3(new_n938_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n932_), .A2(new_n937_), .A3(new_n939_), .ZN(G1348gat));
  AOI21_X1  g739(.A(new_n666_), .B1(new_n860_), .B2(new_n856_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n930_), .ZN(new_n942_));
  AND4_X1   g741(.A1(G176gat), .A2(new_n941_), .A3(new_n613_), .A4(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n931_), .A2(new_n613_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n943_), .B1(new_n944_), .B2(new_n491_), .ZN(G1349gat));
  NOR2_X1   g744(.A1(new_n930_), .A2(new_n344_), .ZN(new_n946_));
  AOI21_X1  g745(.A(G183gat), .B1(new_n941_), .B2(new_n946_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n344_), .A2(new_n476_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n947_), .B1(new_n931_), .B2(new_n948_), .ZN(G1350gat));
  NAND3_X1  g748(.A1(new_n931_), .A2(new_n477_), .A3(new_n692_), .ZN(new_n950_));
  OAI211_X1 g749(.A(new_n294_), .B(new_n933_), .C1(new_n845_), .C2(new_n857_), .ZN(new_n951_));
  INV_X1    g750(.A(KEYINPUT125), .ZN(new_n952_));
  AND3_X1   g751(.A1(new_n951_), .A2(new_n952_), .A3(G190gat), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n952_), .B1(new_n951_), .B2(G190gat), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n950_), .B1(new_n953_), .B2(new_n954_), .ZN(G1351gat));
  NAND2_X1  g754(.A1(new_n882_), .A2(new_n689_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n569_), .A2(new_n649_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n956_), .A2(new_n957_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n958_), .A2(new_n641_), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n959_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g759(.A1(new_n958_), .A2(new_n613_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n961_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g761(.A1(new_n958_), .A2(new_n644_), .ZN(new_n963_));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n964_));
  NOR2_X1   g763(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n965_));
  NAND3_X1  g764(.A1(new_n963_), .A2(new_n964_), .A3(new_n965_), .ZN(new_n966_));
  NOR3_X1   g765(.A1(new_n956_), .A2(new_n344_), .A3(new_n957_), .ZN(new_n967_));
  INV_X1    g766(.A(new_n965_), .ZN(new_n968_));
  OAI21_X1  g767(.A(KEYINPUT126), .B1(new_n967_), .B2(new_n968_), .ZN(new_n969_));
  XOR2_X1   g768(.A(KEYINPUT63), .B(G211gat), .Z(new_n970_));
  AOI22_X1  g769(.A1(new_n966_), .A2(new_n969_), .B1(new_n967_), .B2(new_n970_), .ZN(G1354gat));
  AOI21_X1  g770(.A(G218gat), .B1(new_n958_), .B2(new_n692_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n294_), .A2(G218gat), .ZN(new_n973_));
  XNOR2_X1  g772(.A(new_n973_), .B(KEYINPUT127), .ZN(new_n974_));
  AOI21_X1  g773(.A(new_n972_), .B1(new_n958_), .B2(new_n974_), .ZN(G1355gat));
endmodule


