//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n798_, new_n799_,
    new_n800_, new_n802_, new_n803_, new_n804_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n821_, new_n822_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n935_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n961_, new_n963_, new_n964_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n972_, new_n973_,
    new_n974_, new_n976_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_,
    new_n989_;
  INV_X1    g000(.A(KEYINPUT83), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT76), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT6), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND3_X1  g005(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n207_));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G106gat), .Z(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT10), .B(G99gat), .ZN(new_n209_));
  OAI211_X1 g008(.A(new_n206_), .B(new_n207_), .C1(new_n208_), .C2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n211_), .B1(G85gat), .B2(G92gat), .ZN(new_n212_));
  INV_X1    g011(.A(G92gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT65), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT65), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(G92gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n216_), .A3(G85gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT9), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT66), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n212_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(G92gat), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT9), .B1(new_n222_), .B2(G85gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT66), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n210_), .B1(new_n221_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT7), .ZN(new_n226_));
  INV_X1    g025(.A(G99gat), .ZN(new_n227_));
  INV_X1    g026(.A(G106gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n229_), .A2(new_n206_), .A3(new_n207_), .A4(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT8), .ZN(new_n232_));
  INV_X1    g031(.A(G85gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n233_), .A2(new_n213_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(G85gat), .A2(G92gat), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  AND3_X1   g035(.A1(new_n231_), .A2(new_n232_), .A3(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n232_), .B1(new_n231_), .B2(new_n236_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  XOR2_X1   g038(.A(G43gat), .B(G50gat), .Z(new_n240_));
  XNOR2_X1  g039(.A(G29gat), .B(G36gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  NOR3_X1   g041(.A1(new_n225_), .A2(new_n239_), .A3(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n244_), .B1(new_n225_), .B2(new_n239_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n231_), .A2(new_n236_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT8), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n231_), .A2(new_n232_), .A3(new_n236_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n217_), .A2(KEYINPUT66), .A3(new_n218_), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT66), .B1(new_n217_), .B2(new_n218_), .ZN(new_n251_));
  NOR3_X1   g050(.A1(new_n250_), .A2(new_n251_), .A3(new_n212_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n249_), .B(KEYINPUT67), .C1(new_n252_), .C2(new_n210_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n245_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT15), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n242_), .B(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n243_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n258_), .A2(KEYINPUT35), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT34), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n260_), .B1(new_n257_), .B2(KEYINPUT73), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n242_), .B(KEYINPUT15), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n262_), .B1(new_n245_), .B2(new_n253_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT73), .ZN(new_n264_));
  NOR4_X1   g063(.A1(new_n263_), .A2(new_n264_), .A3(KEYINPUT34), .A4(new_n243_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G232gat), .A2(G233gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NOR3_X1   g066(.A1(new_n261_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n268_));
  NOR3_X1   g067(.A1(new_n225_), .A2(new_n239_), .A3(new_n244_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n210_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n212_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n271_), .B1(new_n223_), .B2(KEYINPUT66), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n270_), .B1(new_n272_), .B2(new_n250_), .ZN(new_n273_));
  AOI21_X1  g072(.A(KEYINPUT67), .B1(new_n273_), .B2(new_n249_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n256_), .B1(new_n269_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n243_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(KEYINPUT73), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT34), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n257_), .A2(KEYINPUT73), .A3(new_n260_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n266_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n259_), .B1(new_n268_), .B2(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n267_), .B1(new_n261_), .B2(new_n265_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n278_), .A2(new_n266_), .A3(new_n279_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n282_), .A2(new_n283_), .A3(KEYINPUT35), .ZN(new_n284_));
  XOR2_X1   g083(.A(G190gat), .B(G218gat), .Z(new_n285_));
  XNOR2_X1  g084(.A(G134gat), .B(G162gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT36), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT74), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n281_), .A2(new_n284_), .A3(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n287_), .B(KEYINPUT36), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n293_), .B1(new_n281_), .B2(new_n284_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT75), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n291_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n282_), .A2(new_n283_), .A3(KEYINPUT35), .ZN(new_n297_));
  INV_X1    g096(.A(new_n259_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n298_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n292_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n300_), .A2(KEYINPUT75), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n203_), .B(KEYINPUT37), .C1(new_n296_), .C2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n300_), .A2(KEYINPUT75), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n281_), .A2(new_n284_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n305_), .A2(new_n295_), .A3(new_n292_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n304_), .A2(new_n306_), .A3(new_n291_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n203_), .B1(new_n307_), .B2(KEYINPUT37), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(KEYINPUT77), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT77), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n281_), .A2(new_n310_), .A3(new_n284_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(new_n292_), .A3(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT37), .ZN(new_n313_));
  AND3_X1   g112(.A1(new_n312_), .A2(new_n313_), .A3(new_n291_), .ZN(new_n314_));
  NOR3_X1   g113(.A1(new_n303_), .A2(new_n308_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(G57gat), .ZN(new_n316_));
  INV_X1    g115(.A(G64gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G57gat), .A2(G64gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n320_), .A2(KEYINPUT11), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G71gat), .B(G78gat), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n322_), .B1(KEYINPUT11), .B2(new_n320_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n320_), .A2(new_n322_), .A3(KEYINPUT11), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT79), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G231gat), .A2(G233gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(G15gat), .B(G22gat), .Z(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT78), .B(G1gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(G8gat), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n330_), .B1(new_n332_), .B2(KEYINPUT14), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G1gat), .B(G8gat), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n333_), .A2(new_n334_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n329_), .B(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G127gat), .B(G155gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G183gat), .B(G211gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT17), .ZN(new_n344_));
  OR2_X1    g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n344_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n338_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT82), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT81), .B1(new_n338_), .B2(new_n345_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n202_), .B1(new_n315_), .B2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT37), .B1(new_n296_), .B2(new_n301_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n293_), .B1(new_n305_), .B2(KEYINPUT77), .ZN(new_n354_));
  INV_X1    g153(.A(new_n305_), .ZN(new_n355_));
  AOI22_X1  g154(.A1(new_n354_), .A2(new_n311_), .B1(new_n355_), .B2(new_n290_), .ZN(new_n356_));
  AOI22_X1  g155(.A1(new_n353_), .A2(KEYINPUT76), .B1(new_n356_), .B2(new_n313_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n351_), .B1(new_n357_), .B2(new_n302_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT83), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n352_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT13), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT72), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT68), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n326_), .B1(new_n273_), .B2(new_n249_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n363_), .B1(new_n364_), .B2(KEYINPUT12), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT12), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n225_), .A2(new_n239_), .ZN(new_n367_));
  OAI211_X1 g166(.A(KEYINPUT68), .B(new_n366_), .C1(new_n367_), .C2(new_n326_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n365_), .A2(new_n368_), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n273_), .A2(new_n249_), .A3(new_n326_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n326_), .A2(new_n366_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n370_), .B1(new_n254_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G230gat), .A2(G233gat), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n369_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT69), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n369_), .A2(new_n372_), .A3(KEYINPUT69), .A4(new_n373_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n370_), .A2(new_n364_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n379_), .A2(new_n373_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  XOR2_X1   g180(.A(G176gat), .B(G204gat), .Z(new_n382_));
  XNOR2_X1  g181(.A(G120gat), .B(G148gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n385_));
  XOR2_X1   g184(.A(new_n384_), .B(new_n385_), .Z(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n378_), .A2(new_n381_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT71), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n380_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT71), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(new_n391_), .A3(new_n387_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n389_), .A2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n387_), .B1(new_n378_), .B2(new_n381_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n362_), .B1(new_n393_), .B2(new_n395_), .ZN(new_n396_));
  AOI211_X1 g195(.A(KEYINPUT72), .B(new_n394_), .C1(new_n389_), .C2(new_n392_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n361_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  AND4_X1   g197(.A1(new_n391_), .A2(new_n378_), .A3(new_n381_), .A4(new_n387_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n391_), .B1(new_n390_), .B2(new_n387_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n395_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT72), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n393_), .A2(new_n362_), .A3(new_n395_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(new_n403_), .A3(KEYINPUT13), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n398_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n337_), .A2(new_n242_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n242_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n408_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G229gat), .A2(G233gat), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT84), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT86), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT85), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n256_), .A2(new_n337_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n416_), .B1(new_n417_), .B2(new_n409_), .ZN(new_n418_));
  AOI21_X1  g217(.A(KEYINPUT85), .B1(new_n256_), .B2(new_n337_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n415_), .B1(new_n420_), .B2(new_n411_), .ZN(new_n421_));
  NOR4_X1   g220(.A1(new_n418_), .A2(KEYINPUT86), .A3(new_n412_), .A4(new_n419_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n414_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G113gat), .B(G141gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G169gat), .B(G197gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT87), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n423_), .A2(new_n428_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n427_), .B(new_n414_), .C1(new_n421_), .C2(new_n422_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n406_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G127gat), .B(G134gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G113gat), .B(G120gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT31), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT23), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n437_), .A2(G183gat), .A3(G190gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G183gat), .A2(G190gat), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT89), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n439_), .A2(new_n440_), .A3(KEYINPUT23), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n440_), .B1(new_n439_), .B2(KEYINPUT23), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n438_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT26), .B(G190gat), .ZN(new_n444_));
  INV_X1    g243(.A(G183gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT25), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT88), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n447_), .B1(new_n445_), .B2(KEYINPUT25), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT25), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(KEYINPUT88), .A3(G183gat), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n444_), .A2(new_n446_), .A3(new_n448_), .A4(new_n450_), .ZN(new_n451_));
  NOR3_X1   g250(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G169gat), .A2(G176gat), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n452_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n443_), .A2(new_n451_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n439_), .A2(KEYINPUT23), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n438_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n459_), .B1(G183gat), .B2(G190gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(KEYINPUT90), .A2(KEYINPUT22), .ZN(new_n461_));
  INV_X1    g260(.A(G176gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(G169gat), .A2(G176gat), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n463_), .A2(G169gat), .B1(new_n461_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n460_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n457_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT91), .B(G43gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(G71gat), .B(G99gat), .Z(new_n470_));
  NAND2_X1  g269(.A1(G227gat), .A2(G233gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT30), .B(G15gat), .ZN(new_n473_));
  XOR2_X1   g272(.A(new_n472_), .B(new_n473_), .Z(new_n474_));
  OR2_X1    g273(.A1(new_n469_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT92), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n469_), .A2(new_n474_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n476_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n436_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n481_), .B1(new_n479_), .B2(new_n436_), .ZN(new_n482_));
  XOR2_X1   g281(.A(new_n433_), .B(new_n434_), .Z(new_n483_));
  INV_X1    g282(.A(KEYINPUT3), .ZN(new_n484_));
  INV_X1    g283(.A(G141gat), .ZN(new_n485_));
  INV_X1    g284(.A(G148gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n484_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G141gat), .A2(G148gat), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT2), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n487_), .A2(new_n490_), .A3(new_n491_), .A4(new_n492_), .ZN(new_n493_));
  OR2_X1    g292(.A1(G155gat), .A2(G162gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G155gat), .A2(G162gat), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(KEYINPUT1), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT1), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n499_), .A2(G155gat), .A3(G162gat), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n498_), .A2(new_n500_), .A3(new_n494_), .ZN(new_n501_));
  XOR2_X1   g300(.A(G141gat), .B(G148gat), .Z(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n497_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT100), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n483_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  AOI22_X1  g305(.A1(new_n493_), .A2(new_n496_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n435_), .A2(new_n507_), .A3(KEYINPUT100), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n506_), .A2(KEYINPUT4), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G225gat), .A2(G233gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  OR3_X1    g310(.A1(new_n435_), .A2(new_n507_), .A3(KEYINPUT4), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n509_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n506_), .A2(new_n510_), .A3(new_n508_), .ZN(new_n514_));
  XOR2_X1   g313(.A(G1gat), .B(G29gat), .Z(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT101), .B(G85gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT0), .B(G57gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n513_), .A2(new_n514_), .A3(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n520_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n482_), .A2(new_n524_), .ZN(new_n525_));
  OR3_X1    g324(.A1(new_n504_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n526_));
  OAI21_X1  g325(.A(KEYINPUT28), .B1(new_n504_), .B2(KEYINPUT29), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G22gat), .B(G50gat), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n526_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n528_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(G211gat), .ZN(new_n532_));
  INV_X1    g331(.A(G218gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G211gat), .A2(G218gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G197gat), .B(G204gat), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT21), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n536_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(G204gat), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n540_), .A2(KEYINPUT95), .A3(G197gat), .ZN(new_n541_));
  INV_X1    g340(.A(G197gat), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n542_), .A2(G204gat), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(KEYINPUT95), .B1(new_n540_), .B2(G197gat), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n541_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n539_), .B1(new_n538_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT96), .ZN(new_n548_));
  INV_X1    g347(.A(new_n535_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(G211gat), .A2(G218gat), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n548_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n534_), .A2(KEYINPUT96), .A3(new_n535_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(new_n552_), .A3(KEYINPUT21), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n553_), .A2(new_n546_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT29), .ZN(new_n555_));
  OAI22_X1  g354(.A1(new_n547_), .A2(new_n554_), .B1(new_n507_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT93), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n557_), .B1(new_n547_), .B2(new_n554_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT94), .ZN(new_n559_));
  OAI21_X1  g358(.A(G228gat), .B1(new_n559_), .B2(G233gat), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n560_), .B1(new_n559_), .B2(G233gat), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n556_), .A2(new_n558_), .A3(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n504_), .A2(KEYINPUT29), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n540_), .A2(G197gat), .ZN(new_n565_));
  OAI21_X1  g364(.A(KEYINPUT21), .B1(new_n543_), .B2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n540_), .A2(KEYINPUT95), .A3(G197gat), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT95), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n568_), .B1(new_n542_), .B2(G204gat), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n567_), .B1(new_n569_), .B2(new_n543_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n536_), .B(new_n566_), .C1(new_n570_), .C2(KEYINPUT21), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n570_), .A2(KEYINPUT21), .A3(new_n551_), .A4(new_n552_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n564_), .B(new_n573_), .C1(new_n557_), .C2(new_n561_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n563_), .A2(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(G78gat), .B(G106gat), .Z(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n576_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n563_), .A2(new_n574_), .A3(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n531_), .A2(new_n577_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT98), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT97), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n579_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n577_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n575_), .A2(new_n582_), .A3(new_n576_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n531_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n581_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  AOI211_X1 g387(.A(KEYINPUT98), .B(new_n531_), .C1(new_n584_), .C2(new_n585_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n580_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G8gat), .B(G36gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(G92gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(KEYINPUT18), .B(G64gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G226gat), .A2(G233gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT19), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT22), .B(G169gat), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(new_n462_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n458_), .A2(KEYINPUT89), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n439_), .A2(new_n440_), .A3(KEYINPUT23), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n445_), .A2(KEYINPUT23), .ZN(new_n602_));
  AOI22_X1  g401(.A1(new_n600_), .A2(new_n601_), .B1(G190gat), .B2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(G183gat), .A2(G190gat), .ZN(new_n604_));
  OAI211_X1 g403(.A(new_n455_), .B(new_n599_), .C1(new_n603_), .C2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n444_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n449_), .A2(G183gat), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n446_), .A2(new_n607_), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n456_), .B(new_n459_), .C1(new_n606_), .C2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n605_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT103), .ZN(new_n611_));
  INV_X1    g410(.A(new_n573_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT103), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n605_), .A2(new_n613_), .A3(new_n609_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n611_), .A2(new_n612_), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT20), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n616_), .B1(new_n573_), .B2(new_n467_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n597_), .B1(new_n615_), .B2(new_n617_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n571_), .A2(new_n457_), .A3(new_n466_), .A4(new_n572_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT20), .ZN(new_n620_));
  AOI22_X1  g419(.A1(new_n605_), .A2(new_n609_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n620_), .A2(new_n621_), .A3(new_n596_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n594_), .B1(new_n618_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n594_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n620_), .A2(new_n621_), .A3(new_n597_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n605_), .A2(new_n571_), .A3(new_n572_), .A4(new_n609_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n596_), .B1(new_n617_), .B2(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n624_), .B1(new_n625_), .B2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n623_), .A2(KEYINPUT27), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT27), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n625_), .A2(new_n627_), .A3(new_n624_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n573_), .A2(new_n467_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n626_), .A2(new_n632_), .A3(KEYINPUT20), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(new_n597_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n610_), .A2(new_n573_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n635_), .A2(KEYINPUT20), .A3(new_n596_), .A4(new_n619_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n594_), .B1(new_n634_), .B2(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n630_), .B1(new_n631_), .B2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n629_), .A2(new_n638_), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n525_), .A2(new_n590_), .A3(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n629_), .A2(new_n524_), .A3(new_n638_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n590_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n644_), .B1(new_n631_), .B2(new_n637_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n521_), .A2(KEYINPUT33), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT33), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n513_), .A2(new_n647_), .A3(new_n514_), .A4(new_n520_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n506_), .A2(KEYINPUT102), .A3(new_n508_), .ZN(new_n650_));
  AOI21_X1  g449(.A(KEYINPUT102), .B1(new_n506_), .B2(new_n508_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n511_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n509_), .A2(new_n510_), .A3(new_n512_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(new_n519_), .A3(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n634_), .A2(new_n594_), .A3(new_n636_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n628_), .A2(new_n655_), .A3(KEYINPUT99), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n645_), .A2(new_n649_), .A3(new_n654_), .A4(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n624_), .A2(KEYINPUT32), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n658_), .B1(new_n625_), .B2(new_n627_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n618_), .A2(new_n622_), .ZN(new_n660_));
  OAI221_X1 g459(.A(new_n659_), .B1(new_n522_), .B2(new_n523_), .C1(new_n660_), .C2(new_n658_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n657_), .A2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n578_), .B1(new_n563_), .B2(new_n574_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(new_n582_), .B2(new_n579_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n585_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n587_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT98), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n586_), .A2(new_n581_), .A3(new_n587_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n662_), .A2(new_n669_), .A3(new_n580_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n482_), .B1(new_n643_), .B2(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n640_), .B1(new_n671_), .B2(KEYINPUT104), .ZN(new_n672_));
  INV_X1    g471(.A(new_n482_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n662_), .A2(new_n669_), .A3(new_n580_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n641_), .B1(new_n669_), .B2(new_n580_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n673_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n672_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n432_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n360_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n524_), .A2(new_n331_), .ZN(new_n684_));
  AOI21_X1  g483(.A(KEYINPUT38), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n356_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n679_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n431_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n405_), .A2(new_n690_), .A3(new_n351_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n524_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n685_), .B1(G1gat), .B2(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n683_), .A2(KEYINPUT38), .A3(new_n684_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n697_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n695_), .A2(new_n698_), .A3(new_n699_), .ZN(G1324gat));
  INV_X1    g499(.A(new_n639_), .ZN(new_n701_));
  OR3_X1    g500(.A1(new_n682_), .A2(G8gat), .A3(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n689_), .A2(new_n639_), .A3(new_n691_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(G8gat), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(new_n705_), .A3(KEYINPUT39), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT39), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n703_), .A2(new_n707_), .A3(G8gat), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n705_), .B1(new_n704_), .B2(KEYINPUT39), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n702_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT40), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  OAI211_X1 g512(.A(KEYINPUT40), .B(new_n702_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1325gat));
  NAND2_X1  g514(.A1(new_n692_), .A2(new_n482_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(G15gat), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT41), .ZN(new_n718_));
  OR3_X1    g517(.A1(new_n682_), .A2(G15gat), .A3(new_n673_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT41), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n716_), .A2(new_n720_), .A3(G15gat), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n718_), .A2(new_n719_), .A3(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT108), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n718_), .A2(new_n719_), .A3(KEYINPUT108), .A4(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1326gat));
  NAND2_X1  g525(.A1(new_n692_), .A2(new_n590_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(G22gat), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT42), .ZN(new_n729_));
  INV_X1    g528(.A(new_n590_), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n730_), .A2(G22gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n729_), .B1(new_n682_), .B2(new_n731_), .ZN(G1327gat));
  INV_X1    g531(.A(new_n351_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n733_), .A2(new_n686_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n681_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(G29gat), .B1(new_n736_), .B2(new_n693_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n353_), .A2(KEYINPUT76), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n356_), .A2(new_n313_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n738_), .A2(new_n679_), .A3(new_n302_), .A4(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT43), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n357_), .A2(new_n742_), .A3(new_n679_), .A4(new_n302_), .ZN(new_n743_));
  AOI211_X1 g542(.A(new_n733_), .B(new_n432_), .C1(new_n741_), .C2(new_n743_), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n744_), .A2(KEYINPUT44), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n745_), .A2(G29gat), .A3(new_n693_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(KEYINPUT44), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n737_), .B1(new_n746_), .B2(new_n747_), .ZN(G1328gat));
  INV_X1    g547(.A(new_n747_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n639_), .B1(new_n744_), .B2(KEYINPUT44), .ZN(new_n750_));
  OAI21_X1  g549(.A(G36gat), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n701_), .A2(G36gat), .ZN(new_n752_));
  OR3_X1    g551(.A1(new_n735_), .A2(KEYINPUT45), .A3(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT45), .B1(new_n735_), .B2(new_n752_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n751_), .A2(new_n755_), .A3(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n751_), .B2(new_n755_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1329gat));
  INV_X1    g558(.A(G43gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n760_), .B1(new_n735_), .B2(new_n673_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  OAI211_X1 g562(.A(KEYINPUT110), .B(new_n760_), .C1(new_n735_), .C2(new_n673_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  OAI211_X1 g564(.A(G43gat), .B(new_n482_), .C1(new_n744_), .C2(KEYINPUT44), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n749_), .B2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT47), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT47), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n765_), .B(new_n769_), .C1(new_n749_), .C2(new_n766_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(G1330gat));
  OR3_X1    g570(.A1(new_n735_), .A2(G50gat), .A3(new_n730_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n745_), .A2(new_n590_), .A3(new_n747_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n773_), .B1(new_n774_), .B2(G50gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n590_), .B1(new_n744_), .B2(KEYINPUT44), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n773_), .B(G50gat), .C1(new_n749_), .C2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n772_), .B1(new_n775_), .B2(new_n778_), .ZN(G1331gat));
  NAND3_X1  g578(.A1(new_n352_), .A2(new_n359_), .A3(new_n405_), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n780_), .A2(KEYINPUT112), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(KEYINPUT112), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n680_), .A2(new_n431_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n781_), .A2(new_n693_), .A3(new_n782_), .A4(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n784_), .A2(KEYINPUT113), .A3(new_n316_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n405_), .A2(new_n690_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n786_), .A2(new_n351_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n689_), .A2(G57gat), .A3(new_n693_), .A4(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n785_), .A2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT113), .B1(new_n784_), .B2(new_n316_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n789_), .A2(new_n790_), .ZN(G1332gat));
  NAND2_X1  g590(.A1(new_n689_), .A2(new_n787_), .ZN(new_n792_));
  OAI21_X1  g591(.A(G64gat), .B1(new_n792_), .B2(new_n701_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT48), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n781_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n639_), .A2(new_n317_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n794_), .B1(new_n795_), .B2(new_n796_), .ZN(G1333gat));
  OAI21_X1  g596(.A(G71gat), .B1(new_n792_), .B2(new_n673_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT49), .ZN(new_n799_));
  OR2_X1    g598(.A1(new_n673_), .A2(G71gat), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n799_), .B1(new_n795_), .B2(new_n800_), .ZN(G1334gat));
  OAI21_X1  g600(.A(G78gat), .B1(new_n792_), .B2(new_n730_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT50), .ZN(new_n803_));
  OR2_X1    g602(.A1(new_n730_), .A2(G78gat), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n803_), .B1(new_n795_), .B2(new_n804_), .ZN(G1335gat));
  NAND2_X1  g604(.A1(new_n741_), .A2(new_n743_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n402_), .A2(KEYINPUT13), .A3(new_n403_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT13), .B1(new_n402_), .B2(new_n403_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n690_), .B(new_n351_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n405_), .A2(KEYINPUT114), .A3(new_n690_), .A4(new_n351_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n806_), .A2(new_n813_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(KEYINPUT115), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n524_), .A2(new_n233_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n786_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n680_), .A2(new_n686_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n693_), .A4(new_n351_), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n815_), .A2(new_n816_), .B1(new_n233_), .B2(new_n819_), .ZN(G1336gat));
  AND2_X1   g619(.A1(new_n639_), .A2(new_n222_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n817_), .A2(new_n818_), .A3(new_n639_), .A4(new_n351_), .ZN(new_n822_));
  AOI22_X1  g621(.A1(new_n815_), .A2(new_n821_), .B1(new_n213_), .B2(new_n822_), .ZN(G1337gat));
  AOI21_X1  g622(.A(new_n227_), .B1(new_n814_), .B2(new_n482_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n673_), .A2(new_n209_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n817_), .A2(new_n818_), .A3(new_n351_), .A4(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  OAI22_X1  g626(.A1(new_n824_), .A2(new_n827_), .B1(KEYINPUT116), .B2(KEYINPUT51), .ZN(new_n828_));
  NAND2_X1  g627(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n828_), .B(new_n829_), .ZN(G1338gat));
  NOR2_X1   g629(.A1(new_n730_), .A2(new_n208_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n817_), .A2(new_n818_), .A3(new_n351_), .A4(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n806_), .A2(new_n590_), .A3(new_n813_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(KEYINPUT117), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n806_), .A2(new_n813_), .A3(new_n836_), .A4(new_n590_), .ZN(new_n837_));
  AND4_X1   g636(.A1(new_n833_), .A2(new_n835_), .A3(G106gat), .A4(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n228_), .B1(new_n834_), .B2(KEYINPUT117), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n833_), .B1(new_n839_), .B2(new_n837_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n832_), .B1(new_n838_), .B2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT53), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n843_), .B(new_n832_), .C1(new_n838_), .C2(new_n840_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n844_), .ZN(G1339gat));
  NOR3_X1   g644(.A1(new_n673_), .A2(new_n590_), .A3(new_n524_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n420_), .A2(new_n412_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n426_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n848_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n847_), .A2(KEYINPUT119), .A3(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n847_), .A2(new_n849_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT119), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n850_), .B(new_n853_), .C1(new_n423_), .C2(new_n426_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  OAI211_X1 g654(.A(KEYINPUT120), .B(new_n855_), .C1(new_n396_), .C2(new_n397_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n431_), .B1(new_n400_), .B2(new_n399_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(KEYINPUT55), .B1(new_n376_), .B2(new_n377_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n369_), .A2(new_n372_), .A3(KEYINPUT55), .A4(new_n373_), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n369_), .A2(new_n372_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n862_), .B2(new_n373_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n386_), .B1(new_n860_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT56), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  OAI211_X1 g665(.A(KEYINPUT56), .B(new_n386_), .C1(new_n860_), .C2(new_n863_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n393_), .A2(KEYINPUT118), .A3(new_n431_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n859_), .A2(new_n868_), .A3(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n856_), .A2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n402_), .A2(new_n403_), .ZN(new_n872_));
  AOI21_X1  g671(.A(KEYINPUT120), .B1(new_n872_), .B2(new_n855_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n686_), .B1(new_n871_), .B2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n875_));
  AND3_X1   g674(.A1(new_n868_), .A2(new_n393_), .A3(new_n855_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT58), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n876_), .B(new_n877_), .ZN(new_n878_));
  AOI22_X1  g677(.A1(new_n874_), .A2(new_n875_), .B1(new_n315_), .B2(new_n878_), .ZN(new_n879_));
  OAI211_X1 g678(.A(KEYINPUT57), .B(new_n686_), .C1(new_n871_), .C2(new_n873_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n733_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n398_), .A2(new_n690_), .A3(new_n404_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n358_), .B2(new_n883_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n738_), .A2(new_n302_), .A3(new_n739_), .ZN(new_n885_));
  AND4_X1   g684(.A1(new_n882_), .A2(new_n885_), .A3(new_n883_), .A4(new_n733_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n884_), .A2(new_n886_), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n701_), .B(new_n846_), .C1(new_n881_), .C2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(KEYINPUT59), .ZN(new_n889_));
  OR2_X1    g688(.A1(new_n876_), .A2(KEYINPUT58), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n876_), .A2(KEYINPUT58), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n357_), .A2(new_n890_), .A3(new_n302_), .A4(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n854_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n893_));
  AOI22_X1  g692(.A1(new_n857_), .A2(new_n858_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n894_));
  AOI22_X1  g693(.A1(new_n893_), .A2(KEYINPUT120), .B1(new_n869_), .B2(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n855_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n356_), .B1(new_n895_), .B2(new_n898_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n892_), .B1(new_n899_), .B2(KEYINPUT57), .ZN(new_n900_));
  INV_X1    g699(.A(new_n880_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n351_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n885_), .A2(new_n883_), .A3(new_n733_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(KEYINPUT54), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n905_), .A2(new_n906_), .A3(new_n701_), .A4(new_n846_), .ZN(new_n907_));
  AND4_X1   g706(.A1(G113gat), .A2(new_n889_), .A3(new_n431_), .A4(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n888_), .ZN(new_n909_));
  AOI21_X1  g708(.A(G113gat), .B1(new_n909_), .B2(new_n431_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n908_), .A2(new_n910_), .ZN(G1340gat));
  INV_X1    g710(.A(G120gat), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(KEYINPUT60), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n406_), .B2(KEYINPUT60), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT121), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n913_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n916_));
  OAI211_X1 g715(.A(new_n909_), .B(new_n916_), .C1(new_n915_), .C2(new_n914_), .ZN(new_n917_));
  AND3_X1   g716(.A1(new_n889_), .A2(new_n907_), .A3(new_n405_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n918_), .B2(new_n912_), .ZN(G1341gat));
  NAND4_X1  g718(.A1(new_n889_), .A2(new_n907_), .A3(G127gat), .A4(new_n733_), .ZN(new_n920_));
  INV_X1    g719(.A(G127gat), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n921_), .B1(new_n888_), .B2(new_n351_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT122), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  OAI211_X1 g723(.A(KEYINPUT122), .B(new_n921_), .C1(new_n888_), .C2(new_n351_), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n920_), .A2(new_n924_), .A3(new_n925_), .ZN(G1342gat));
  AND4_X1   g725(.A1(G134gat), .A2(new_n889_), .A3(new_n315_), .A4(new_n907_), .ZN(new_n927_));
  AOI21_X1  g726(.A(G134gat), .B1(new_n909_), .B2(new_n356_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n927_), .A2(new_n928_), .ZN(G1343gat));
  NAND2_X1  g728(.A1(new_n673_), .A2(new_n590_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n930_), .A2(new_n524_), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n701_), .B(new_n931_), .C1(new_n881_), .C2(new_n887_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n932_), .A2(new_n690_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(new_n485_), .ZN(G1344gat));
  NOR2_X1   g733(.A1(new_n932_), .A2(new_n406_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(new_n486_), .ZN(G1345gat));
  OAI21_X1  g735(.A(KEYINPUT123), .B1(new_n932_), .B2(new_n351_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(KEYINPUT61), .B(G155gat), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n639_), .B1(new_n902_), .B2(new_n904_), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT123), .ZN(new_n940_));
  NAND4_X1  g739(.A1(new_n939_), .A2(new_n940_), .A3(new_n733_), .A4(new_n931_), .ZN(new_n941_));
  AND3_X1   g740(.A1(new_n937_), .A2(new_n938_), .A3(new_n941_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n938_), .B1(new_n937_), .B2(new_n941_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n942_), .A2(new_n943_), .ZN(G1346gat));
  INV_X1    g743(.A(new_n932_), .ZN(new_n945_));
  AOI21_X1  g744(.A(G162gat), .B1(new_n945_), .B2(new_n356_), .ZN(new_n946_));
  INV_X1    g745(.A(G162gat), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n885_), .A2(new_n947_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(KEYINPUT124), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n946_), .B1(new_n945_), .B2(new_n949_), .ZN(G1347gat));
  NAND3_X1  g749(.A1(new_n730_), .A2(new_n482_), .A3(new_n524_), .ZN(new_n951_));
  INV_X1    g750(.A(new_n951_), .ZN(new_n952_));
  OAI211_X1 g751(.A(new_n639_), .B(new_n952_), .C1(new_n881_), .C2(new_n887_), .ZN(new_n953_));
  OAI21_X1  g752(.A(G169gat), .B1(new_n953_), .B2(new_n690_), .ZN(new_n954_));
  INV_X1    g753(.A(KEYINPUT62), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n954_), .A2(new_n955_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n701_), .B1(new_n902_), .B2(new_n904_), .ZN(new_n957_));
  NAND4_X1  g756(.A1(new_n957_), .A2(new_n431_), .A3(new_n598_), .A4(new_n952_), .ZN(new_n958_));
  OAI211_X1 g757(.A(KEYINPUT62), .B(G169gat), .C1(new_n953_), .C2(new_n690_), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n956_), .A2(new_n958_), .A3(new_n959_), .ZN(G1348gat));
  NOR2_X1   g759(.A1(new_n953_), .A2(new_n406_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n961_), .B(new_n462_), .ZN(G1349gat));
  NOR2_X1   g761(.A1(new_n953_), .A2(new_n351_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n963_), .A2(G183gat), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n964_), .B1(new_n608_), .B2(new_n963_), .ZN(G1350gat));
  NAND3_X1  g764(.A1(new_n957_), .A2(new_n952_), .A3(new_n315_), .ZN(new_n966_));
  AOI21_X1  g765(.A(KEYINPUT125), .B1(new_n966_), .B2(G190gat), .ZN(new_n967_));
  OAI211_X1 g766(.A(KEYINPUT125), .B(G190gat), .C1(new_n953_), .C2(new_n885_), .ZN(new_n968_));
  INV_X1    g767(.A(new_n968_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n356_), .A2(new_n444_), .ZN(new_n970_));
  OAI22_X1  g769(.A1(new_n967_), .A2(new_n969_), .B1(new_n953_), .B2(new_n970_), .ZN(G1351gat));
  NOR2_X1   g770(.A1(new_n930_), .A2(new_n693_), .ZN(new_n972_));
  OAI211_X1 g771(.A(new_n639_), .B(new_n972_), .C1(new_n881_), .C2(new_n887_), .ZN(new_n973_));
  NOR2_X1   g772(.A1(new_n973_), .A2(new_n690_), .ZN(new_n974_));
  XNOR2_X1  g773(.A(new_n974_), .B(new_n542_), .ZN(G1352gat));
  NOR2_X1   g774(.A1(new_n973_), .A2(new_n406_), .ZN(new_n976_));
  XNOR2_X1  g775(.A(new_n976_), .B(new_n540_), .ZN(G1353gat));
  NOR2_X1   g776(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n978_));
  AND2_X1   g777(.A1(new_n978_), .A2(KEYINPUT126), .ZN(new_n979_));
  AOI211_X1 g778(.A(new_n979_), .B(new_n351_), .C1(KEYINPUT63), .C2(G211gat), .ZN(new_n980_));
  NAND3_X1  g779(.A1(new_n957_), .A2(new_n972_), .A3(new_n980_), .ZN(new_n981_));
  NOR2_X1   g780(.A1(new_n978_), .A2(KEYINPUT126), .ZN(new_n982_));
  XNOR2_X1  g781(.A(new_n981_), .B(new_n982_), .ZN(G1354gat));
  OAI21_X1  g782(.A(new_n533_), .B1(new_n973_), .B2(new_n686_), .ZN(new_n984_));
  NAND4_X1  g783(.A1(new_n957_), .A2(G218gat), .A3(new_n315_), .A4(new_n972_), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n984_), .A2(new_n985_), .ZN(new_n986_));
  NAND2_X1  g785(.A1(new_n986_), .A2(KEYINPUT127), .ZN(new_n987_));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n988_));
  NAND3_X1  g787(.A1(new_n984_), .A2(new_n985_), .A3(new_n988_), .ZN(new_n989_));
  NAND2_X1  g788(.A1(new_n987_), .A2(new_n989_), .ZN(G1355gat));
endmodule


