//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1 1 0 0 1 0 0 0 1 1 1 0 0 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0 0 0 1 1 1 0 1 0 1 1 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n780_, new_n781_, new_n782_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_, new_n945_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n955_, new_n956_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n967_, new_n968_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n976_,
    new_n977_;
  INV_X1    g000(.A(KEYINPUT38), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G230gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT68), .B(KEYINPUT12), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT6), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n208_), .A2(G99gat), .A3(G106gat), .ZN(new_n209_));
  AND2_X1   g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT7), .ZN(new_n211_));
  INV_X1    g010(.A(G99gat), .ZN(new_n212_));
  INV_X1    g011(.A(G106gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n205_), .B1(new_n210_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n207_), .A2(new_n209_), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n218_), .A2(KEYINPUT64), .A3(new_n214_), .A4(new_n215_), .ZN(new_n219_));
  OR2_X1    g018(.A1(G85gat), .A2(G92gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n217_), .A2(new_n219_), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT8), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  OR2_X1    g025(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n213_), .A3(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n220_), .A2(KEYINPUT9), .A3(new_n221_), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n221_), .A2(KEYINPUT9), .ZN(new_n231_));
  AND4_X1   g030(.A1(new_n218_), .A2(new_n229_), .A3(new_n230_), .A4(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n218_), .A2(KEYINPUT65), .ZN(new_n233_));
  INV_X1    g032(.A(new_n215_), .ZN(new_n234_));
  NOR3_X1   g033(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT66), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n214_), .A2(new_n237_), .A3(new_n215_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n207_), .A2(new_n209_), .A3(new_n239_), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n233_), .A2(new_n236_), .A3(new_n238_), .A4(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n222_), .A2(new_n225_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n232_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n226_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G57gat), .B(G64gat), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n245_), .A2(KEYINPUT11), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(KEYINPUT11), .ZN(new_n247_));
  XOR2_X1   g046(.A(G71gat), .B(G78gat), .Z(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n247_), .A2(new_n248_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n204_), .B1(new_n244_), .B2(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n251_), .B1(new_n226_), .B2(new_n243_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n254_), .A2(KEYINPUT67), .A3(KEYINPUT12), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(KEYINPUT67), .B1(new_n254_), .B2(KEYINPUT12), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n203_), .B(new_n256_), .C1(new_n258_), .C2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n203_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n244_), .A2(new_n252_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n261_), .B1(new_n262_), .B2(new_n254_), .ZN(new_n263_));
  XOR2_X1   g062(.A(G120gat), .B(G148gat), .Z(new_n264_));
  XNOR2_X1  g063(.A(G176gat), .B(G204gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n267_));
  XOR2_X1   g066(.A(new_n266_), .B(new_n267_), .Z(new_n268_));
  NAND3_X1  g067(.A1(new_n260_), .A2(new_n263_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n268_), .B1(new_n260_), .B2(new_n263_), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT13), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT71), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n274_), .B(KEYINPUT13), .C1(new_n270_), .C2(new_n271_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n260_), .A2(new_n263_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n268_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT13), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(new_n280_), .A3(new_n269_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT70), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n279_), .A2(new_n283_), .A3(new_n280_), .A4(new_n269_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n276_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT76), .B(G15gat), .ZN(new_n287_));
  INV_X1    g086(.A(G22gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(G1gat), .B(G8gat), .Z(new_n290_));
  INV_X1    g089(.A(G1gat), .ZN(new_n291_));
  INV_X1    g090(.A(G8gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT14), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  AND3_X1   g092(.A1(new_n289_), .A2(new_n290_), .A3(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n290_), .B1(new_n289_), .B2(new_n293_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(new_n252_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G231gat), .A2(G233gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G127gat), .B(G155gat), .Z(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G183gat), .B(G211gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT17), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n299_), .A2(new_n305_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n304_), .A2(KEYINPUT17), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n299_), .A2(new_n305_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G190gat), .B(G218gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G134gat), .B(G162gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n313_), .A2(KEYINPUT36), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G232gat), .A2(G233gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT34), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n316_), .A2(KEYINPUT35), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G29gat), .B(G36gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G43gat), .B(G50gat), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n319_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n226_), .A2(new_n243_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT73), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n226_), .A2(new_n243_), .A3(KEYINPUT73), .A4(new_n322_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n317_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n320_), .A2(KEYINPUT15), .A3(new_n321_), .ZN(new_n328_));
  AOI21_X1  g127(.A(KEYINPUT15), .B1(new_n320_), .B2(new_n321_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n241_), .A2(new_n242_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n232_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n218_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n222_), .B1(new_n334_), .B2(new_n205_), .ZN(new_n335_));
  AOI21_X1  g134(.A(KEYINPUT8), .B1(new_n335_), .B2(new_n219_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n330_), .B1(new_n333_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n244_), .A2(KEYINPUT72), .A3(new_n330_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n316_), .A2(KEYINPUT35), .ZN(new_n342_));
  AND3_X1   g141(.A1(new_n327_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n342_), .B1(new_n327_), .B2(new_n341_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n314_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT74), .B1(new_n343_), .B2(new_n344_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n313_), .A2(KEYINPUT36), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n345_), .A2(new_n346_), .A3(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT75), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT37), .ZN(new_n351_));
  OAI221_X1 g150(.A(KEYINPUT74), .B1(new_n347_), .B2(new_n314_), .C1(new_n343_), .C2(new_n344_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n349_), .A2(new_n350_), .A3(new_n351_), .A4(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n349_), .A2(new_n352_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(KEYINPUT75), .A2(KEYINPUT37), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(KEYINPUT75), .A2(KEYINPUT37), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n354_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n286_), .A2(new_n310_), .A3(new_n353_), .A4(new_n358_), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n359_), .A2(KEYINPUT78), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(KEYINPUT78), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n320_), .A2(new_n321_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n362_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n289_), .A2(new_n293_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n290_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n289_), .A2(new_n290_), .A3(new_n293_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(new_n367_), .A3(new_n322_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n363_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT79), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n363_), .A2(new_n368_), .A3(KEYINPUT79), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n371_), .A2(G229gat), .A3(G233gat), .A4(new_n372_), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n328_), .A2(new_n329_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n368_), .B1(new_n296_), .B2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G229gat), .A2(G233gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT80), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n375_), .A2(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G113gat), .B(G141gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT81), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G169gat), .B(G197gat), .ZN(new_n382_));
  XOR2_X1   g181(.A(new_n381_), .B(new_n382_), .Z(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n373_), .A2(new_n379_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n384_), .B1(new_n373_), .B2(new_n379_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT82), .ZN(new_n388_));
  OR3_X1    g187(.A1(new_n386_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n388_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(G183gat), .ZN(new_n393_));
  INV_X1    g192(.A(G190gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G183gat), .A2(G190gat), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT23), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT85), .B(KEYINPUT23), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n395_), .B(new_n398_), .C1(new_n399_), .C2(new_n396_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT88), .ZN(new_n401_));
  INV_X1    g200(.A(new_n396_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT85), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n403_), .A2(KEYINPUT23), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n397_), .A2(KEYINPUT85), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n402_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT88), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n406_), .A2(new_n407_), .A3(new_n395_), .A4(new_n398_), .ZN(new_n408_));
  INV_X1    g207(.A(G169gat), .ZN(new_n409_));
  INV_X1    g208(.A(G176gat), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n409_), .A2(KEYINPUT87), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT86), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT22), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT22), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(G169gat), .ZN(new_n416_));
  AOI22_X1  g215(.A1(new_n412_), .A2(new_n414_), .B1(new_n416_), .B2(KEYINPUT87), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n415_), .A2(KEYINPUT86), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT87), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(G169gat), .ZN(new_n420_));
  AOI21_X1  g219(.A(G176gat), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n411_), .B1(new_n417_), .B2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n401_), .A2(new_n408_), .A3(new_n422_), .ZN(new_n423_));
  NOR3_X1   g222(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n396_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n396_), .A2(KEYINPUT23), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n424_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT24), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n429_), .B1(G169gat), .B2(G176gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n409_), .A2(new_n410_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n430_), .A2(KEYINPUT84), .A3(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT25), .B(G183gat), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT83), .B1(new_n394_), .B2(KEYINPUT26), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT26), .B(G190gat), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n433_), .B(new_n434_), .C1(new_n435_), .C2(KEYINPUT83), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n430_), .A2(new_n431_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT84), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n428_), .A2(new_n432_), .A3(new_n436_), .A4(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n423_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G227gat), .A2(G233gat), .ZN(new_n442_));
  INV_X1    g241(.A(G71gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(G99gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n441_), .B(new_n445_), .ZN(new_n446_));
  XOR2_X1   g245(.A(G127gat), .B(G134gat), .Z(new_n447_));
  XOR2_X1   g246(.A(G113gat), .B(G120gat), .Z(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n446_), .A2(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n446_), .A2(new_n449_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G15gat), .B(G43gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(KEYINPUT89), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT30), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT31), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  OR3_X1    g255(.A1(new_n450_), .A2(new_n451_), .A3(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n456_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G22gat), .B(G50gat), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT28), .ZN(new_n462_));
  INV_X1    g261(.A(G141gat), .ZN(new_n463_));
  INV_X1    g262(.A(G148gat), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n463_), .A2(new_n464_), .A3(KEYINPUT3), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT3), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n466_), .B1(G141gat), .B2(G148gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  AND3_X1   g267(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n469_));
  AOI21_X1  g268(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n468_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT92), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n468_), .A2(new_n471_), .A3(KEYINPUT92), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  OR2_X1    g275(.A1(G155gat), .A2(G162gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G155gat), .A2(G162gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT90), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n481_), .B1(new_n478_), .B2(KEYINPUT1), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT1), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n483_), .A2(KEYINPUT90), .A3(G155gat), .A4(G162gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n478_), .A2(KEYINPUT1), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n482_), .A2(new_n484_), .A3(new_n485_), .A4(new_n477_), .ZN(new_n486_));
  XOR2_X1   g285(.A(G141gat), .B(G148gat), .Z(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT91), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT91), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n486_), .A2(new_n490_), .A3(new_n487_), .ZN(new_n491_));
  AOI22_X1  g290(.A1(new_n476_), .A2(new_n480_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT29), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n462_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n486_), .A2(new_n490_), .A3(new_n487_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n490_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n479_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n498_));
  NOR4_X1   g297(.A1(new_n497_), .A2(new_n498_), .A3(KEYINPUT28), .A4(KEYINPUT29), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n461_), .B1(new_n494_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n489_), .A2(new_n491_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n475_), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT92), .B1(new_n468_), .B2(new_n471_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n480_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n501_), .A2(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT28), .B1(new_n505_), .B2(KEYINPUT29), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n492_), .A2(new_n462_), .A3(new_n493_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n461_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n506_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n500_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(G228gat), .ZN(new_n511_));
  INV_X1    g310(.A(G233gat), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(KEYINPUT96), .B(KEYINPUT29), .Z(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n515_), .B1(new_n501_), .B2(new_n504_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT21), .ZN(new_n517_));
  INV_X1    g316(.A(G218gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(G211gat), .ZN(new_n519_));
  INV_X1    g318(.A(G211gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(G218gat), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n517_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT94), .ZN(new_n523_));
  AND2_X1   g322(.A1(G197gat), .A2(G204gat), .ZN(new_n524_));
  NOR2_X1   g323(.A1(G197gat), .A2(G204gat), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n523_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(G197gat), .ZN(new_n527_));
  INV_X1    g326(.A(G204gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G197gat), .A2(G204gat), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(KEYINPUT94), .A3(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n522_), .A2(new_n526_), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT95), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n522_), .A2(new_n526_), .A3(new_n531_), .A4(KEYINPUT95), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT93), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n536_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n537_), .A2(KEYINPUT21), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n519_), .A2(new_n521_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n539_), .B1(new_n537_), .B2(KEYINPUT21), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n534_), .A2(new_n535_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n513_), .B1(new_n516_), .B2(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(G78gat), .B(G106gat), .Z(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n534_), .A2(new_n535_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n538_), .A2(new_n540_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n513_), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n547_), .B(new_n548_), .C1(new_n492_), .C2(new_n493_), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n542_), .A2(new_n544_), .A3(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n544_), .B1(new_n542_), .B2(new_n549_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n510_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  AOI211_X1 g351(.A(new_n541_), .B(new_n513_), .C1(new_n505_), .C2(KEYINPUT29), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n514_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n548_), .B1(new_n554_), .B2(new_n547_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n543_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n542_), .A2(new_n549_), .A3(new_n544_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n556_), .A2(new_n509_), .A3(new_n557_), .A4(new_n500_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n552_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G8gat), .B(G36gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT18), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G64gat), .B(G92gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT32), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G226gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT19), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  AOI22_X1  g368(.A1(new_n423_), .A2(new_n440_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n397_), .A2(KEYINPUT85), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n403_), .A2(KEYINPUT23), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n571_), .A2(new_n572_), .B1(G183gat), .B2(G190gat), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n395_), .B1(new_n573_), .B2(new_n426_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT22), .B(G169gat), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n411_), .B1(new_n575_), .B2(new_n410_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n406_), .A2(new_n398_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n424_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n433_), .A2(new_n435_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n577_), .B1(new_n578_), .B2(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(KEYINPUT20), .B1(new_n547_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT99), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n570_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT20), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n579_), .A2(new_n580_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n578_), .ZN(new_n588_));
  AOI22_X1  g387(.A1(new_n587_), .A2(new_n588_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n586_), .B1(new_n541_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(KEYINPUT99), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n569_), .B1(new_n585_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT97), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n593_), .B1(new_n541_), .B2(new_n589_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n547_), .A2(KEYINPUT97), .A3(new_n582_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n423_), .A2(new_n440_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n586_), .B1(new_n597_), .B2(new_n541_), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n596_), .A2(new_n569_), .A3(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n566_), .B1(new_n592_), .B2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT100), .ZN(new_n601_));
  INV_X1    g400(.A(new_n449_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n602_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n501_), .A2(new_n449_), .A3(new_n504_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G225gat), .A2(G233gat), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n603_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n603_), .A2(KEYINPUT4), .A3(new_n604_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n605_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n608_), .B1(new_n603_), .B2(KEYINPUT4), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n606_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(G1gat), .B(G29gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT98), .B(KEYINPUT0), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G57gat), .B(G85gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n610_), .A2(new_n616_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n606_), .B(new_n615_), .C1(new_n607_), .C2(new_n609_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n441_), .A2(new_n547_), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n590_), .A2(new_n619_), .A3(new_n569_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n596_), .A2(new_n598_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n620_), .B1(new_n621_), .B2(new_n568_), .ZN(new_n622_));
  AOI22_X1  g421(.A1(new_n617_), .A2(new_n618_), .B1(new_n622_), .B2(new_n565_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT100), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n624_), .B(new_n566_), .C1(new_n592_), .C2(new_n599_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n601_), .A2(new_n623_), .A3(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n618_), .A2(KEYINPUT33), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT4), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n505_), .A2(new_n628_), .A3(new_n602_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n603_), .A2(new_n604_), .ZN(new_n630_));
  OAI211_X1 g429(.A(new_n608_), .B(new_n629_), .C1(new_n630_), .C2(new_n628_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT33), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n631_), .A2(new_n632_), .A3(new_n606_), .A4(new_n615_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n627_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n629_), .A2(new_n605_), .ZN(new_n635_));
  OAI221_X1 g434(.A(new_n616_), .B1(new_n630_), .B2(new_n605_), .C1(new_n607_), .C2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n590_), .A2(new_n619_), .A3(new_n569_), .ZN(new_n637_));
  OAI21_X1  g436(.A(KEYINPUT20), .B1(new_n441_), .B2(new_n547_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n638_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n564_), .B(new_n637_), .C1(new_n639_), .C2(new_n569_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n569_), .B1(new_n596_), .B2(new_n598_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n563_), .B1(new_n641_), .B2(new_n620_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n634_), .A2(new_n636_), .A3(new_n640_), .A4(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n559_), .B1(new_n626_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n618_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n615_), .B1(new_n631_), .B2(new_n606_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n559_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n640_), .A2(KEYINPUT27), .ZN(new_n649_));
  INV_X1    g448(.A(new_n591_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n619_), .B1(new_n590_), .B2(KEYINPUT99), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n568_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n596_), .A2(new_n598_), .A3(new_n569_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n564_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n649_), .A2(new_n654_), .ZN(new_n655_));
  XOR2_X1   g454(.A(KEYINPUT101), .B(KEYINPUT27), .Z(new_n656_));
  AOI21_X1  g455(.A(new_n656_), .B1(new_n642_), .B2(new_n640_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n648_), .A2(new_n655_), .A3(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n460_), .B1(new_n644_), .B2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n655_), .A2(new_n657_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n559_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n660_), .A2(new_n647_), .A3(new_n661_), .A4(new_n459_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n392_), .B1(new_n659_), .B2(new_n662_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n360_), .A2(new_n361_), .A3(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n665_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n647_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(new_n291_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n202_), .B1(new_n668_), .B2(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n647_), .A2(G1gat), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n666_), .A2(KEYINPUT38), .A3(new_n667_), .A4(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n286_), .A2(new_n391_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n674_), .A2(new_n309_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n354_), .B1(new_n659_), .B2(new_n662_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(G1gat), .B1(new_n677_), .B2(new_n647_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n671_), .A2(new_n673_), .A3(new_n678_), .ZN(G1324gat));
  INV_X1    g478(.A(KEYINPUT40), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n660_), .A2(G8gat), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n666_), .A2(new_n667_), .A3(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT39), .ZN(new_n683_));
  INV_X1    g482(.A(new_n677_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n660_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n683_), .B1(new_n686_), .B2(G8gat), .ZN(new_n687_));
  AOI211_X1 g486(.A(KEYINPUT39), .B(new_n292_), .C1(new_n684_), .C2(new_n685_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n680_), .B1(new_n682_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n681_), .ZN(new_n691_));
  OAI221_X1 g490(.A(KEYINPUT40), .B1(new_n688_), .B2(new_n687_), .C1(new_n668_), .C2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(G1325gat));
  OAI21_X1  g492(.A(G15gat), .B1(new_n677_), .B2(new_n460_), .ZN(new_n694_));
  XOR2_X1   g493(.A(new_n694_), .B(KEYINPUT41), .Z(new_n695_));
  OR2_X1    g494(.A1(new_n460_), .A2(G15gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n668_), .B2(new_n696_), .ZN(G1326gat));
  OAI21_X1  g496(.A(G22gat), .B1(new_n677_), .B2(new_n661_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT42), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n559_), .A2(new_n288_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n699_), .B1(new_n668_), .B2(new_n700_), .ZN(G1327gat));
  INV_X1    g500(.A(new_n354_), .ZN(new_n702_));
  AOI211_X1 g501(.A(new_n310_), .B(new_n702_), .C1(new_n276_), .C2(new_n285_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(new_n663_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT103), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n703_), .A2(new_n663_), .A3(new_n706_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n705_), .A2(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(G29gat), .B1(new_n708_), .B2(new_n669_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n674_), .A2(new_n310_), .ZN(new_n710_));
  AOI221_X4 g509(.A(KEYINPUT43), .B1(new_n358_), .B2(new_n353_), .C1(new_n659_), .C2(new_n662_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n659_), .A2(new_n662_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n358_), .A2(new_n353_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n712_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n710_), .B1(new_n711_), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  OAI211_X1 g517(.A(KEYINPUT44), .B(new_n710_), .C1(new_n711_), .C2(new_n715_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n669_), .A2(G29gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n709_), .B1(new_n720_), .B2(new_n721_), .ZN(G1328gat));
  NAND3_X1  g521(.A1(new_n718_), .A2(new_n685_), .A3(new_n719_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G36gat), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n660_), .A2(G36gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n705_), .A2(new_n707_), .A3(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT104), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT45), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT104), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n705_), .A2(new_n729_), .A3(new_n707_), .A4(new_n725_), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n727_), .A2(new_n728_), .A3(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n728_), .B1(new_n727_), .B2(new_n730_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n724_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  OAI221_X1 g534(.A(new_n724_), .B1(KEYINPUT105), .B2(KEYINPUT46), .C1(new_n731_), .C2(new_n732_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1329gat));
  INV_X1    g536(.A(G43gat), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n460_), .A2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n718_), .A2(new_n719_), .A3(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n708_), .A2(new_n459_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(new_n738_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n718_), .A2(KEYINPUT106), .A3(new_n719_), .A4(new_n739_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n742_), .A2(new_n744_), .A3(new_n745_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g546(.A(G50gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n708_), .A2(new_n748_), .A3(new_n559_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT108), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT107), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n718_), .A2(new_n751_), .A3(new_n559_), .A4(new_n719_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n752_), .A2(G50gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n718_), .A2(new_n559_), .A3(new_n719_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT107), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n750_), .B1(new_n753_), .B2(new_n755_), .ZN(new_n756_));
  AND4_X1   g555(.A1(new_n750_), .A2(new_n755_), .A3(G50gat), .A4(new_n752_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n749_), .B1(new_n756_), .B2(new_n757_), .ZN(G1331gat));
  INV_X1    g557(.A(G57gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n669_), .B2(KEYINPUT110), .ZN(new_n760_));
  INV_X1    g559(.A(new_n286_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n676_), .A2(new_n761_), .A3(new_n310_), .A4(new_n392_), .ZN(new_n762_));
  AOI211_X1 g561(.A(new_n760_), .B(new_n762_), .C1(KEYINPUT110), .C2(new_n759_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n714_), .A2(new_n309_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n761_), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n765_), .A2(KEYINPUT109), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(KEYINPUT109), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n391_), .B1(new_n659_), .B2(new_n662_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n766_), .A2(new_n767_), .A3(new_n768_), .ZN(new_n769_));
  OR2_X1    g568(.A1(new_n769_), .A2(new_n647_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n763_), .B1(new_n770_), .B2(new_n759_), .ZN(G1332gat));
  OAI21_X1  g570(.A(G64gat), .B1(new_n762_), .B2(new_n660_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT48), .ZN(new_n773_));
  OR2_X1    g572(.A1(new_n660_), .A2(G64gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n769_), .B2(new_n774_), .ZN(G1333gat));
  OAI21_X1  g574(.A(G71gat), .B1(new_n762_), .B2(new_n460_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT49), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n459_), .A2(new_n443_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n769_), .B2(new_n778_), .ZN(G1334gat));
  OAI21_X1  g578(.A(G78gat), .B1(new_n762_), .B2(new_n661_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT50), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n661_), .A2(G78gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n781_), .B1(new_n769_), .B2(new_n782_), .ZN(G1335gat));
  NOR3_X1   g582(.A1(new_n286_), .A2(new_n310_), .A3(new_n702_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n768_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n785_), .A2(G85gat), .A3(new_n647_), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n711_), .A2(new_n715_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n286_), .A2(new_n310_), .A3(new_n391_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n669_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n786_), .B1(new_n790_), .B2(G85gat), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT111), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n791_), .B(new_n792_), .ZN(G1336gat));
  NOR2_X1   g592(.A1(new_n785_), .A2(new_n660_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n794_), .A2(G92gat), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n685_), .A2(G92gat), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT112), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n795_), .B1(new_n789_), .B2(new_n797_), .ZN(G1337gat));
  INV_X1    g597(.A(KEYINPUT113), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT51), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n459_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n800_), .B1(new_n785_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n789_), .A2(new_n459_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n803_), .B2(G99gat), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n799_), .A2(KEYINPUT51), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n804_), .B(new_n805_), .ZN(G1338gat));
  OAI211_X1 g605(.A(new_n559_), .B(new_n788_), .C1(new_n711_), .C2(new_n715_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(G106gat), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT52), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n784_), .A2(new_n768_), .A3(new_n213_), .A4(new_n559_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n809_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n811_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n813_), .A2(new_n814_), .ZN(G1339gat));
  NOR4_X1   g614(.A1(new_n685_), .A2(new_n647_), .A3(new_n559_), .A4(new_n460_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT58), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n818_), .B1(new_n261_), .B2(KEYINPUT116), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n819_), .B1(new_n818_), .B2(new_n261_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n256_), .B(new_n820_), .C1(new_n258_), .C2(new_n259_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n244_), .A2(KEYINPUT12), .A3(new_n252_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT67), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  AOI22_X1  g623(.A1(new_n824_), .A2(new_n257_), .B1(new_n255_), .B2(new_n253_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n819_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n821_), .B(new_n278_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT56), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n828_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT121), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT121), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n827_), .A2(new_n832_), .A3(new_n828_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n829_), .B1(new_n831_), .B2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n371_), .A2(new_n372_), .A3(new_n377_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n375_), .A2(KEYINPUT119), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n378_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n375_), .A2(KEYINPUT119), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n383_), .B(new_n835_), .C1(new_n837_), .C2(new_n838_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n839_), .A2(new_n385_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n269_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n817_), .B1(new_n834_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n829_), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n827_), .A2(new_n832_), .A3(new_n828_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n832_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n843_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n846_), .A2(KEYINPUT58), .A3(new_n269_), .A4(new_n840_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n842_), .A2(new_n714_), .A3(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n840_), .B1(new_n271_), .B2(new_n270_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT120), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT120), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n840_), .B(new_n851_), .C1(new_n271_), .C2(new_n270_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT56), .B1(new_n827_), .B2(KEYINPUT117), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n256_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n819_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT117), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n856_), .A2(new_n857_), .A3(new_n278_), .A4(new_n821_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n854_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(KEYINPUT118), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n827_), .A2(KEYINPUT117), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n861_), .A2(new_n862_), .A3(new_n828_), .A4(new_n858_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n860_), .A2(new_n843_), .A3(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n270_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n853_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n702_), .A2(KEYINPUT57), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n848_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n863_), .A2(new_n843_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n862_), .B1(new_n854_), .B2(new_n858_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n865_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n850_), .A2(new_n852_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(KEYINPUT57), .B1(new_n873_), .B2(new_n702_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n309_), .B1(new_n868_), .B2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(KEYINPUT115), .B1(new_n359_), .B2(new_n391_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT115), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n764_), .A2(new_n877_), .A3(new_n286_), .A4(new_n392_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n876_), .A2(new_n878_), .A3(KEYINPUT54), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n875_), .A2(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(KEYINPUT54), .B1(new_n876_), .B2(new_n878_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n816_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(G113gat), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n883_), .A2(new_n884_), .A3(new_n391_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n882_), .A2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n876_), .A2(new_n878_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n890_), .A2(new_n875_), .A3(new_n879_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n891_), .A2(KEYINPUT59), .A3(new_n816_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n392_), .B1(new_n887_), .B2(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n885_), .B1(new_n893_), .B2(new_n884_), .ZN(G1340gat));
  INV_X1    g693(.A(G120gat), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n895_), .B1(new_n286_), .B2(KEYINPUT60), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n883_), .B(new_n896_), .C1(KEYINPUT60), .C2(new_n895_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n286_), .B1(new_n887_), .B2(new_n892_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n898_), .B2(new_n895_), .ZN(G1341gat));
  AOI21_X1  g698(.A(G127gat), .B1(new_n883_), .B2(new_n310_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n887_), .A2(new_n892_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n310_), .A2(G127gat), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(KEYINPUT122), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n900_), .B1(new_n901_), .B2(new_n903_), .ZN(G1342gat));
  INV_X1    g703(.A(G134gat), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n883_), .A2(new_n905_), .A3(new_n354_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n714_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n907_), .B1(new_n887_), .B2(new_n892_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n906_), .B1(new_n908_), .B2(new_n905_), .ZN(G1343gat));
  NOR2_X1   g708(.A1(new_n880_), .A2(new_n881_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n460_), .A2(new_n669_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n685_), .A2(new_n911_), .A3(new_n661_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n910_), .A2(new_n392_), .A3(new_n913_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(new_n463_), .ZN(G1344gat));
  NOR3_X1   g714(.A1(new_n910_), .A2(new_n286_), .A3(new_n913_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(new_n464_), .ZN(G1345gat));
  OAI211_X1 g716(.A(new_n310_), .B(new_n912_), .C1(new_n880_), .C2(new_n881_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  NAND4_X1  g719(.A1(new_n891_), .A2(KEYINPUT123), .A3(new_n310_), .A4(new_n912_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(KEYINPUT61), .B(G155gat), .ZN(new_n922_));
  AND3_X1   g721(.A1(new_n920_), .A2(new_n921_), .A3(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n922_), .B1(new_n920_), .B2(new_n921_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1346gat));
  INV_X1    g724(.A(G162gat), .ZN(new_n926_));
  NAND4_X1  g725(.A1(new_n891_), .A2(new_n926_), .A3(new_n354_), .A4(new_n912_), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n910_), .A2(new_n907_), .A3(new_n913_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n927_), .B1(new_n928_), .B2(new_n926_), .ZN(G1347gat));
  NOR3_X1   g728(.A1(new_n660_), .A2(new_n460_), .A3(new_n669_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(new_n391_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n931_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n891_), .A2(new_n661_), .A3(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(G169gat), .ZN(new_n934_));
  XOR2_X1   g733(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n910_), .A2(new_n559_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n937_), .A2(new_n575_), .A3(new_n932_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n935_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n933_), .A2(G169gat), .A3(new_n939_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n936_), .A2(new_n938_), .A3(new_n940_), .ZN(G1348gat));
  NAND4_X1  g740(.A1(new_n891_), .A2(new_n761_), .A3(new_n661_), .A4(new_n930_), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n942_), .A2(new_n943_), .A3(G176gat), .ZN(new_n944_));
  XOR2_X1   g743(.A(KEYINPUT125), .B(G176gat), .Z(new_n945_));
  OAI21_X1  g744(.A(new_n944_), .B1(new_n942_), .B2(new_n945_), .ZN(G1349gat));
  NAND2_X1  g745(.A1(new_n930_), .A2(new_n310_), .ZN(new_n947_));
  NOR3_X1   g746(.A1(new_n910_), .A2(new_n559_), .A3(new_n947_), .ZN(new_n948_));
  INV_X1    g747(.A(new_n433_), .ZN(new_n949_));
  INV_X1    g748(.A(new_n947_), .ZN(new_n950_));
  NAND4_X1  g749(.A1(new_n891_), .A2(new_n949_), .A3(new_n661_), .A4(new_n950_), .ZN(new_n951_));
  OAI22_X1  g750(.A1(new_n948_), .A2(G183gat), .B1(new_n951_), .B2(KEYINPUT126), .ZN(new_n952_));
  AND2_X1   g751(.A1(new_n951_), .A2(KEYINPUT126), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n952_), .A2(new_n953_), .ZN(G1350gat));
  NAND4_X1  g753(.A1(new_n937_), .A2(new_n354_), .A3(new_n435_), .A4(new_n930_), .ZN(new_n955_));
  AND3_X1   g754(.A1(new_n937_), .A2(new_n714_), .A3(new_n930_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n955_), .B1(new_n956_), .B2(new_n394_), .ZN(G1351gat));
  NAND3_X1  g756(.A1(new_n460_), .A2(new_n647_), .A3(new_n559_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n958_), .A2(new_n660_), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n891_), .A2(new_n391_), .A3(new_n959_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n960_), .A2(new_n527_), .ZN(new_n961_));
  NAND4_X1  g760(.A1(new_n891_), .A2(G197gat), .A3(new_n391_), .A4(new_n959_), .ZN(new_n962_));
  INV_X1    g761(.A(KEYINPUT127), .ZN(new_n963_));
  OAI21_X1  g762(.A(new_n961_), .B1(new_n962_), .B2(new_n963_), .ZN(new_n964_));
  AND2_X1   g763(.A1(new_n962_), .A2(new_n963_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n964_), .A2(new_n965_), .ZN(G1352gat));
  INV_X1    g765(.A(new_n959_), .ZN(new_n967_));
  NOR3_X1   g766(.A1(new_n910_), .A2(new_n286_), .A3(new_n967_), .ZN(new_n968_));
  XNOR2_X1  g767(.A(new_n968_), .B(new_n528_), .ZN(G1353gat));
  NOR2_X1   g768(.A1(new_n910_), .A2(new_n967_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n970_), .A2(new_n310_), .ZN(new_n971_));
  OAI21_X1  g770(.A(new_n971_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n972_));
  XNOR2_X1  g771(.A(KEYINPUT63), .B(G211gat), .ZN(new_n973_));
  NAND3_X1  g772(.A1(new_n970_), .A2(new_n310_), .A3(new_n973_), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n972_), .A2(new_n974_), .ZN(G1354gat));
  NAND3_X1  g774(.A1(new_n970_), .A2(new_n518_), .A3(new_n354_), .ZN(new_n976_));
  NOR3_X1   g775(.A1(new_n910_), .A2(new_n907_), .A3(new_n967_), .ZN(new_n977_));
  OAI21_X1  g776(.A(new_n976_), .B1(new_n518_), .B2(new_n977_), .ZN(G1355gat));
endmodule


