//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 0 0 0 0 0 1 1 0 0 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 1 1 1 1 0 1 1 1 0 1 0 1 0 1 0 1 0 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n793_, new_n794_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n806_, new_n807_, new_n808_, new_n809_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n957_,
    new_n958_, new_n959_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_,
    new_n973_, new_n975_, new_n976_, new_n978_, new_n979_, new_n980_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n993_, new_n994_,
    new_n995_, new_n996_, new_n997_, new_n998_, new_n1000_, new_n1001_,
    new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1011_, new_n1012_, new_n1014_, new_n1015_,
    new_n1016_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1028_, new_n1029_;
  NOR2_X1   g000(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G169gat), .ZN(new_n203_));
  INV_X1    g002(.A(G190gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT81), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT81), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G190gat), .ZN(new_n207_));
  INV_X1    g006(.A(G183gat), .ZN(new_n208_));
  AND3_X1   g007(.A1(new_n205_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n203_), .B1(new_n209_), .B2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n208_), .A2(KEYINPUT25), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT25), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(G183gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n206_), .A2(G190gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n204_), .A2(KEYINPUT81), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT26), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n219_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  OR3_X1    g028(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n229_), .A2(new_n212_), .A3(new_n213_), .A4(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n215_), .B1(new_n225_), .B2(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n232_), .A2(KEYINPUT82), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT82), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n230_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n226_), .B1(G169gat), .B2(G176gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n216_), .A2(new_n218_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT26), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n239_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n238_), .B1(new_n240_), .B2(new_n223_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n237_), .A2(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n234_), .B1(new_n242_), .B2(new_n215_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G71gat), .B(G99gat), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(G227gat), .ZN(new_n246_));
  INV_X1    g045(.A(G233gat), .ZN(new_n247_));
  OAI21_X1  g046(.A(G15gat), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(G43gat), .ZN(new_n249_));
  INV_X1    g048(.A(G15gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n250_), .A2(G227gat), .A3(G233gat), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n248_), .A2(new_n249_), .A3(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n249_), .B1(new_n248_), .B2(new_n251_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n245_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT30), .ZN(new_n255_));
  INV_X1    g054(.A(new_n251_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n250_), .B1(G227gat), .B2(G233gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(G43gat), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n248_), .A2(new_n249_), .A3(new_n251_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(new_n244_), .A3(new_n259_), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n254_), .A2(new_n255_), .A3(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n255_), .B1(new_n254_), .B2(new_n260_), .ZN(new_n262_));
  OAI22_X1  g061(.A1(new_n233_), .A2(new_n243_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n254_), .A2(new_n260_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT30), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n232_), .A2(KEYINPUT82), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n242_), .A2(new_n234_), .A3(new_n215_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n254_), .A2(new_n255_), .A3(new_n260_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .A4(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n263_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G113gat), .B(G120gat), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(G134gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(G127gat), .ZN(new_n274_));
  INV_X1    g073(.A(G127gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(G134gat), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n274_), .A2(new_n276_), .A3(KEYINPUT83), .ZN(new_n277_));
  AOI21_X1  g076(.A(KEYINPUT83), .B1(new_n274_), .B2(new_n276_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n272_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT83), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n275_), .A2(G134gat), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n273_), .A2(G127gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n280_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n274_), .A2(new_n276_), .A3(KEYINPUT83), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n283_), .A2(new_n284_), .A3(new_n271_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n279_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT84), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n279_), .A2(new_n285_), .A3(KEYINPUT84), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT31), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n288_), .A2(KEYINPUT31), .A3(new_n289_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n270_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT85), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n270_), .A2(KEYINPUT85), .A3(new_n294_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT87), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n292_), .A2(new_n293_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n301_), .A2(KEYINPUT86), .A3(new_n269_), .A4(new_n263_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT86), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n303_), .B1(new_n270_), .B2(new_n294_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n299_), .A2(new_n300_), .A3(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n300_), .B1(new_n299_), .B2(new_n305_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G225gat), .A2(G233gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  OR2_X1    g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G155gat), .A2(G162gat), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n315_), .A2(KEYINPUT90), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G141gat), .A2(G148gat), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT2), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n317_), .A2(KEYINPUT90), .A3(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  OR3_X1    g119(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n322_));
  NAND3_X1  g121(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n314_), .B1(new_n320_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n313_), .A2(KEYINPUT1), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT1), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n327_), .A2(G155gat), .A3(G162gat), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(new_n328_), .A3(new_n312_), .ZN(new_n329_));
  XOR2_X1   g128(.A(G141gat), .B(G148gat), .Z(new_n330_));
  AOI21_X1  g129(.A(KEYINPUT89), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n329_), .A2(new_n330_), .A3(KEYINPUT89), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n325_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n279_), .A2(new_n285_), .A3(KEYINPUT84), .ZN(new_n335_));
  AOI21_X1  g134(.A(KEYINPUT84), .B1(new_n279_), .B2(new_n285_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n334_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT4), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n329_), .A2(new_n330_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT89), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n322_), .A2(new_n323_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n343_), .B(new_n321_), .C1(new_n316_), .C2(new_n319_), .ZN(new_n344_));
  AOI22_X1  g143(.A1(new_n342_), .A2(new_n332_), .B1(new_n344_), .B2(new_n314_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n345_), .A2(new_n285_), .A3(new_n279_), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n337_), .A2(new_n346_), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n311_), .B(new_n339_), .C1(new_n347_), .C2(new_n338_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n337_), .A2(new_n346_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(new_n310_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G1gat), .B(G29gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G57gat), .B(G85gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n351_), .B(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G22gat), .B(G50gat), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT29), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n325_), .B(new_n361_), .C1(new_n331_), .C2(new_n333_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT28), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT28), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n345_), .A2(new_n364_), .A3(new_n361_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G228gat), .A2(G233gat), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT95), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n363_), .A2(new_n365_), .A3(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n368_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n360_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n363_), .A2(new_n365_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n368_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n363_), .A2(new_n365_), .A3(new_n368_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(new_n359_), .A3(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n345_), .A2(new_n361_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(G78gat), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT21), .ZN(new_n380_));
  AND2_X1   g179(.A1(G197gat), .A2(G204gat), .ZN(new_n381_));
  NOR2_X1   g180(.A1(G197gat), .A2(G204gat), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT94), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n380_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT93), .ZN(new_n386_));
  INV_X1    g185(.A(G218gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(G211gat), .ZN(new_n388_));
  INV_X1    g187(.A(G211gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(G218gat), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n386_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n388_), .A2(new_n390_), .A3(new_n386_), .ZN(new_n393_));
  OR2_X1    g192(.A1(G197gat), .A2(G204gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G197gat), .A2(G204gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT94), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n385_), .A2(new_n392_), .A3(new_n393_), .A4(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n394_), .A2(KEYINPUT21), .A3(new_n395_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT91), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  XOR2_X1   g200(.A(KEYINPUT92), .B(KEYINPUT21), .Z(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n396_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n393_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n403_), .B1(new_n404_), .B2(new_n391_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n398_), .B1(new_n401_), .B2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(KEYINPUT95), .A2(G228gat), .A3(G233gat), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n378_), .A2(new_n379_), .A3(new_n406_), .A4(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n406_), .B1(new_n367_), .B2(new_n366_), .ZN(new_n409_));
  OAI21_X1  g208(.A(G78gat), .B1(new_n409_), .B2(new_n377_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n371_), .A2(new_n376_), .A3(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n411_), .B1(new_n371_), .B2(new_n376_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT96), .B(G106gat), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NOR3_X1   g214(.A1(new_n412_), .A2(new_n413_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n411_), .ZN(new_n417_));
  NOR3_X1   g216(.A1(new_n369_), .A2(new_n370_), .A3(new_n360_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n359_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n417_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n371_), .A2(new_n376_), .A3(new_n411_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n414_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n416_), .A2(new_n422_), .ZN(new_n423_));
  XOR2_X1   g222(.A(G8gat), .B(G36gat), .Z(new_n424_));
  XNOR2_X1  g223(.A(G64gat), .B(G92gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  AOI22_X1  g227(.A1(new_n392_), .A2(new_n393_), .B1(new_n402_), .B2(new_n396_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n399_), .B(KEYINPUT91), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT21), .B1(new_n396_), .B2(KEYINPUT94), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n383_), .A2(new_n384_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n404_), .A2(new_n391_), .ZN(new_n434_));
  AOI22_X1  g233(.A1(new_n429_), .A2(new_n430_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n435_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n212_), .B(new_n213_), .C1(G183gat), .C2(G190gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n203_), .A2(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n219_), .A2(KEYINPUT97), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT97), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n440_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n239_), .A2(new_n204_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n442_), .A2(new_n223_), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n439_), .A2(new_n441_), .A3(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n438_), .B1(new_n444_), .B2(new_n231_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT20), .B1(new_n406_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G226gat), .A2(G233gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT19), .ZN(new_n448_));
  NOR3_X1   g247(.A1(new_n436_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n448_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n266_), .A2(new_n435_), .A3(new_n267_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT20), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n452_), .B1(new_n406_), .B2(new_n445_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n450_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n428_), .B1(new_n449_), .B2(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n406_), .B1(new_n233_), .B2(new_n243_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n238_), .A2(new_n440_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n441_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n457_), .B(new_n458_), .C1(new_n223_), .C2(new_n442_), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n459_), .A2(new_n237_), .B1(new_n203_), .B2(new_n437_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n452_), .B1(new_n460_), .B2(new_n435_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n456_), .A2(new_n461_), .A3(new_n450_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n428_), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n451_), .A2(new_n453_), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n462_), .B(new_n463_), .C1(new_n464_), .C2(new_n450_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n455_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT27), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n450_), .B1(new_n456_), .B2(new_n461_), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n451_), .A2(new_n453_), .A3(new_n450_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n428_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(new_n465_), .A3(KEYINPUT27), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n468_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n309_), .A2(new_n358_), .A3(new_n423_), .A4(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n473_), .B1(new_n416_), .B2(new_n422_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n357_), .B1(new_n416_), .B2(new_n422_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT88), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n478_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n299_), .A2(new_n305_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT87), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n299_), .A2(new_n300_), .A3(new_n305_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n481_), .A2(KEYINPUT88), .A3(new_n482_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n476_), .A2(new_n477_), .A3(new_n479_), .A4(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n416_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n338_), .B1(new_n337_), .B2(new_n346_), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT4), .B1(new_n290_), .B2(new_n334_), .ZN(new_n487_));
  NOR3_X1   g286(.A1(new_n486_), .A2(new_n487_), .A3(new_n310_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n350_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n356_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT33), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT100), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n356_), .B1(new_n347_), .B2(new_n311_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n310_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n495_), .A2(new_n455_), .A3(new_n465_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT100), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n351_), .A2(new_n497_), .A3(KEYINPUT33), .A4(new_n356_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n490_), .A2(new_n491_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n492_), .A2(new_n496_), .A3(new_n498_), .A4(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n422_), .ZN(new_n501_));
  OAI211_X1 g300(.A(KEYINPUT32), .B(new_n463_), .C1(new_n469_), .C2(new_n470_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n463_), .A2(KEYINPUT32), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n462_), .B(new_n503_), .C1(new_n464_), .C2(new_n450_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n351_), .A2(new_n356_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n490_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n502_), .B(new_n504_), .C1(new_n505_), .C2(new_n506_), .ZN(new_n507_));
  AND4_X1   g306(.A1(new_n485_), .A2(new_n500_), .A3(new_n501_), .A4(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n475_), .B1(new_n484_), .B2(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(G1gat), .B(G8gat), .Z(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(G22gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n250_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G15gat), .A2(G22gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G1gat), .A2(G8gat), .ZN(new_n515_));
  AOI22_X1  g314(.A1(new_n513_), .A2(new_n514_), .B1(KEYINPUT14), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT76), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  AND2_X1   g317(.A1(G15gat), .A2(G22gat), .ZN(new_n519_));
  NOR2_X1   g318(.A1(G15gat), .A2(G22gat), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n515_), .A2(KEYINPUT14), .ZN(new_n522_));
  NOR3_X1   g321(.A1(new_n521_), .A2(new_n522_), .A3(KEYINPUT76), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n511_), .B1(new_n518_), .B2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G29gat), .B(G36gat), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G43gat), .B(G50gat), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n525_), .A2(new_n527_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n516_), .A2(new_n517_), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT76), .B1(new_n521_), .B2(new_n522_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(new_n533_), .A3(new_n510_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n524_), .A2(new_n531_), .A3(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G229gat), .A2(G233gat), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n529_), .A2(KEYINPUT15), .A3(new_n530_), .ZN(new_n537_));
  AOI21_X1  g336(.A(KEYINPUT15), .B1(new_n529_), .B2(new_n530_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n532_), .A2(new_n533_), .A3(new_n510_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n510_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n535_), .B(new_n536_), .C1(new_n540_), .C2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n531_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n545_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n535_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n536_), .ZN(new_n548_));
  AOI21_X1  g347(.A(KEYINPUT78), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT78), .ZN(new_n550_));
  AOI211_X1 g349(.A(new_n550_), .B(new_n536_), .C1(new_n546_), .C2(new_n535_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n544_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(G113gat), .B(G141gat), .Z(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT79), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G169gat), .B(G197gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n552_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n556_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n544_), .B(new_n558_), .C1(new_n549_), .C2(new_n551_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT80), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n509_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G120gat), .B(G148gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT5), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G176gat), .B(G204gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G57gat), .B(G64gat), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT11), .ZN(new_n569_));
  XOR2_X1   g368(.A(G71gat), .B(G78gat), .Z(new_n570_));
  OR2_X1    g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n568_), .A2(KEYINPUT11), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n570_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n571_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(G106gat), .ZN(new_n575_));
  OR2_X1    g374(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n576_));
  NAND2_X1  g375(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n576_), .A2(KEYINPUT64), .A3(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(KEYINPUT64), .B1(new_n576_), .B2(new_n577_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n575_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT9), .ZN(new_n581_));
  INV_X1    g380(.A(G85gat), .ZN(new_n582_));
  INV_X1    g381(.A(G92gat), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G85gat), .A2(G92gat), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n581_), .B(new_n584_), .C1(new_n586_), .C2(KEYINPUT65), .ZN(new_n587_));
  INV_X1    g386(.A(new_n586_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT65), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(new_n589_), .A3(KEYINPUT9), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G99gat), .A2(G106gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT6), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n580_), .A2(new_n587_), .A3(new_n590_), .A4(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT8), .ZN(new_n594_));
  INV_X1    g393(.A(new_n591_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT67), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n596_), .A2(KEYINPUT6), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT6), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n598_), .A2(KEYINPUT67), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n595_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT66), .ZN(new_n601_));
  INV_X1    g400(.A(G99gat), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(new_n602_), .A3(new_n575_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT7), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT7), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n601_), .A2(new_n605_), .A3(new_n602_), .A4(new_n575_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n598_), .A2(KEYINPUT67), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n596_), .A2(KEYINPUT6), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n607_), .A2(new_n608_), .A3(new_n591_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n600_), .A2(new_n604_), .A3(new_n606_), .A4(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n594_), .B1(new_n610_), .B2(new_n588_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n588_), .A2(new_n594_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n604_), .A2(new_n606_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n612_), .B1(new_n613_), .B2(new_n592_), .ZN(new_n614_));
  OAI211_X1 g413(.A(new_n574_), .B(new_n593_), .C1(new_n611_), .C2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G230gat), .A2(G233gat), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n593_), .B1(new_n611_), .B2(new_n614_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT12), .ZN(new_n619_));
  INV_X1    g418(.A(new_n574_), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n618_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n619_), .B1(new_n618_), .B2(new_n620_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n617_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n618_), .A2(new_n620_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n616_), .B1(new_n624_), .B2(new_n615_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n623_), .A2(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n567_), .B1(new_n627_), .B2(KEYINPUT68), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n628_), .B1(KEYINPUT68), .B2(new_n627_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n624_), .A2(KEYINPUT12), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n618_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n625_), .B1(new_n632_), .B2(new_n617_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n633_), .A2(KEYINPUT69), .A3(new_n567_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n623_), .A2(new_n626_), .A3(new_n567_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT69), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n634_), .A2(new_n637_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n629_), .A2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n641_), .B1(new_n639_), .B2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(KEYINPUT75), .B(KEYINPUT37), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(G232gat), .A2(G233gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT34), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n647_), .A2(KEYINPUT35), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n648_), .B1(new_n618_), .B2(new_n539_), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n607_), .A2(new_n608_), .A3(new_n591_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n591_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n586_), .B1(new_n652_), .B2(new_n613_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n592_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n604_), .A2(new_n606_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  OAI22_X1  g455(.A1(new_n653_), .A2(new_n594_), .B1(new_n656_), .B2(new_n612_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT71), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n657_), .A2(new_n658_), .A3(new_n531_), .A4(new_n593_), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n593_), .B(new_n531_), .C1(new_n611_), .C2(new_n614_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT71), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT74), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n649_), .A2(new_n659_), .A3(new_n661_), .A4(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT72), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n647_), .A2(KEYINPUT35), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT72), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n649_), .A2(new_n659_), .A3(new_n661_), .A4(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n664_), .A2(new_n666_), .A3(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n663_), .A2(KEYINPUT72), .A3(new_n665_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(G190gat), .B(G218gat), .ZN(new_n671_));
  XNOR2_X1  g470(.A(G134gat), .B(G162gat), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT36), .Z(new_n674_));
  AND3_X1   g473(.A1(new_n669_), .A2(new_n670_), .A3(new_n674_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(KEYINPUT73), .B(KEYINPUT36), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n673_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n679_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n645_), .B1(new_n675_), .B2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n669_), .A2(new_n670_), .A3(new_n674_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n663_), .A2(KEYINPUT72), .A3(new_n665_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n668_), .A2(new_n666_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n664_), .B2(new_n684_), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n682_), .B(new_n644_), .C1(new_n685_), .C2(new_n679_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n681_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(G231gat), .A2(G233gat), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n574_), .B(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(new_n543_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT77), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(G127gat), .B(G155gat), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT16), .ZN(new_n694_));
  XNOR2_X1  g493(.A(G183gat), .B(G211gat), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n694_), .B(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(KEYINPUT17), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n692_), .B(new_n697_), .ZN(new_n698_));
  OR3_X1    g497(.A1(new_n690_), .A2(KEYINPUT17), .A3(new_n696_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n687_), .A2(new_n701_), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n563_), .A2(new_n643_), .A3(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(G1gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n703_), .A2(new_n704_), .A3(new_n357_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n706_), .A2(KEYINPUT38), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n706_), .A2(KEYINPUT38), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n705_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT101), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n682_), .B1(new_n685_), .B2(new_n679_), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n509_), .A2(new_n710_), .A3(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n710_), .B1(new_n509_), .B2(new_n711_), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n643_), .A2(new_n700_), .A3(new_n560_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT102), .B1(new_n714_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n714_), .A2(KEYINPUT102), .A3(new_n716_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n358_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  OAI221_X1 g519(.A(new_n709_), .B1(new_n707_), .B2(new_n705_), .C1(new_n720_), .C2(new_n704_), .ZN(G1324gat));
  INV_X1    g520(.A(G8gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n703_), .A2(new_n722_), .A3(new_n473_), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n473_), .B(new_n716_), .C1(new_n712_), .C2(new_n713_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n724_), .A2(new_n725_), .A3(G8gat), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n725_), .B1(new_n724_), .B2(G8gat), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n727_), .A2(new_n728_), .A3(KEYINPUT39), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT39), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n724_), .A2(G8gat), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT104), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n730_), .B1(new_n732_), .B2(new_n726_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n723_), .B1(new_n729_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT40), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  OAI211_X1 g535(.A(KEYINPUT40), .B(new_n723_), .C1(new_n729_), .C2(new_n733_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(G1325gat));
  NAND2_X1  g537(.A1(new_n479_), .A2(new_n483_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n703_), .A2(new_n250_), .A3(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n719_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n739_), .B1(new_n741_), .B2(new_n717_), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n742_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(KEYINPUT41), .B1(new_n742_), .B2(G15gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(G1326gat));
  INV_X1    g544(.A(new_n423_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n703_), .A2(new_n512_), .A3(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n741_), .B2(new_n717_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT42), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n748_), .A2(new_n749_), .A3(G22gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n748_), .B2(G22gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n747_), .B1(new_n750_), .B2(new_n751_), .ZN(G1327gat));
  INV_X1    g551(.A(new_n643_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n711_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n701_), .A2(new_n754_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n563_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(G29gat), .B1(new_n758_), .B2(new_n357_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n509_), .A2(new_n687_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT43), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n700_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n560_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n753_), .A2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n509_), .A2(KEYINPUT43), .A3(new_n687_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n762_), .A2(new_n764_), .A3(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT44), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n762_), .A2(KEYINPUT44), .A3(new_n764_), .A4(new_n765_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n357_), .A2(G29gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n759_), .B1(new_n770_), .B2(new_n771_), .ZN(G1328gat));
  OR2_X1    g571(.A1(new_n473_), .A2(KEYINPUT105), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n473_), .A2(KEYINPUT105), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n757_), .A2(G36gat), .A3(new_n776_), .ZN(new_n777_));
  XOR2_X1   g576(.A(new_n777_), .B(KEYINPUT45), .Z(new_n778_));
  NAND3_X1  g577(.A1(new_n768_), .A2(new_n473_), .A3(new_n769_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(G36gat), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n778_), .B(new_n780_), .C1(KEYINPUT106), .C2(KEYINPUT46), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(G1329gat));
  NAND3_X1  g584(.A1(new_n770_), .A2(G43gat), .A3(new_n309_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n739_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n249_), .B1(new_n757_), .B2(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n786_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n786_), .B2(new_n788_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n790_), .A2(new_n791_), .ZN(G1330gat));
  AOI21_X1  g591(.A(G50gat), .B1(new_n758_), .B2(new_n746_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n746_), .A2(G50gat), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n770_), .B2(new_n794_), .ZN(G1331gat));
  AND2_X1   g594(.A1(new_n509_), .A2(new_n763_), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n643_), .A2(new_n701_), .A3(new_n687_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n358_), .B1(new_n798_), .B2(KEYINPUT108), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n799_), .B1(KEYINPUT108), .B2(new_n798_), .ZN(new_n800_));
  INV_X1    g599(.A(G57gat), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n643_), .A2(new_n701_), .A3(new_n562_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n714_), .A2(new_n802_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n358_), .A2(new_n801_), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n800_), .A2(new_n801_), .B1(new_n803_), .B2(new_n804_), .ZN(G1332gat));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n775_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(G64gat), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT48), .ZN(new_n808_));
  OR3_X1    g607(.A1(new_n798_), .A2(G64gat), .A3(new_n776_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(G1333gat));
  NAND2_X1  g609(.A1(new_n803_), .A2(new_n739_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(G71gat), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(KEYINPUT49), .ZN(new_n813_));
  OR3_X1    g612(.A1(new_n798_), .A2(G71gat), .A3(new_n787_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(G1334gat));
  AOI21_X1  g614(.A(new_n379_), .B1(new_n803_), .B2(new_n746_), .ZN(new_n816_));
  XOR2_X1   g615(.A(new_n816_), .B(KEYINPUT50), .Z(new_n817_));
  NAND4_X1  g616(.A1(new_n796_), .A2(new_n379_), .A3(new_n746_), .A4(new_n797_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(G1335gat));
  NOR2_X1   g618(.A1(new_n643_), .A2(new_n755_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n796_), .A2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n582_), .B1(new_n821_), .B2(new_n358_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n762_), .A2(new_n765_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n643_), .A2(new_n560_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n357_), .A2(G85gat), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(KEYINPUT109), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n822_), .B1(new_n825_), .B2(new_n827_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(KEYINPUT110), .ZN(G1336gat));
  INV_X1    g628(.A(new_n821_), .ZN(new_n830_));
  AOI21_X1  g629(.A(G92gat), .B1(new_n830_), .B2(new_n473_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n825_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n775_), .A2(G92gat), .ZN(new_n833_));
  XOR2_X1   g632(.A(new_n833_), .B(KEYINPUT111), .Z(new_n834_));
  AOI21_X1  g633(.A(new_n831_), .B1(new_n832_), .B2(new_n834_), .ZN(G1337gat));
  OAI21_X1  g634(.A(G99gat), .B1(new_n825_), .B2(new_n787_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n309_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n821_), .B2(new_n837_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g638(.A1(new_n830_), .A2(new_n575_), .A3(new_n746_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n823_), .A2(new_n746_), .A3(new_n824_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n841_), .A2(new_n842_), .A3(G106gat), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n842_), .B1(new_n841_), .B2(G106gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n840_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n840_), .B(new_n846_), .C1(new_n843_), .C2(new_n844_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(G1339gat));
  NAND3_X1  g649(.A1(new_n643_), .A2(new_n561_), .A3(new_n702_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(KEYINPUT54), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n643_), .A2(new_n702_), .A3(new_n853_), .A4(new_n561_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n535_), .B(new_n548_), .C1(new_n540_), .C2(new_n543_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n547_), .A2(new_n536_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n857_), .A2(new_n556_), .A3(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n559_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT114), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT114), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n559_), .A2(new_n862_), .A3(new_n859_), .ZN(new_n863_));
  AOI22_X1  g662(.A1(new_n861_), .A2(new_n863_), .B1(new_n634_), .B2(new_n637_), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n617_), .B(KEYINPUT55), .C1(new_n621_), .C2(new_n622_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT113), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n632_), .A2(KEYINPUT113), .A3(KEYINPUT55), .A4(new_n617_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT55), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n623_), .A2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n615_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n616_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n867_), .A2(new_n868_), .A3(new_n870_), .A4(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n567_), .ZN(new_n875_));
  AND3_X1   g674(.A1(new_n874_), .A2(KEYINPUT56), .A3(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(KEYINPUT56), .B1(new_n874_), .B2(new_n875_), .ZN(new_n877_));
  OAI211_X1 g676(.A(KEYINPUT58), .B(new_n864_), .C1(new_n876_), .C2(new_n877_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n878_), .A2(new_n687_), .ZN(new_n879_));
  XOR2_X1   g678(.A(KEYINPUT117), .B(KEYINPUT58), .Z(new_n880_));
  AOI21_X1  g679(.A(KEYINPUT69), .B1(new_n633_), .B2(new_n567_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n635_), .A2(new_n636_), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n559_), .A2(new_n862_), .A3(new_n859_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n862_), .B1(new_n559_), .B2(new_n859_), .ZN(new_n884_));
  OAI22_X1  g683(.A1(new_n881_), .A2(new_n882_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n874_), .A2(new_n875_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT56), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n874_), .A2(KEYINPUT56), .A3(new_n875_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n885_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT116), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n880_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n891_), .B(new_n864_), .C1(new_n876_), .C2(new_n877_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n879_), .B1(new_n892_), .B2(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n876_), .A2(new_n877_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n638_), .A2(new_n560_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n883_), .A2(new_n884_), .ZN(new_n898_));
  OAI22_X1  g697(.A1(new_n896_), .A2(new_n897_), .B1(new_n639_), .B2(new_n898_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n899_), .A2(KEYINPUT57), .A3(new_n711_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n897_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n898_), .B1(new_n638_), .B2(new_n629_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n711_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  XOR2_X1   g702(.A(KEYINPUT115), .B(KEYINPUT57), .Z(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n895_), .A2(new_n900_), .A3(new_n905_), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n906_), .A2(KEYINPUT118), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n700_), .B1(new_n906_), .B2(KEYINPUT118), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n856_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n309_), .A2(new_n357_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n423_), .A2(new_n474_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  OAI21_X1  g712(.A(KEYINPUT59), .B1(new_n909_), .B2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT119), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n878_), .A2(new_n687_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n880_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n864_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(new_n918_), .B2(KEYINPUT116), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n916_), .B1(new_n919_), .B2(new_n893_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n904_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n921_), .B1(new_n899_), .B2(new_n711_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n915_), .B1(new_n920_), .B2(new_n922_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n895_), .A2(KEYINPUT119), .A3(new_n905_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n923_), .A2(new_n924_), .A3(new_n900_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n701_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n855_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n913_), .A2(KEYINPUT59), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n914_), .A2(new_n562_), .A3(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(G113gat), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n909_), .A2(new_n913_), .ZN(new_n932_));
  INV_X1    g731(.A(new_n932_), .ZN(new_n933_));
  OR2_X1    g732(.A1(new_n763_), .A2(G113gat), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n931_), .B1(new_n933_), .B2(new_n934_), .ZN(G1340gat));
  INV_X1    g734(.A(G120gat), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n643_), .B1(new_n927_), .B2(new_n928_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n936_), .B1(new_n937_), .B2(new_n914_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n643_), .A2(KEYINPUT60), .ZN(new_n939_));
  MUX2_X1   g738(.A(KEYINPUT60), .B(new_n939_), .S(new_n936_), .Z(new_n940_));
  AND2_X1   g739(.A1(new_n932_), .A2(new_n940_), .ZN(new_n941_));
  OAI21_X1  g740(.A(KEYINPUT120), .B1(new_n938_), .B2(new_n941_), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT59), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n906_), .A2(KEYINPUT118), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(new_n701_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n906_), .A2(KEYINPUT118), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n855_), .B1(new_n945_), .B2(new_n946_), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n943_), .B1(new_n947_), .B2(new_n912_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n856_), .B1(new_n925_), .B2(new_n701_), .ZN(new_n949_));
  INV_X1    g748(.A(new_n928_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n753_), .B1(new_n949_), .B2(new_n950_), .ZN(new_n951_));
  OAI21_X1  g750(.A(G120gat), .B1(new_n948_), .B2(new_n951_), .ZN(new_n952_));
  INV_X1    g751(.A(KEYINPUT120), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n932_), .A2(new_n940_), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n952_), .A2(new_n953_), .A3(new_n954_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n942_), .A2(new_n955_), .ZN(G1341gat));
  NAND3_X1  g755(.A1(new_n914_), .A2(new_n700_), .A3(new_n929_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n957_), .A2(G127gat), .ZN(new_n958_));
  NAND3_X1  g757(.A1(new_n932_), .A2(new_n275_), .A3(new_n700_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n958_), .A2(new_n959_), .ZN(G1342gat));
  AOI21_X1  g759(.A(G134gat), .B1(new_n932_), .B2(new_n754_), .ZN(new_n961_));
  AND2_X1   g760(.A1(new_n914_), .A2(new_n929_), .ZN(new_n962_));
  INV_X1    g761(.A(new_n687_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(KEYINPUT121), .B(G134gat), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n963_), .A2(new_n964_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n961_), .B1(new_n962_), .B2(new_n965_), .ZN(G1343gat));
  NOR3_X1   g765(.A1(new_n775_), .A2(new_n739_), .A3(new_n477_), .ZN(new_n967_));
  XNOR2_X1  g766(.A(new_n967_), .B(KEYINPUT122), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n947_), .A2(new_n968_), .ZN(new_n969_));
  INV_X1    g768(.A(new_n969_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n970_), .A2(new_n560_), .ZN(new_n971_));
  XNOR2_X1  g770(.A(new_n971_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g771(.A1(new_n970_), .A2(new_n753_), .ZN(new_n973_));
  XNOR2_X1  g772(.A(new_n973_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g773(.A1(new_n969_), .A2(new_n701_), .ZN(new_n975_));
  XOR2_X1   g774(.A(KEYINPUT61), .B(G155gat), .Z(new_n976_));
  XNOR2_X1  g775(.A(new_n975_), .B(new_n976_), .ZN(G1346gat));
  AOI21_X1  g776(.A(G162gat), .B1(new_n970_), .B2(new_n754_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n687_), .A2(G162gat), .ZN(new_n979_));
  XOR2_X1   g778(.A(new_n979_), .B(KEYINPUT123), .Z(new_n980_));
  AOI21_X1  g779(.A(new_n978_), .B1(new_n970_), .B2(new_n980_), .ZN(G1347gat));
  NOR2_X1   g780(.A1(new_n776_), .A2(new_n357_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n982_), .A2(new_n739_), .ZN(new_n983_));
  NOR2_X1   g782(.A1(new_n983_), .A2(new_n746_), .ZN(new_n984_));
  NAND3_X1  g783(.A1(new_n927_), .A2(new_n560_), .A3(new_n984_), .ZN(new_n985_));
  INV_X1    g784(.A(KEYINPUT62), .ZN(new_n986_));
  AND4_X1   g785(.A1(KEYINPUT124), .A2(new_n985_), .A3(new_n986_), .A4(G169gat), .ZN(new_n987_));
  OAI21_X1  g786(.A(G169gat), .B1(new_n986_), .B2(KEYINPUT124), .ZN(new_n988_));
  INV_X1    g787(.A(new_n988_), .ZN(new_n989_));
  AOI22_X1  g788(.A1(new_n985_), .A2(new_n989_), .B1(KEYINPUT124), .B2(new_n986_), .ZN(new_n990_));
  XOR2_X1   g789(.A(KEYINPUT22), .B(G169gat), .Z(new_n991_));
  OAI22_X1  g790(.A1(new_n987_), .A2(new_n990_), .B1(new_n985_), .B2(new_n991_), .ZN(G1348gat));
  NAND2_X1  g791(.A1(new_n927_), .A2(new_n984_), .ZN(new_n993_));
  INV_X1    g792(.A(new_n993_), .ZN(new_n994_));
  AOI21_X1  g793(.A(G176gat), .B1(new_n994_), .B2(new_n753_), .ZN(new_n995_));
  NOR2_X1   g794(.A1(new_n909_), .A2(new_n746_), .ZN(new_n996_));
  INV_X1    g795(.A(G176gat), .ZN(new_n997_));
  NOR3_X1   g796(.A1(new_n983_), .A2(new_n997_), .A3(new_n643_), .ZN(new_n998_));
  AOI21_X1  g797(.A(new_n995_), .B1(new_n996_), .B2(new_n998_), .ZN(G1349gat));
  NOR2_X1   g798(.A1(new_n439_), .A2(new_n441_), .ZN(new_n1000_));
  NOR2_X1   g799(.A1(new_n701_), .A2(new_n1000_), .ZN(new_n1001_));
  NAND2_X1  g800(.A1(new_n994_), .A2(new_n1001_), .ZN(new_n1002_));
  INV_X1    g801(.A(KEYINPUT125), .ZN(new_n1003_));
  NOR2_X1   g802(.A1(new_n983_), .A2(new_n701_), .ZN(new_n1004_));
  AND2_X1   g803(.A1(new_n996_), .A2(new_n1004_), .ZN(new_n1005_));
  OAI211_X1 g804(.A(new_n1002_), .B(new_n1003_), .C1(new_n1005_), .C2(G183gat), .ZN(new_n1006_));
  NOR3_X1   g805(.A1(new_n993_), .A2(new_n1000_), .A3(new_n701_), .ZN(new_n1007_));
  AOI21_X1  g806(.A(G183gat), .B1(new_n996_), .B2(new_n1004_), .ZN(new_n1008_));
  OAI21_X1  g807(.A(KEYINPUT125), .B1(new_n1007_), .B2(new_n1008_), .ZN(new_n1009_));
  NAND2_X1  g808(.A1(new_n1006_), .A2(new_n1009_), .ZN(G1350gat));
  OAI21_X1  g809(.A(G190gat), .B1(new_n993_), .B2(new_n963_), .ZN(new_n1011_));
  OR2_X1    g810(.A1(new_n711_), .A2(new_n443_), .ZN(new_n1012_));
  OAI21_X1  g811(.A(new_n1011_), .B1(new_n993_), .B2(new_n1012_), .ZN(G1351gat));
  NAND4_X1  g812(.A1(new_n947_), .A2(new_n746_), .A3(new_n787_), .A4(new_n982_), .ZN(new_n1014_));
  NOR2_X1   g813(.A1(new_n1014_), .A2(new_n763_), .ZN(new_n1015_));
  INV_X1    g814(.A(G197gat), .ZN(new_n1016_));
  XNOR2_X1  g815(.A(new_n1015_), .B(new_n1016_), .ZN(G1352gat));
  NOR2_X1   g816(.A1(new_n1014_), .A2(new_n643_), .ZN(new_n1018_));
  NAND2_X1  g817(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n1019_));
  NAND2_X1  g818(.A1(new_n1018_), .A2(new_n1019_), .ZN(new_n1020_));
  XOR2_X1   g819(.A(KEYINPUT126), .B(G204gat), .Z(new_n1021_));
  OAI21_X1  g820(.A(new_n1020_), .B1(new_n1018_), .B2(new_n1021_), .ZN(G1353gat));
  AOI21_X1  g821(.A(new_n701_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n1023_));
  XNOR2_X1  g822(.A(new_n1023_), .B(KEYINPUT127), .ZN(new_n1024_));
  NOR2_X1   g823(.A1(new_n1014_), .A2(new_n1024_), .ZN(new_n1025_));
  NOR2_X1   g824(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1026_));
  XNOR2_X1  g825(.A(new_n1025_), .B(new_n1026_), .ZN(G1354gat));
  OAI21_X1  g826(.A(G218gat), .B1(new_n1014_), .B2(new_n963_), .ZN(new_n1028_));
  NAND2_X1  g827(.A1(new_n754_), .A2(new_n387_), .ZN(new_n1029_));
  OAI21_X1  g828(.A(new_n1028_), .B1(new_n1014_), .B2(new_n1029_), .ZN(G1355gat));
endmodule


