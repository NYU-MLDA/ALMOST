//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n627_, new_n628_, new_n629_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n902_, new_n903_, new_n905_, new_n906_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT21), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G218gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G211gat), .ZN(new_n206_));
  INV_X1    g005(.A(G211gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G218gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT84), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n206_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n207_), .A2(G218gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n205_), .A2(G211gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT84), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n204_), .A2(new_n210_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n202_), .A2(new_n203_), .ZN(new_n215_));
  AND3_X1   g014(.A1(new_n206_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n209_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n215_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G197gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n219_), .A2(KEYINPUT83), .A3(G204gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT21), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT83), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n221_), .B1(new_n222_), .B2(new_n202_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n214_), .B1(new_n218_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G228gat), .A2(G233gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT81), .ZN(new_n226_));
  XOR2_X1   g025(.A(new_n226_), .B(KEYINPUT82), .Z(new_n227_));
  OR2_X1    g026(.A1(G155gat), .A2(G162gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G155gat), .A2(G162gat), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G141gat), .A2(G148gat), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT78), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT2), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n235_));
  INV_X1    g034(.A(G141gat), .ZN(new_n236_));
  INV_X1    g035(.A(G148gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n234_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n233_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n230_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT1), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n228_), .A2(new_n243_), .A3(new_n229_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n236_), .A2(new_n237_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n244_), .A2(new_n231_), .A3(new_n245_), .A4(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n242_), .A2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT80), .B1(new_n248_), .B2(KEYINPUT29), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT80), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT29), .ZN(new_n251_));
  AOI211_X1 g050(.A(new_n250_), .B(new_n251_), .C1(new_n242_), .C2(new_n247_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n224_), .B(new_n227_), .C1(new_n249_), .C2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n224_), .A2(KEYINPUT86), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n213_), .A2(new_n210_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n219_), .A2(G204gat), .ZN(new_n256_));
  INV_X1    g055(.A(G204gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(G197gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  OAI211_X1 g058(.A(KEYINPUT21), .B(new_n220_), .C1(new_n259_), .C2(KEYINPUT83), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n255_), .A2(new_n260_), .A3(new_n215_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT86), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n261_), .A2(new_n262_), .A3(new_n214_), .ZN(new_n263_));
  XOR2_X1   g062(.A(KEYINPUT85), .B(KEYINPUT29), .Z(new_n264_));
  AOI22_X1  g063(.A1(new_n254_), .A2(new_n263_), .B1(new_n248_), .B2(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n253_), .B1(new_n265_), .B2(new_n226_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G78gat), .B(G106gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n267_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n253_), .B(new_n269_), .C1(new_n265_), .C2(new_n226_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT87), .B1(new_n266_), .B2(new_n267_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n242_), .A2(new_n251_), .A3(new_n247_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT79), .B(KEYINPUT28), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(G22gat), .B(G50gat), .Z(new_n278_));
  NAND2_X1  g077(.A1(new_n273_), .A2(new_n275_), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n277_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n278_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n271_), .B1(new_n272_), .B2(new_n283_), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n268_), .A2(new_n282_), .A3(KEYINPUT87), .A4(new_n270_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT4), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G127gat), .B(G134gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G113gat), .B(G120gat), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n289_), .A2(new_n290_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n248_), .A2(new_n288_), .A3(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G225gat), .A2(G233gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT94), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n242_), .A2(KEYINPUT93), .A3(new_n247_), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n291_), .A2(new_n292_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n293_), .A2(KEYINPUT93), .A3(new_n242_), .A4(new_n247_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n298_), .B1(new_n303_), .B2(KEYINPUT4), .ZN(new_n304_));
  AOI211_X1 g103(.A(KEYINPUT94), .B(new_n288_), .C1(new_n301_), .C2(new_n302_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n297_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(new_n295_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G1gat), .B(G29gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(G85gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT0), .B(G57gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n309_), .B(new_n310_), .Z(new_n311_));
  AND3_X1   g110(.A1(new_n306_), .A2(new_n307_), .A3(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n311_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NOR3_X1   g113(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n315_));
  AND2_X1   g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316_));
  NOR2_X1   g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n315_), .B1(new_n318_), .B2(KEYINPUT24), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT26), .B(G190gat), .ZN(new_n320_));
  INV_X1    g119(.A(G183gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT25), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT25), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(KEYINPUT73), .A3(G183gat), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT73), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n325_), .B1(new_n321_), .B2(KEYINPUT25), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n320_), .A2(new_n322_), .A3(new_n324_), .A4(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n319_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G183gat), .A2(G190gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT75), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n331_), .A2(G183gat), .A3(G190gat), .ZN(new_n332_));
  AOI21_X1  g131(.A(KEYINPUT23), .B1(new_n330_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT74), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT23), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n337_));
  AOI22_X1  g136(.A1(new_n336_), .A2(new_n337_), .B1(G183gat), .B2(G190gat), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n333_), .A2(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(G183gat), .A2(G190gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n330_), .A2(new_n332_), .A3(KEYINPUT23), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n336_), .A2(G183gat), .A3(G190gat), .A4(new_n337_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n340_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(G169gat), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  OAI22_X1  g145(.A1(new_n328_), .A2(new_n339_), .B1(new_n343_), .B2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G71gat), .B(G99gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(G43gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n347_), .B(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G227gat), .A2(G233gat), .ZN(new_n351_));
  INV_X1    g150(.A(G15gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT30), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n350_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n350_), .A2(new_n354_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT76), .B(KEYINPUT31), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n300_), .B(new_n358_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n356_), .A2(KEYINPUT77), .A3(new_n357_), .A4(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT77), .ZN(new_n361_));
  INV_X1    g160(.A(new_n357_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n361_), .B1(new_n362_), .B2(new_n355_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n356_), .A2(KEYINPUT77), .A3(new_n357_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n359_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n363_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n314_), .A2(new_n360_), .A3(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n287_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT24), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT89), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT89), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT24), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(new_n372_), .A3(new_n317_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G169gat), .B(G176gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n373_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(G190gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT26), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT26), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(G190gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n323_), .A2(G183gat), .ZN(new_n381_));
  AND4_X1   g180(.A1(new_n378_), .A2(new_n380_), .A3(new_n322_), .A4(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n376_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n341_), .A2(new_n342_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n340_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n385_), .B1(new_n333_), .B2(new_n338_), .ZN(new_n386_));
  AOI22_X1  g185(.A1(new_n383_), .A2(new_n384_), .B1(new_n386_), .B2(new_n345_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n254_), .A2(new_n263_), .A3(new_n387_), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n347_), .A2(KEYINPUT91), .A3(new_n224_), .ZN(new_n389_));
  AOI21_X1  g188(.A(KEYINPUT91), .B1(new_n347_), .B2(new_n224_), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n388_), .B(KEYINPUT20), .C1(new_n389_), .C2(new_n390_), .ZN(new_n391_));
  AND3_X1   g190(.A1(KEYINPUT19), .A2(G226gat), .A3(G233gat), .ZN(new_n392_));
  AOI21_X1  g191(.A(KEYINPUT19), .B1(G226gat), .B2(G233gat), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n391_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT95), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n391_), .A2(KEYINPUT95), .A3(new_n394_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n384_), .A2(new_n385_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n345_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n319_), .B(new_n327_), .C1(new_n338_), .C2(new_n333_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n400_), .A2(new_n261_), .A3(new_n214_), .A4(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n386_), .A2(new_n345_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n370_), .A2(new_n372_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(new_n318_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n320_), .A2(new_n322_), .A3(new_n381_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n384_), .A2(new_n405_), .A3(new_n406_), .A4(new_n373_), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n403_), .A2(new_n407_), .B1(new_n261_), .B2(new_n214_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT90), .ZN(new_n409_));
  OAI211_X1 g208(.A(KEYINPUT20), .B(new_n402_), .C1(new_n408_), .C2(new_n409_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n408_), .A2(new_n409_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n394_), .B(KEYINPUT88), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n397_), .A2(new_n398_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT96), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G8gat), .B(G36gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G64gat), .B(G92gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n416_), .A2(new_n417_), .A3(new_n423_), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n395_), .A2(new_n396_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n422_), .B1(new_n425_), .B2(new_n398_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n403_), .A2(new_n407_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n409_), .B1(new_n427_), .B2(new_n224_), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT20), .B1(new_n347_), .B2(new_n224_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n408_), .A2(new_n409_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n414_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT20), .B1(new_n392_), .B2(new_n393_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n434_), .B1(new_n427_), .B2(new_n224_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n390_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n347_), .A2(KEYINPUT91), .A3(new_n224_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n435_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n432_), .A2(new_n423_), .A3(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n439_), .A2(KEYINPUT96), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n424_), .B(KEYINPUT27), .C1(new_n426_), .C2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT27), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n413_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n435_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n444_), .B1(new_n390_), .B2(new_n389_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n422_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n442_), .B1(new_n439_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT97), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT97), .ZN(new_n449_));
  OAI211_X1 g248(.A(new_n449_), .B(new_n442_), .C1(new_n439_), .C2(new_n446_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n368_), .A2(new_n441_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n313_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n306_), .A2(new_n307_), .A3(new_n311_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n284_), .A2(new_n453_), .A3(new_n454_), .A4(new_n285_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n455_), .B1(new_n448_), .B2(new_n450_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT33), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n454_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n443_), .A2(new_n422_), .A3(new_n445_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n443_), .A2(new_n445_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n423_), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n295_), .B(new_n294_), .C1(new_n304_), .C2(new_n305_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n311_), .B1(new_n303_), .B2(new_n296_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n458_), .A2(new_n459_), .A3(new_n461_), .A4(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n454_), .A2(new_n457_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n422_), .A2(KEYINPUT32), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  OAI22_X1  g267(.A1(new_n312_), .A2(new_n313_), .B1(new_n468_), .B2(new_n460_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n467_), .B1(new_n425_), .B2(new_n398_), .ZN(new_n470_));
  OAI22_X1  g269(.A1(new_n465_), .A2(new_n466_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n456_), .A2(new_n441_), .B1(new_n471_), .B2(new_n286_), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n366_), .A2(new_n360_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n452_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT69), .B(G8gat), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(G1gat), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT14), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G15gat), .B(G22gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G1gat), .B(G8gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  XOR2_X1   g282(.A(G29gat), .B(G36gat), .Z(new_n484_));
  XOR2_X1   g283(.A(G43gat), .B(G50gat), .Z(new_n485_));
  XOR2_X1   g284(.A(new_n484_), .B(new_n485_), .Z(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n483_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT72), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n482_), .A2(new_n486_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n491_), .A2(G229gat), .A3(G233gat), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n486_), .B(KEYINPUT15), .Z(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n482_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G229gat), .A2(G233gat), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n494_), .A2(new_n495_), .A3(new_n488_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n492_), .A2(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(G113gat), .B(G141gat), .Z(new_n498_));
  XNOR2_X1  g297(.A(G169gat), .B(G197gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n497_), .B(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n474_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT37), .ZN(new_n504_));
  XOR2_X1   g303(.A(G85gat), .B(G92gat), .Z(new_n505_));
  NOR2_X1   g304(.A1(G99gat), .A2(G106gat), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT7), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G99gat), .A2(G106gat), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT6), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n505_), .B1(new_n508_), .B2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT8), .ZN(new_n513_));
  XOR2_X1   g312(.A(KEYINPUT10), .B(G99gat), .Z(new_n514_));
  INV_X1    g313(.A(G106gat), .ZN(new_n515_));
  AOI22_X1  g314(.A1(KEYINPUT9), .A2(new_n505_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(G85gat), .ZN(new_n517_));
  INV_X1    g316(.A(G92gat), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n517_), .A2(new_n518_), .A3(KEYINPUT9), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n511_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n516_), .A2(new_n520_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n513_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT64), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n513_), .A2(new_n521_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT64), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n523_), .A2(new_n526_), .A3(new_n493_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT35), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G232gat), .A2(G233gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT34), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  AOI22_X1  g330(.A1(new_n522_), .A2(new_n487_), .B1(new_n528_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n527_), .A2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n531_), .A2(new_n528_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G190gat), .B(G218gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G134gat), .B(G162gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n538_), .A2(KEYINPUT36), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n527_), .B(new_n532_), .C1(new_n528_), .C2(new_n531_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n535_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n538_), .B(KEYINPUT36), .Z(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n544_), .B1(new_n535_), .B2(new_n540_), .ZN(new_n545_));
  OAI211_X1 g344(.A(KEYINPUT68), .B(new_n504_), .C1(new_n542_), .C2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n535_), .A2(new_n540_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n543_), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n504_), .A2(KEYINPUT68), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n504_), .A2(KEYINPUT68), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n548_), .A2(new_n541_), .A3(new_n549_), .A4(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G57gat), .B(G64gat), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n552_), .A2(KEYINPUT11), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(KEYINPUT11), .ZN(new_n554_));
  XOR2_X1   g353(.A(G71gat), .B(G78gat), .Z(new_n555_));
  NAND3_X1  g354(.A1(new_n553_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n554_), .A2(new_n555_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G231gat), .A2(G233gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT70), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n558_), .B(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(new_n482_), .ZN(new_n562_));
  XOR2_X1   g361(.A(G127gat), .B(G155gat), .Z(new_n563_));
  XNOR2_X1  g362(.A(G183gat), .B(G211gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT71), .B(KEYINPUT16), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT17), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n567_), .A2(new_n568_), .ZN(new_n570_));
  NOR3_X1   g369(.A1(new_n562_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n562_), .A2(new_n569_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n546_), .A2(new_n551_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT66), .ZN(new_n575_));
  INV_X1    g374(.A(new_n558_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT12), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n523_), .A2(new_n526_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G230gat), .A2(G233gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n522_), .A2(new_n558_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT65), .B(KEYINPUT12), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n582_), .B1(new_n524_), .B2(new_n576_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .A4(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n524_), .A2(new_n576_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n581_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n587_), .A2(G230gat), .A3(G233gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G120gat), .B(G148gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT5), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G176gat), .B(G204gat), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n590_), .B(new_n591_), .Z(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n585_), .A2(new_n588_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n593_), .B1(new_n585_), .B2(new_n588_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n575_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n585_), .A2(new_n588_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(new_n592_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n599_), .A2(KEYINPUT66), .A3(new_n594_), .ZN(new_n600_));
  XOR2_X1   g399(.A(KEYINPUT67), .B(KEYINPUT13), .Z(new_n601_));
  NAND3_X1  g400(.A1(new_n597_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n595_), .A2(new_n575_), .A3(new_n596_), .ZN(new_n603_));
  AOI21_X1  g402(.A(KEYINPUT66), .B1(new_n599_), .B2(new_n594_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT13), .ZN(new_n605_));
  OAI22_X1  g404(.A1(new_n603_), .A2(new_n604_), .B1(KEYINPUT67), .B2(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n574_), .B1(new_n602_), .B2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n503_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n314_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n609_), .A2(new_n477_), .A3(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT38), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n548_), .A2(new_n541_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n474_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n606_), .A2(new_n602_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n614_), .A2(new_n573_), .A3(new_n502_), .A4(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT98), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n617_), .A2(new_n610_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n612_), .B1(new_n618_), .B2(new_n477_), .ZN(G1324gat));
  NAND2_X1  g418(.A1(new_n441_), .A2(new_n451_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(G8gat), .B1(new_n616_), .B2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT39), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n609_), .A2(new_n620_), .A3(new_n476_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT40), .Z(G1325gat));
  AOI21_X1  g425(.A(new_n352_), .B1(new_n617_), .B2(new_n473_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT41), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n609_), .A2(new_n352_), .A3(new_n473_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1326gat));
  INV_X1    g429(.A(G22gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n286_), .B(KEYINPUT99), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n631_), .B1(new_n617_), .B2(new_n632_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT42), .Z(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n631_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT100), .Z(new_n636_));
  OAI21_X1  g435(.A(new_n634_), .B1(new_n608_), .B2(new_n636_), .ZN(G1327gat));
  INV_X1    g436(.A(new_n615_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n638_), .A2(new_n613_), .A3(new_n573_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(new_n503_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(G29gat), .B1(new_n641_), .B2(new_n610_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n546_), .A2(new_n551_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n644_), .A2(KEYINPUT43), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(new_n474_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n647_));
  INV_X1    g446(.A(new_n455_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n441_), .A2(new_n451_), .A3(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n471_), .A2(new_n286_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n473_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n452_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n647_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  OAI211_X1 g452(.A(KEYINPUT101), .B(new_n452_), .C1(new_n472_), .C2(new_n473_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n653_), .A2(new_n643_), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT102), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n655_), .A2(new_n656_), .A3(KEYINPUT43), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n656_), .B1(new_n655_), .B2(KEYINPUT43), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n646_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n638_), .A2(new_n573_), .A3(new_n501_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  OR2_X1    g460(.A1(KEYINPUT103), .A2(KEYINPUT44), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n610_), .A2(G29gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n642_), .B1(new_n663_), .B2(new_n664_), .ZN(G1328gat));
  INV_X1    g464(.A(G36gat), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n641_), .A2(new_n666_), .A3(new_n620_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT45), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n663_), .A2(new_n620_), .ZN(new_n669_));
  OAI211_X1 g468(.A(KEYINPUT46), .B(new_n668_), .C1(new_n669_), .C2(new_n666_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT46), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n666_), .B1(new_n663_), .B2(new_n620_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n668_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n671_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n670_), .A2(new_n674_), .ZN(G1329gat));
  INV_X1    g474(.A(G43gat), .ZN(new_n676_));
  INV_X1    g475(.A(new_n473_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n676_), .B1(new_n640_), .B2(new_n677_), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT104), .Z(new_n679_));
  NOR2_X1   g478(.A1(new_n677_), .A2(new_n676_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n663_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT47), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n681_), .B(new_n682_), .ZN(G1330gat));
  AOI21_X1  g482(.A(G50gat), .B1(new_n641_), .B2(new_n632_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n287_), .A2(G50gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n663_), .B2(new_n685_), .ZN(G1331gat));
  NAND4_X1  g485(.A1(new_n614_), .A2(new_n573_), .A3(new_n501_), .A4(new_n638_), .ZN(new_n687_));
  INV_X1    g486(.A(G57gat), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n687_), .A2(new_n688_), .A3(new_n314_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n474_), .A2(new_n501_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT105), .Z(new_n691_));
  INV_X1    g490(.A(new_n574_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n691_), .A2(new_n638_), .A3(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n314_), .B1(new_n693_), .B2(KEYINPUT106), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n694_), .B1(KEYINPUT106), .B2(new_n693_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n689_), .B1(new_n695_), .B2(new_n688_), .ZN(G1332gat));
  OAI21_X1  g495(.A(G64gat), .B1(new_n687_), .B2(new_n621_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT48), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n621_), .A2(G64gat), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n698_), .B1(new_n693_), .B2(new_n699_), .ZN(G1333gat));
  NOR2_X1   g499(.A1(new_n677_), .A2(G71gat), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT108), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n693_), .A2(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(G71gat), .B1(new_n687_), .B2(new_n677_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT107), .Z(new_n705_));
  AOI21_X1  g504(.A(new_n703_), .B1(new_n705_), .B2(KEYINPUT49), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n706_), .B1(KEYINPUT49), .B2(new_n705_), .ZN(G1334gat));
  INV_X1    g506(.A(new_n632_), .ZN(new_n708_));
  OAI21_X1  g507(.A(G78gat), .B1(new_n687_), .B2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT50), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n708_), .A2(G78gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n710_), .B1(new_n693_), .B2(new_n711_), .ZN(G1335gat));
  INV_X1    g511(.A(new_n613_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n573_), .ZN(new_n714_));
  AND4_X1   g513(.A1(new_n713_), .A2(new_n691_), .A3(new_n714_), .A4(new_n638_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n715_), .A2(new_n517_), .A3(new_n610_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n638_), .A2(new_n714_), .A3(new_n501_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n659_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n659_), .A2(new_n718_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n717_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n721_), .A2(new_n610_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n716_), .B1(new_n722_), .B2(new_n517_), .ZN(G1336gat));
  NAND3_X1  g522(.A1(new_n715_), .A2(new_n518_), .A3(new_n620_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n721_), .A2(new_n620_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n725_), .B2(new_n518_), .ZN(G1337gat));
  INV_X1    g525(.A(G99gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n727_), .B1(new_n721_), .B2(new_n473_), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n715_), .A2(new_n473_), .A3(new_n514_), .ZN(new_n729_));
  OR3_X1    g528(.A1(new_n728_), .A2(KEYINPUT51), .A3(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(KEYINPUT51), .B1(new_n728_), .B2(new_n729_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1338gat));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n717_), .A2(new_n286_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n659_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(G106gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n733_), .B1(new_n659_), .B2(new_n734_), .ZN(new_n737_));
  OAI21_X1  g536(.A(KEYINPUT111), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n659_), .A2(new_n734_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT110), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT111), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n740_), .A2(new_n741_), .A3(G106gat), .A4(new_n735_), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n738_), .A2(KEYINPUT52), .A3(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT52), .ZN(new_n744_));
  OAI211_X1 g543(.A(KEYINPUT111), .B(new_n744_), .C1(new_n736_), .C2(new_n737_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n715_), .A2(new_n515_), .A3(new_n287_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(KEYINPUT53), .B1(new_n743_), .B2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n738_), .A2(KEYINPUT52), .A3(new_n742_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT53), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n749_), .A2(new_n750_), .A3(new_n745_), .A4(new_n746_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n748_), .A2(new_n751_), .ZN(G1339gat));
  AOI21_X1  g551(.A(KEYINPUT113), .B1(new_n607_), .B2(new_n501_), .ZN(new_n753_));
  AND4_X1   g552(.A1(KEYINPUT113), .A2(new_n615_), .A3(new_n692_), .A4(new_n501_), .ZN(new_n754_));
  OAI21_X1  g553(.A(KEYINPUT112), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n615_), .A2(new_n692_), .A3(new_n501_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT113), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n607_), .A2(KEYINPUT113), .A3(new_n501_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT112), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n758_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n755_), .A2(KEYINPUT54), .A3(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(KEYINPUT54), .B1(new_n755_), .B2(new_n761_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n501_), .A2(new_n595_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT56), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n583_), .B1(new_n522_), .B2(new_n558_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n580_), .B1(new_n768_), .B2(new_n579_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n585_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n768_), .A2(KEYINPUT55), .A3(new_n580_), .A4(new_n579_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n593_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n767_), .B1(new_n773_), .B2(KEYINPUT114), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n775_));
  AOI211_X1 g574(.A(new_n775_), .B(new_n593_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n774_), .A2(new_n776_), .ZN(new_n777_));
  AOI22_X1  g576(.A1(new_n777_), .A2(KEYINPUT115), .B1(KEYINPUT56), .B2(new_n773_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT115), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n779_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n766_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n492_), .A2(new_n496_), .A3(new_n500_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n491_), .A2(new_n495_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n495_), .B1(new_n483_), .B2(new_n487_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n500_), .B1(new_n784_), .B2(new_n494_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n782_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT116), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n782_), .A2(new_n786_), .A3(KEYINPUT116), .ZN(new_n790_));
  AOI211_X1 g589(.A(new_n603_), .B(new_n604_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n791_));
  OAI211_X1 g590(.A(KEYINPUT57), .B(new_n613_), .C1(new_n781_), .C2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT57), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n771_), .A2(new_n772_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n592_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n775_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n773_), .A2(KEYINPUT114), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n796_), .A2(KEYINPUT115), .A3(new_n767_), .A4(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n773_), .A2(KEYINPUT56), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n780_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n791_), .B1(new_n800_), .B2(new_n765_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n793_), .B1(new_n801_), .B2(new_n713_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n595_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n795_), .A2(new_n767_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n799_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n803_), .A2(new_n805_), .A3(KEYINPUT58), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT58), .B1(new_n803_), .B2(new_n805_), .ZN(new_n808_));
  OR3_X1    g607(.A1(new_n807_), .A2(new_n644_), .A3(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n792_), .A2(new_n802_), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n714_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n764_), .A2(new_n811_), .ZN(new_n812_));
  NOR4_X1   g611(.A1(new_n620_), .A2(new_n314_), .A3(new_n287_), .A4(new_n677_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(G113gat), .B1(new_n815_), .B2(new_n502_), .ZN(new_n816_));
  OR2_X1    g615(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n817_));
  NAND2_X1  g616(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n814_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n812_), .A2(KEYINPUT117), .A3(KEYINPUT59), .A4(new_n813_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n501_), .A2(KEYINPUT118), .ZN(new_n822_));
  MUX2_X1   g621(.A(KEYINPUT118), .B(new_n822_), .S(G113gat), .Z(new_n823_));
  AOI21_X1  g622(.A(new_n816_), .B1(new_n821_), .B2(new_n823_), .ZN(G1340gat));
  INV_X1    g623(.A(KEYINPUT60), .ZN(new_n825_));
  AOI21_X1  g624(.A(G120gat), .B1(new_n638_), .B2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n826_), .B1(new_n825_), .B2(G120gat), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n812_), .A2(new_n813_), .A3(new_n827_), .ZN(new_n828_));
  XOR2_X1   g627(.A(new_n828_), .B(KEYINPUT119), .Z(new_n829_));
  AOI21_X1  g628(.A(new_n615_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n830_));
  INV_X1    g629(.A(G120gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n829_), .B1(new_n830_), .B2(new_n831_), .ZN(G1341gat));
  INV_X1    g631(.A(G127gat), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n815_), .A2(new_n833_), .A3(new_n573_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n714_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(new_n833_), .ZN(G1342gat));
  INV_X1    g635(.A(G134gat), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n815_), .A2(new_n837_), .A3(new_n713_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n644_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n839_), .B2(new_n837_), .ZN(G1343gat));
  XNOR2_X1  g639(.A(KEYINPUT121), .B(G141gat), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n620_), .A2(new_n314_), .A3(new_n286_), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n807_), .A2(new_n644_), .A3(new_n808_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n613_), .B1(new_n781_), .B2(new_n791_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(new_n793_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n573_), .B1(new_n845_), .B2(new_n792_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n755_), .A2(new_n761_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n755_), .A2(KEYINPUT54), .A3(new_n761_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n677_), .B(new_n842_), .C1(new_n846_), .C2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n473_), .B1(new_n764_), .B2(new_n811_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n855_), .A2(KEYINPUT120), .A3(new_n842_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n841_), .B1(new_n857_), .B2(new_n502_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n841_), .ZN(new_n859_));
  AOI211_X1 g658(.A(new_n501_), .B(new_n859_), .C1(new_n854_), .C2(new_n856_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n858_), .A2(new_n860_), .ZN(G1344gat));
  XNOR2_X1  g660(.A(KEYINPUT122), .B(G148gat), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n862_), .B1(new_n857_), .B2(new_n638_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n862_), .ZN(new_n864_));
  AOI211_X1 g663(.A(new_n615_), .B(new_n864_), .C1(new_n854_), .C2(new_n856_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n863_), .A2(new_n865_), .ZN(G1345gat));
  NOR2_X1   g665(.A1(new_n852_), .A2(new_n853_), .ZN(new_n867_));
  AOI21_X1  g666(.A(KEYINPUT120), .B1(new_n855_), .B2(new_n842_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n573_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(KEYINPUT61), .B(G155gat), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n870_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n857_), .A2(new_n573_), .A3(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n873_), .ZN(G1346gat));
  NAND2_X1  g673(.A1(new_n857_), .A2(new_n713_), .ZN(new_n875_));
  INV_X1    g674(.A(G162gat), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n643_), .A2(G162gat), .ZN(new_n877_));
  XOR2_X1   g676(.A(new_n877_), .B(KEYINPUT123), .Z(new_n878_));
  AOI22_X1  g677(.A1(new_n875_), .A2(new_n876_), .B1(new_n857_), .B2(new_n878_), .ZN(G1347gat));
  XNOR2_X1  g678(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n621_), .A2(new_n367_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n882_), .B1(new_n764_), .B2(new_n811_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n883_), .A2(new_n502_), .A3(new_n708_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n880_), .B1(new_n884_), .B2(KEYINPUT22), .ZN(new_n885_));
  OAI21_X1  g684(.A(G169gat), .B1(new_n884_), .B2(new_n880_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(G169gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n888_), .B2(new_n885_), .ZN(G1348gat));
  NAND2_X1  g688(.A1(new_n812_), .A2(new_n881_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n632_), .ZN(new_n891_));
  AOI21_X1  g690(.A(G176gat), .B1(new_n891_), .B2(new_n638_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n890_), .A2(new_n287_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n638_), .A2(G176gat), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n892_), .B1(new_n893_), .B2(new_n894_), .ZN(G1349gat));
  NAND3_X1  g694(.A1(new_n883_), .A2(new_n286_), .A3(new_n573_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(KEYINPUT125), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(G183gat), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n896_), .A2(KEYINPUT125), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n714_), .B1(new_n322_), .B2(new_n381_), .ZN(new_n900_));
  AOI22_X1  g699(.A1(new_n898_), .A2(new_n899_), .B1(new_n891_), .B2(new_n900_), .ZN(G1350gat));
  NAND3_X1  g700(.A1(new_n891_), .A2(new_n320_), .A3(new_n713_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n890_), .A2(new_n644_), .A3(new_n632_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n377_), .B2(new_n903_), .ZN(G1351gat));
  NAND3_X1  g703(.A1(new_n855_), .A2(new_n648_), .A3(new_n620_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n905_), .A2(new_n501_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(new_n219_), .ZN(G1352gat));
  NOR2_X1   g706(.A1(new_n905_), .A2(new_n615_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(new_n257_), .ZN(G1353gat));
  NOR2_X1   g708(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n910_));
  AND2_X1   g709(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n911_));
  NOR4_X1   g710(.A1(new_n905_), .A2(new_n714_), .A3(new_n910_), .A4(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n910_), .B1(new_n905_), .B2(new_n714_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT126), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  OAI211_X1 g714(.A(KEYINPUT126), .B(new_n910_), .C1(new_n905_), .C2(new_n714_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n912_), .B1(new_n915_), .B2(new_n916_), .ZN(G1354gat));
  XNOR2_X1  g716(.A(KEYINPUT127), .B(G218gat), .ZN(new_n918_));
  NOR3_X1   g717(.A1(new_n905_), .A2(new_n644_), .A3(new_n918_), .ZN(new_n919_));
  OR2_X1    g718(.A1(new_n905_), .A2(new_n613_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n919_), .B1(new_n920_), .B2(new_n918_), .ZN(G1355gat));
endmodule


