//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 0 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 0 1 1 0 0 1 0 0 1 0 1 1 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n866_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n896_, new_n897_, new_n899_, new_n900_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT15), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G29gat), .B(G36gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G43gat), .B(G50gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n206_), .A2(new_n208_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n203_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  XOR2_X1   g011(.A(new_n204_), .B(new_n205_), .Z(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(new_n207_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(KEYINPUT15), .A3(new_n209_), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G99gat), .A2(G106gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT6), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT7), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n222_), .B(new_n223_), .C1(G99gat), .C2(G106gat), .ZN(new_n224_));
  INV_X1    g023(.A(G99gat), .ZN(new_n225_));
  INV_X1    g024(.A(G106gat), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n225_), .B(new_n226_), .C1(KEYINPUT64), .C2(KEYINPUT7), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n221_), .B1(new_n224_), .B2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G85gat), .A2(G92gat), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G85gat), .A2(G92gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT65), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G85gat), .ZN(new_n233_));
  INV_X1    g032(.A(G92gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n236_), .A3(new_n229_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT8), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n232_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n228_), .A2(new_n239_), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n232_), .A2(new_n237_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n224_), .A2(new_n227_), .A3(new_n242_), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n219_), .A2(new_n220_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n242_), .B1(new_n224_), .B2(new_n227_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n241_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n240_), .B1(new_n247_), .B2(KEYINPUT8), .ZN(new_n248_));
  XOR2_X1   g047(.A(KEYINPUT10), .B(G99gat), .Z(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(new_n226_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n235_), .A2(KEYINPUT9), .A3(new_n229_), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n229_), .A2(KEYINPUT9), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n250_), .A2(new_n251_), .A3(new_n252_), .A4(new_n244_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n248_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n216_), .A2(KEYINPUT73), .A3(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n258_), .B1(new_n248_), .B2(new_n254_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n214_), .A2(new_n209_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n224_), .A2(new_n227_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT66), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n262_), .A2(new_n244_), .A3(new_n243_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n238_), .B1(new_n263_), .B2(new_n241_), .ZN(new_n264_));
  OAI211_X1 g063(.A(KEYINPUT67), .B(new_n253_), .C1(new_n264_), .C2(new_n240_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n259_), .A2(new_n260_), .A3(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT73), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n212_), .A2(new_n215_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n267_), .B1(new_n268_), .B2(new_n255_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n257_), .A2(new_n266_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G232gat), .A2(G233gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT34), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT35), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n274_), .A2(KEYINPUT75), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(KEYINPUT75), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n275_), .B(new_n276_), .C1(KEYINPUT35), .C2(new_n272_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n277_), .B1(new_n216_), .B2(new_n256_), .ZN(new_n278_));
  AOI22_X1  g077(.A1(new_n270_), .A2(new_n274_), .B1(new_n266_), .B2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G190gat), .B(G218gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT74), .ZN(new_n281_));
  XOR2_X1   g080(.A(G134gat), .B(G162gat), .Z(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT36), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n279_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n283_), .A2(KEYINPUT36), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n279_), .A2(KEYINPUT76), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(KEYINPUT76), .B1(new_n279_), .B2(new_n288_), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n202_), .B(new_n286_), .C1(new_n290_), .C2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT76), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n270_), .A2(new_n274_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n278_), .A2(new_n266_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n293_), .B1(new_n296_), .B2(new_n287_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n284_), .B(KEYINPUT77), .ZN(new_n298_));
  AOI22_X1  g097(.A1(new_n297_), .A2(new_n289_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n292_), .B1(new_n299_), .B2(new_n202_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G57gat), .B(G64gat), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n301_), .A2(KEYINPUT11), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(KEYINPUT11), .ZN(new_n303_));
  XOR2_X1   g102(.A(G71gat), .B(G78gat), .Z(new_n304_));
  NAND3_X1  g103(.A1(new_n302_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n303_), .A2(new_n304_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G231gat), .A2(G233gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT79), .ZN(new_n310_));
  INV_X1    g109(.A(G1gat), .ZN(new_n311_));
  INV_X1    g110(.A(G8gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT14), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT78), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT78), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n315_), .B(KEYINPUT14), .C1(new_n311_), .C2(new_n312_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G15gat), .B(G22gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n314_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(G1gat), .B(G8gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n310_), .B(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(G127gat), .B(G155gat), .Z(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT16), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G183gat), .B(G211gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT17), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n322_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n326_), .A2(new_n327_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n322_), .A2(new_n328_), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n300_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G230gat), .A2(G233gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n259_), .A2(new_n307_), .A3(new_n265_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n307_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n247_), .A2(KEYINPUT8), .ZN(new_n341_));
  INV_X1    g140(.A(new_n240_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(KEYINPUT67), .B1(new_n343_), .B2(new_n253_), .ZN(new_n344_));
  NOR3_X1   g143(.A1(new_n248_), .A2(new_n258_), .A3(new_n254_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n340_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n339_), .B1(new_n346_), .B2(KEYINPUT68), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n307_), .B1(new_n259_), .B2(new_n265_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT68), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n338_), .B1(new_n347_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT12), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n346_), .A2(new_n352_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n340_), .B(KEYINPUT12), .C1(new_n248_), .C2(new_n254_), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n339_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n353_), .A2(new_n355_), .A3(new_n337_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n351_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G120gat), .B(G148gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT5), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G176gat), .B(G204gat), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n359_), .B(new_n360_), .Z(new_n361_));
  XOR2_X1   g160(.A(new_n361_), .B(KEYINPUT69), .Z(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n357_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n361_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n351_), .A2(new_n356_), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n336_), .B1(new_n365_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT13), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n364_), .B(new_n367_), .C1(KEYINPUT70), .C2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n334_), .A2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT80), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G71gat), .B(G99gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(G43gat), .ZN(new_n377_));
  XOR2_X1   g176(.A(KEYINPUT89), .B(KEYINPUT30), .Z(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  XOR2_X1   g178(.A(G127gat), .B(G134gat), .Z(new_n380_));
  XNOR2_X1  g179(.A(G113gat), .B(G120gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n379_), .B(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G183gat), .A2(G190gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT23), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT86), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT87), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n385_), .B(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n387_), .B1(KEYINPUT23), .B2(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(G169gat), .A2(G176gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT85), .ZN(new_n392_));
  INV_X1    g191(.A(G169gat), .ZN(new_n393_));
  INV_X1    g192(.A(G176gat), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT24), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT25), .B(G183gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT26), .B(G190gat), .ZN(new_n399_));
  AOI22_X1  g198(.A1(new_n392_), .A2(new_n397_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n392_), .A2(KEYINPUT24), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n390_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G227gat), .A2(G233gat), .ZN(new_n403_));
  INV_X1    g202(.A(G15gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n385_), .A2(KEYINPUT23), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n389_), .A2(KEYINPUT23), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n407_), .B1(new_n408_), .B2(KEYINPUT88), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n409_), .B1(KEYINPUT88), .B2(new_n408_), .ZN(new_n410_));
  OR2_X1    g209(.A1(G183gat), .A2(G190gat), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT22), .B(G169gat), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n395_), .B1(new_n413_), .B2(new_n394_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n402_), .B(new_n406_), .C1(new_n412_), .C2(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n415_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n402_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n405_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT31), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n416_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n420_), .B1(new_n416_), .B2(new_n419_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n384_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n423_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(new_n421_), .A3(new_n383_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n424_), .A2(new_n426_), .A3(KEYINPUT90), .ZN(new_n427_));
  AOI21_X1  g226(.A(KEYINPUT90), .B1(new_n424_), .B2(new_n426_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT3), .ZN(new_n431_));
  INV_X1    g230(.A(G141gat), .ZN(new_n432_));
  INV_X1    g231(.A(G148gat), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G141gat), .A2(G148gat), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT2), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n434_), .A2(new_n437_), .A3(new_n438_), .A4(new_n439_), .ZN(new_n440_));
  AND2_X1   g239(.A1(G155gat), .A2(G162gat), .ZN(new_n441_));
  NOR2_X1   g240(.A1(G155gat), .A2(G162gat), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n440_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT91), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT1), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n442_), .B1(new_n441_), .B2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n448_), .B1(new_n447_), .B2(new_n441_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n432_), .A2(new_n433_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(new_n435_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n446_), .A2(new_n451_), .ZN(new_n452_));
  OR2_X1    g251(.A1(new_n452_), .A2(KEYINPUT29), .ZN(new_n453_));
  XOR2_X1   g252(.A(G22gat), .B(G50gat), .Z(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  AND2_X1   g254(.A1(KEYINPUT93), .A2(G228gat), .ZN(new_n456_));
  NOR2_X1   g255(.A1(KEYINPUT93), .A2(G228gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(G233gat), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  XOR2_X1   g257(.A(new_n458_), .B(G78gat), .Z(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(new_n226_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n455_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n454_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n453_), .B(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n460_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n461_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n452_), .A2(KEYINPUT29), .ZN(new_n467_));
  INV_X1    g266(.A(G197gat), .ZN(new_n468_));
  OR3_X1    g267(.A1(new_n468_), .A2(KEYINPUT94), .A3(G204gat), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT94), .B1(new_n468_), .B2(G204gat), .ZN(new_n470_));
  INV_X1    g269(.A(G204gat), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n469_), .B(new_n470_), .C1(G197gat), .C2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT21), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G211gat), .B(G218gat), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT95), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n475_), .B1(new_n468_), .B2(G204gat), .ZN(new_n476_));
  NOR3_X1   g275(.A1(new_n471_), .A2(KEYINPUT95), .A3(G197gat), .ZN(new_n477_));
  OAI22_X1  g276(.A1(new_n476_), .A2(new_n477_), .B1(new_n468_), .B2(G204gat), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n473_), .B(new_n474_), .C1(new_n478_), .C2(KEYINPUT21), .ZN(new_n479_));
  INV_X1    g278(.A(new_n474_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(KEYINPUT21), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n467_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n484_));
  XOR2_X1   g283(.A(new_n483_), .B(new_n484_), .Z(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n466_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n461_), .A2(new_n465_), .A3(new_n485_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n430_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT4), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT99), .B1(new_n452_), .B2(new_n382_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n493_), .B1(new_n382_), .B2(new_n452_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT99), .ZN(new_n495_));
  OR3_X1    g294(.A1(new_n452_), .A2(new_n495_), .A3(new_n382_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n492_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n452_), .A2(new_n492_), .A3(new_n382_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT101), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G225gat), .A2(G233gat), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n501_), .B(KEYINPUT100), .Z(new_n502_));
  NAND3_X1  g301(.A1(new_n498_), .A2(new_n500_), .A3(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(G1gat), .B(G29gat), .Z(new_n504_));
  XNOR2_X1  g303(.A(KEYINPUT102), .B(KEYINPUT0), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G57gat), .B(G85gat), .ZN(new_n507_));
  XOR2_X1   g306(.A(new_n506_), .B(new_n507_), .Z(new_n508_));
  NAND2_X1  g307(.A1(new_n494_), .A2(new_n496_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n501_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n503_), .A2(KEYINPUT33), .A3(new_n508_), .A4(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n508_), .B1(new_n509_), .B2(new_n502_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n500_), .A2(new_n501_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n512_), .B1(new_n513_), .B2(new_n497_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT104), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n512_), .B(KEYINPUT104), .C1(new_n497_), .C2(new_n513_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n511_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n500_), .A2(new_n502_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n508_), .B(new_n510_), .C1(new_n519_), .C2(new_n497_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(KEYINPUT103), .B1(new_n521_), .B2(KEYINPUT33), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT103), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT33), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n520_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n518_), .B1(new_n522_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G226gat), .A2(G233gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT19), .ZN(new_n528_));
  INV_X1    g327(.A(new_n482_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT96), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n410_), .A2(new_n530_), .A3(new_n401_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n530_), .B1(new_n410_), .B2(new_n401_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n400_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n390_), .A2(new_n411_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n415_), .B1(new_n534_), .B2(KEYINPUT97), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n535_), .B1(KEYINPUT97), .B2(new_n534_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n529_), .B1(new_n533_), .B2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n402_), .B1(new_n412_), .B2(new_n415_), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT20), .B1(new_n538_), .B2(new_n482_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n528_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT98), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n533_), .A2(new_n529_), .A3(new_n536_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT20), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n543_), .B1(new_n538_), .B2(new_n482_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n528_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT98), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n548_), .B(new_n528_), .C1(new_n537_), .C2(new_n539_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n541_), .A2(new_n547_), .A3(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G8gat), .B(G36gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT18), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G64gat), .B(G92gat), .ZN(new_n553_));
  XOR2_X1   g352(.A(new_n552_), .B(new_n553_), .Z(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n550_), .A2(new_n555_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n541_), .A2(new_n547_), .A3(new_n554_), .A4(new_n549_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n526_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n503_), .A2(new_n510_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n508_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(new_n520_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n554_), .A2(KEYINPUT32), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n550_), .A2(new_n566_), .ZN(new_n567_));
  OR3_X1    g366(.A1(new_n537_), .A2(new_n539_), .A3(new_n528_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n568_), .B1(new_n546_), .B2(new_n545_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n569_), .A2(KEYINPUT105), .A3(new_n566_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(KEYINPUT105), .B1(new_n569_), .B2(new_n566_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n564_), .B(new_n567_), .C1(new_n571_), .C2(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n491_), .B1(new_n560_), .B2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n489_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n424_), .A2(new_n426_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n577_), .A2(new_n488_), .A3(new_n487_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n564_), .B1(new_n575_), .B2(new_n578_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n557_), .A2(KEYINPUT106), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n557_), .A2(KEYINPUT106), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT27), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n582_), .B1(new_n569_), .B2(new_n555_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n580_), .A2(new_n581_), .A3(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(KEYINPUT107), .B(KEYINPUT27), .Z(new_n585_));
  OAI21_X1  g384(.A(new_n585_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n586_));
  AND3_X1   g385(.A1(new_n579_), .A2(new_n584_), .A3(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n574_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT81), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n260_), .A2(new_n589_), .A3(new_n320_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n589_), .B1(new_n260_), .B2(new_n320_), .ZN(new_n591_));
  OAI22_X1  g390(.A1(new_n590_), .A2(new_n591_), .B1(new_n320_), .B2(new_n260_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G229gat), .A2(G233gat), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n212_), .A2(new_n321_), .A3(new_n215_), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n596_), .B(new_n593_), .C1(new_n590_), .C2(new_n591_), .ZN(new_n597_));
  XOR2_X1   g396(.A(G113gat), .B(G141gat), .Z(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT82), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G169gat), .B(G197gat), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n599_), .B(new_n600_), .Z(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n595_), .A2(new_n597_), .A3(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT83), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT83), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n595_), .A2(new_n605_), .A3(new_n597_), .A4(new_n602_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n595_), .A2(new_n597_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(new_n601_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT84), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n588_), .A2(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n564_), .B(KEYINPUT108), .Z(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n614_), .A2(G1gat), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n375_), .A2(new_n612_), .A3(new_n615_), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n616_), .A2(KEYINPUT109), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(KEYINPUT109), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n617_), .A2(KEYINPUT38), .A3(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(KEYINPUT38), .B1(new_n617_), .B2(new_n618_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n564_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n286_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n588_), .A2(new_n623_), .ZN(new_n624_));
  AOI22_X1  g423(.A1(new_n604_), .A2(new_n606_), .B1(new_n608_), .B2(new_n601_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n373_), .A2(new_n625_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n624_), .A2(KEYINPUT110), .A3(new_n333_), .A4(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT110), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n579_), .A2(new_n584_), .A3(new_n586_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n571_), .A2(new_n572_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n567_), .A2(new_n564_), .ZN(new_n631_));
  AOI22_X1  g430(.A1(new_n630_), .A2(new_n631_), .B1(new_n526_), .B2(new_n559_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n629_), .B1(new_n632_), .B2(new_n491_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(new_n622_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n626_), .A2(new_n333_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n628_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n621_), .B1(new_n627_), .B2(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n637_), .A2(new_n311_), .ZN(new_n638_));
  OR3_X1    g437(.A1(new_n619_), .A2(new_n620_), .A3(new_n638_), .ZN(G1324gat));
  NAND2_X1  g438(.A1(new_n584_), .A2(new_n586_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n375_), .A2(new_n312_), .A3(new_n612_), .A4(new_n640_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT111), .Z(new_n642_));
  NAND4_X1  g441(.A1(new_n624_), .A2(new_n640_), .A3(new_n333_), .A4(new_n626_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(G8gat), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT39), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n643_), .A2(KEYINPUT39), .A3(G8gat), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n642_), .A2(KEYINPUT40), .A3(new_n646_), .A4(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT40), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n647_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n641_), .B(KEYINPUT111), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n649_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n648_), .A2(new_n652_), .ZN(G1325gat));
  NAND4_X1  g452(.A1(new_n375_), .A2(new_n404_), .A3(new_n612_), .A4(new_n429_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n430_), .B1(new_n627_), .B2(new_n636_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n655_), .A2(new_n404_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n656_), .A2(KEYINPUT41), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n656_), .A2(KEYINPUT41), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n654_), .B1(new_n657_), .B2(new_n658_), .ZN(G1326gat));
  INV_X1    g458(.A(G22gat), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n375_), .A2(new_n660_), .A3(new_n612_), .A4(new_n489_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n490_), .B1(new_n627_), .B2(new_n636_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(new_n660_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT42), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n662_), .A2(KEYINPUT42), .A3(new_n660_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n661_), .B1(new_n665_), .B2(new_n666_), .ZN(G1327gat));
  INV_X1    g466(.A(new_n611_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n622_), .A2(new_n333_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n372_), .A2(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n633_), .A2(new_n668_), .A3(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(G29gat), .B1(new_n672_), .B2(new_n564_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n626_), .A2(new_n332_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n300_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n675_), .B1(new_n574_), .B2(new_n587_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT43), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT43), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n678_), .B(new_n675_), .C1(new_n574_), .C2(new_n587_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n674_), .B1(new_n677_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT44), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n681_), .A2(G29gat), .A3(new_n613_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n680_), .A2(KEYINPUT44), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n673_), .B1(new_n682_), .B2(new_n684_), .ZN(G1328gat));
  INV_X1    g484(.A(KEYINPUT46), .ZN(new_n686_));
  INV_X1    g485(.A(G36gat), .ZN(new_n687_));
  INV_X1    g486(.A(new_n640_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n680_), .B2(KEYINPUT44), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n687_), .B1(new_n684_), .B2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(KEYINPUT112), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT112), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n640_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n672_), .A2(new_n687_), .A3(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT45), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n695_), .B(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n686_), .B1(new_n690_), .B2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n681_), .A2(new_n640_), .ZN(new_n699_));
  OAI21_X1  g498(.A(G36gat), .B1(new_n699_), .B2(new_n683_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n695_), .B(KEYINPUT45), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n700_), .A2(KEYINPUT46), .A3(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n698_), .A2(new_n702_), .ZN(G1329gat));
  XOR2_X1   g502(.A(KEYINPUT113), .B(G43gat), .Z(new_n704_));
  OAI21_X1  g503(.A(new_n704_), .B1(new_n671_), .B2(new_n430_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT114), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n705_), .B(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n681_), .A2(G43gat), .A3(new_n577_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n707_), .B1(new_n708_), .B2(new_n683_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT47), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT47), .ZN(new_n711_));
  OAI211_X1 g510(.A(new_n707_), .B(new_n711_), .C1(new_n708_), .C2(new_n683_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(G1330gat));
  AOI21_X1  g512(.A(G50gat), .B1(new_n672_), .B2(new_n489_), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n681_), .A2(G50gat), .A3(new_n489_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n715_), .B2(new_n684_), .ZN(G1331gat));
  NOR3_X1   g515(.A1(new_n668_), .A2(new_n372_), .A3(new_n332_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n624_), .A2(new_n564_), .A3(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(G57gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(KEYINPUT115), .B1(new_n588_), .B2(new_n610_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT115), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n633_), .A2(new_n721_), .A3(new_n625_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n334_), .A2(new_n372_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n614_), .A2(G57gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n719_), .B1(new_n725_), .B2(new_n726_), .ZN(G1332gat));
  NAND3_X1  g526(.A1(new_n624_), .A2(new_n694_), .A3(new_n717_), .ZN(new_n728_));
  XOR2_X1   g527(.A(KEYINPUT116), .B(KEYINPUT48), .Z(new_n729_));
  AND3_X1   g528(.A1(new_n728_), .A2(G64gat), .A3(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n728_), .B2(G64gat), .ZN(new_n731_));
  INV_X1    g530(.A(new_n694_), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n732_), .A2(G64gat), .ZN(new_n733_));
  OAI22_X1  g532(.A1(new_n730_), .A2(new_n731_), .B1(new_n725_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT117), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n734_), .B(new_n735_), .ZN(G1333gat));
  NAND3_X1  g535(.A1(new_n624_), .A2(new_n429_), .A3(new_n717_), .ZN(new_n737_));
  XOR2_X1   g536(.A(KEYINPUT118), .B(KEYINPUT49), .Z(new_n738_));
  AND3_X1   g537(.A1(new_n737_), .A2(G71gat), .A3(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n737_), .B2(G71gat), .ZN(new_n740_));
  OR2_X1    g539(.A1(new_n430_), .A2(G71gat), .ZN(new_n741_));
  OAI22_X1  g540(.A1(new_n739_), .A2(new_n740_), .B1(new_n725_), .B2(new_n741_), .ZN(G1334gat));
  NAND3_X1  g541(.A1(new_n624_), .A2(new_n489_), .A3(new_n717_), .ZN(new_n743_));
  XOR2_X1   g542(.A(KEYINPUT119), .B(KEYINPUT50), .Z(new_n744_));
  AND3_X1   g543(.A1(new_n743_), .A2(G78gat), .A3(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n743_), .B2(G78gat), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n490_), .A2(G78gat), .ZN(new_n747_));
  OAI22_X1  g546(.A1(new_n745_), .A2(new_n746_), .B1(new_n725_), .B2(new_n747_), .ZN(G1335gat));
  NAND2_X1  g547(.A1(new_n373_), .A2(new_n669_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n720_), .B2(new_n722_), .ZN(new_n750_));
  AOI21_X1  g549(.A(G85gat), .B1(new_n750_), .B2(new_n613_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n373_), .A2(new_n625_), .A3(new_n332_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(new_n677_), .B2(new_n679_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT120), .Z(new_n754_));
  NOR2_X1   g553(.A1(new_n621_), .A2(new_n233_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(G1336gat));
  AOI21_X1  g555(.A(G92gat), .B1(new_n750_), .B2(new_n640_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n732_), .A2(new_n234_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n754_), .B2(new_n758_), .ZN(G1337gat));
  NAND2_X1  g558(.A1(new_n753_), .A2(new_n429_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(G99gat), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n577_), .A2(new_n249_), .ZN(new_n762_));
  AOI22_X1  g561(.A1(new_n750_), .A2(new_n762_), .B1(KEYINPUT121), .B2(KEYINPUT51), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(KEYINPUT121), .A2(KEYINPUT51), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT122), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n764_), .B(new_n766_), .ZN(G1338gat));
  NAND3_X1  g566(.A1(new_n750_), .A2(new_n226_), .A3(new_n489_), .ZN(new_n768_));
  AOI211_X1 g567(.A(KEYINPUT52), .B(new_n226_), .C1(new_n753_), .C2(new_n489_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n677_), .A2(new_n679_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n752_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n489_), .A3(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n770_), .B1(new_n773_), .B2(G106gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n768_), .B1(new_n769_), .B2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT53), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n777_), .B(new_n768_), .C1(new_n769_), .C2(new_n774_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(G1339gat));
  NOR3_X1   g578(.A1(new_n614_), .A2(new_n640_), .A3(new_n578_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n781_), .A2(KEYINPUT59), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n625_), .A2(new_n368_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n337_), .B1(new_n353_), .B2(new_n355_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n356_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n339_), .B(new_n354_), .C1(new_n348_), .C2(KEYINPUT12), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n787_), .A2(new_n785_), .A3(new_n338_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n786_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT56), .B1(new_n790_), .B2(new_n363_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT56), .ZN(new_n792_));
  AOI211_X1 g591(.A(new_n792_), .B(new_n362_), .C1(new_n786_), .C2(new_n789_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n783_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n592_), .A2(new_n593_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n596_), .B(new_n594_), .C1(new_n590_), .C2(new_n591_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n601_), .A3(new_n796_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n607_), .B(new_n797_), .C1(new_n365_), .C2(new_n368_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n623_), .B1(new_n794_), .B2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT57), .B1(new_n799_), .B2(KEYINPUT123), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT123), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT57), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n607_), .A2(new_n797_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n803_), .B1(new_n367_), .B2(new_n364_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n785_), .B1(new_n787_), .B2(new_n338_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n787_), .A2(new_n338_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n363_), .B1(new_n807_), .B2(new_n788_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n792_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n790_), .A2(KEYINPUT56), .A3(new_n363_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n804_), .B1(new_n811_), .B2(new_n783_), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n801_), .B(new_n802_), .C1(new_n812_), .C2(new_n623_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n803_), .A2(new_n368_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n811_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT58), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n811_), .A2(KEYINPUT58), .A3(new_n814_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n675_), .A3(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n800_), .A2(new_n813_), .A3(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT124), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n821_), .A3(new_n332_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n300_), .A2(new_n372_), .A3(new_n611_), .A4(new_n333_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n823_), .B(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n822_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n821_), .B1(new_n820_), .B2(new_n332_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n782_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n825_), .B1(new_n332_), .B2(new_n820_), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT59), .B1(new_n830_), .B2(new_n781_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(KEYINPUT125), .B(G113gat), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n611_), .A2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n829_), .A2(new_n831_), .A3(new_n833_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n820_), .A2(new_n332_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n610_), .B(new_n780_), .C1(new_n835_), .C2(new_n825_), .ZN(new_n836_));
  INV_X1    g635(.A(G113gat), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n834_), .A2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT126), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT126), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n834_), .A2(new_n841_), .A3(new_n838_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(G1340gat));
  NOR2_X1   g642(.A1(new_n830_), .A2(new_n781_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n372_), .A2(KEYINPUT60), .ZN(new_n845_));
  MUX2_X1   g644(.A(new_n845_), .B(KEYINPUT60), .S(G120gat), .Z(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT127), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n847_), .B(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n829_), .A2(new_n373_), .A3(new_n831_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(G120gat), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(G1341gat));
  INV_X1    g651(.A(G127gat), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n844_), .A2(new_n853_), .A3(new_n333_), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n829_), .A2(new_n333_), .A3(new_n831_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n853_), .ZN(G1342gat));
  NAND3_X1  g655(.A1(new_n829_), .A2(new_n675_), .A3(new_n831_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(G134gat), .ZN(new_n858_));
  INV_X1    g657(.A(new_n844_), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n622_), .A2(G134gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n858_), .B1(new_n859_), .B2(new_n860_), .ZN(G1343gat));
  NOR2_X1   g660(.A1(new_n830_), .A2(new_n575_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n694_), .A2(new_n614_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n862_), .A2(new_n610_), .A3(new_n863_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g664(.A1(new_n862_), .A2(new_n373_), .A3(new_n863_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g666(.A1(new_n862_), .A2(new_n333_), .A3(new_n863_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(KEYINPUT61), .B(G155gat), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n868_), .B(new_n869_), .ZN(G1346gat));
  INV_X1    g669(.A(G162gat), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n862_), .A2(new_n871_), .A3(new_n623_), .A4(new_n863_), .ZN(new_n872_));
  AND3_X1   g671(.A1(new_n862_), .A2(new_n675_), .A3(new_n863_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(new_n871_), .ZN(G1347gat));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n875_));
  NOR4_X1   g674(.A1(new_n732_), .A2(new_n430_), .A3(new_n489_), .A4(new_n613_), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n876_), .B(new_n610_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n875_), .B1(new_n878_), .B2(new_n393_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n877_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n413_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n879_), .A2(new_n880_), .A3(new_n881_), .ZN(G1348gat));
  NOR3_X1   g681(.A1(new_n732_), .A2(new_n430_), .A3(new_n613_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n883_), .A2(G176gat), .A3(new_n373_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n884_), .A2(new_n489_), .A3(new_n830_), .ZN(new_n885_));
  OR2_X1    g684(.A1(new_n827_), .A2(new_n828_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n886_), .A2(new_n373_), .A3(new_n876_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n885_), .B1(new_n887_), .B2(new_n394_), .ZN(G1349gat));
  AND2_X1   g687(.A1(new_n886_), .A2(new_n876_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n332_), .A2(new_n398_), .ZN(new_n890_));
  INV_X1    g689(.A(G183gat), .ZN(new_n891_));
  INV_X1    g690(.A(new_n830_), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n892_), .A2(new_n490_), .A3(new_n333_), .A4(new_n883_), .ZN(new_n893_));
  AOI22_X1  g692(.A1(new_n889_), .A2(new_n890_), .B1(new_n891_), .B2(new_n893_), .ZN(G1350gat));
  NAND3_X1  g693(.A1(new_n889_), .A2(new_n399_), .A3(new_n623_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n886_), .A2(new_n876_), .ZN(new_n896_));
  OAI21_X1  g695(.A(G190gat), .B1(new_n896_), .B2(new_n300_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n897_), .ZN(G1351gat));
  NOR2_X1   g697(.A1(new_n732_), .A2(new_n564_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n862_), .A2(new_n610_), .A3(new_n899_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g700(.A1(new_n862_), .A2(new_n373_), .A3(new_n899_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g702(.A1(new_n862_), .A2(new_n333_), .A3(new_n899_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n905_));
  AND2_X1   g704(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n904_), .A2(new_n905_), .A3(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n907_), .B1(new_n904_), .B2(new_n905_), .ZN(G1354gat));
  INV_X1    g707(.A(G218gat), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n862_), .A2(new_n909_), .A3(new_n623_), .A4(new_n899_), .ZN(new_n910_));
  AND3_X1   g709(.A1(new_n862_), .A2(new_n675_), .A3(new_n899_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n911_), .B2(new_n909_), .ZN(G1355gat));
endmodule


