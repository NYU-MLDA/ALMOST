//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n644_, new_n645_, new_n646_, new_n647_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n847_, new_n848_, new_n849_, new_n851_, new_n852_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n886_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n911_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT68), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT11), .ZN(new_n205_));
  XOR2_X1   g004(.A(G71gat), .B(G78gat), .Z(new_n206_));
  OR2_X1    g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n202_), .B(KEYINPUT68), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT11), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n205_), .A2(new_n210_), .A3(new_n206_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n207_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT77), .ZN(new_n213_));
  INV_X1    g012(.A(G1gat), .ZN(new_n214_));
  INV_X1    g013(.A(G8gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT14), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n216_), .A2(KEYINPUT75), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(KEYINPUT75), .ZN(new_n218_));
  XOR2_X1   g017(.A(G15gat), .B(G22gat), .Z(new_n219_));
  NOR3_X1   g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(G1gat), .B(G8gat), .Z(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G231gat), .A2(G233gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n213_), .A2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G127gat), .B(G155gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT16), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G183gat), .B(G211gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n229_), .A2(KEYINPUT17), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(KEYINPUT17), .ZN(new_n231_));
  NOR3_X1   g030(.A1(new_n225_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n232_), .B1(new_n224_), .B2(new_n213_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT70), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n212_), .B(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n236_), .A2(new_n224_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n224_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n230_), .B(KEYINPUT76), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n233_), .A2(new_n240_), .ZN(new_n241_));
  XOR2_X1   g040(.A(new_n241_), .B(KEYINPUT78), .Z(new_n242_));
  INV_X1    g041(.A(KEYINPUT37), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n244_));
  XOR2_X1   g043(.A(G85gat), .B(G92gat), .Z(new_n245_));
  INV_X1    g044(.A(G99gat), .ZN(new_n246_));
  INV_X1    g045(.A(G106gat), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT65), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT7), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n246_), .B(new_n247_), .C1(new_n248_), .C2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n250_), .B1(KEYINPUT65), .B2(KEYINPUT7), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G99gat), .A2(G106gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT6), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n248_), .A2(new_n249_), .A3(new_n246_), .A4(new_n247_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n251_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n244_), .B(new_n245_), .C1(new_n255_), .C2(KEYINPUT66), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT8), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(KEYINPUT10), .B(G99gat), .Z(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT64), .B(G106gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n245_), .A2(KEYINPUT9), .ZN(new_n262_));
  INV_X1    g061(.A(G85gat), .ZN(new_n263_));
  INV_X1    g062(.A(G92gat), .ZN(new_n264_));
  OR3_X1    g063(.A1(new_n263_), .A2(new_n264_), .A3(KEYINPUT9), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n261_), .A2(new_n262_), .A3(new_n265_), .A4(new_n253_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n257_), .A2(KEYINPUT67), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n255_), .B(new_n245_), .C1(KEYINPUT66), .C2(new_n267_), .ZN(new_n268_));
  AND3_X1   g067(.A1(new_n258_), .A2(new_n266_), .A3(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G29gat), .B(G36gat), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n270_), .A2(KEYINPUT72), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(KEYINPUT72), .ZN(new_n272_));
  XOR2_X1   g071(.A(G43gat), .B(G50gat), .Z(new_n273_));
  OR3_X1    g072(.A1(new_n271_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n273_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n269_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT73), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n276_), .B(KEYINPUT15), .Z(new_n281_));
  XOR2_X1   g080(.A(new_n266_), .B(KEYINPUT69), .Z(new_n282_));
  NAND3_X1  g081(.A1(new_n282_), .A2(new_n268_), .A3(new_n258_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT35), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G232gat), .A2(G233gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT34), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  AOI22_X1  g086(.A1(new_n281_), .A2(new_n283_), .B1(new_n284_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n280_), .A2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n287_), .A2(new_n284_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(G190gat), .B(G218gat), .Z(new_n292_));
  XNOR2_X1  g091(.A(G134gat), .B(G162gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n295_), .A2(KEYINPUT36), .ZN(new_n296_));
  INV_X1    g095(.A(new_n290_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n280_), .A2(new_n297_), .A3(new_n288_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n291_), .A2(new_n296_), .A3(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n243_), .B1(new_n299_), .B2(KEYINPUT74), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n294_), .B(KEYINPUT36), .ZN(new_n301_));
  INV_X1    g100(.A(new_n298_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n297_), .B1(new_n280_), .B2(new_n288_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n301_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n299_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n300_), .A2(new_n305_), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n304_), .B(new_n299_), .C1(KEYINPUT74), .C2(new_n243_), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n242_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n235_), .A2(KEYINPUT12), .A3(new_n283_), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n269_), .A2(new_n212_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT12), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G230gat), .A2(G233gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n269_), .A2(new_n212_), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n310_), .A2(new_n313_), .A3(new_n314_), .A4(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n311_), .A2(new_n315_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n314_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G120gat), .B(G148gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT5), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G176gat), .B(G204gat), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n321_), .B(new_n322_), .Z(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n316_), .A2(new_n319_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n324_), .B1(new_n316_), .B2(new_n319_), .ZN(new_n327_));
  OR3_X1    g126(.A1(new_n326_), .A2(new_n327_), .A3(KEYINPUT13), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT13), .B1(new_n326_), .B2(new_n327_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT71), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n309_), .A2(new_n331_), .A3(KEYINPUT79), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n222_), .B(new_n276_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G229gat), .A2(G233gat), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n281_), .A2(new_n222_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n336_), .B1(new_n222_), .B2(new_n276_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n335_), .B1(new_n337_), .B2(new_n334_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT80), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G113gat), .B(G141gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G169gat), .B(G197gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n340_), .B(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n332_), .A2(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(KEYINPUT79), .B1(new_n309_), .B2(new_n331_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G127gat), .B(G134gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G113gat), .B(G120gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n351_), .B(KEYINPUT31), .Z(new_n352_));
  NOR2_X1   g151(.A1(new_n352_), .A2(KEYINPUT84), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(G183gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT25), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT25), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(G183gat), .ZN(new_n358_));
  INV_X1    g157(.A(G190gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT26), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT26), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(G190gat), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n356_), .A2(new_n358_), .A3(new_n360_), .A4(new_n362_), .ZN(new_n363_));
  OR2_X1    g162(.A1(G169gat), .A2(G176gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G169gat), .A2(G176gat), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n364_), .A2(KEYINPUT24), .A3(new_n365_), .ZN(new_n366_));
  OR3_X1    g165(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n363_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT23), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n369_), .A2(G183gat), .A3(G190gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G183gat), .A2(G190gat), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n371_), .A2(KEYINPUT81), .A3(KEYINPUT23), .ZN(new_n372_));
  AOI21_X1  g171(.A(KEYINPUT81), .B1(new_n371_), .B2(KEYINPUT23), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n370_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n368_), .A2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(KEYINPUT82), .B1(new_n371_), .B2(KEYINPUT23), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n370_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n355_), .A2(new_n359_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n369_), .A2(KEYINPUT82), .A3(G183gat), .A4(G190gat), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n377_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n365_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT22), .B(G169gat), .ZN(new_n382_));
  INV_X1    g181(.A(G176gat), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n381_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n380_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n375_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT30), .ZN(new_n387_));
  XOR2_X1   g186(.A(G71gat), .B(G99gat), .Z(new_n388_));
  NAND2_X1  g187(.A1(G227gat), .A2(G233gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G15gat), .B(G43gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT83), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n390_), .B(new_n392_), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n387_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n387_), .A2(new_n393_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT85), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n396_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n354_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n394_), .A2(new_n395_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT85), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(new_n397_), .A3(new_n353_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n400_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT98), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT27), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G226gat), .A2(G233gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT19), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT20), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G211gat), .B(G218gat), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT21), .ZN(new_n413_));
  OR2_X1    g212(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n414_), .A2(KEYINPUT93), .A3(G204gat), .A4(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT91), .ZN(new_n417_));
  INV_X1    g216(.A(G204gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(KEYINPUT91), .A2(G204gat), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(G197gat), .A3(new_n420_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n416_), .A2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n414_), .A2(G204gat), .A3(new_n415_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT93), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n413_), .B1(new_n422_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(G197gat), .ZN(new_n427_));
  AND2_X1   g226(.A1(KEYINPUT91), .A2(G204gat), .ZN(new_n428_));
  NOR2_X1   g227(.A1(KEYINPUT91), .A2(G204gat), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n427_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT92), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  OAI211_X1 g231(.A(KEYINPUT92), .B(new_n427_), .C1(new_n428_), .C2(new_n429_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n415_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n418_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n432_), .A2(new_n433_), .A3(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n412_), .B1(new_n437_), .B2(KEYINPUT21), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT94), .B(KEYINPUT21), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n425_), .A2(new_n416_), .A3(new_n421_), .A4(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n426_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n374_), .A2(new_n378_), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n377_), .A2(new_n379_), .ZN(new_n443_));
  AOI22_X1  g242(.A1(new_n384_), .A2(new_n442_), .B1(new_n368_), .B2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n410_), .B1(new_n441_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT96), .ZN(new_n446_));
  AOI21_X1  g245(.A(G197gat), .B1(new_n419_), .B2(new_n420_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n436_), .B1(new_n447_), .B2(KEYINPUT92), .ZN(new_n448_));
  INV_X1    g247(.A(new_n433_), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT21), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n450_), .A2(new_n440_), .A3(new_n411_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n426_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n446_), .B1(new_n453_), .B2(new_n386_), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n368_), .A2(new_n374_), .B1(new_n380_), .B2(new_n384_), .ZN(new_n455_));
  AOI211_X1 g254(.A(KEYINPUT96), .B(new_n455_), .C1(new_n451_), .C2(new_n452_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n409_), .B(new_n445_), .C1(new_n454_), .C2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G8gat), .B(G36gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT18), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G64gat), .B(G92gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT20), .B1(new_n441_), .B2(new_n444_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n453_), .A2(new_n386_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n408_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n457_), .A2(new_n462_), .A3(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n462_), .B1(new_n457_), .B2(new_n465_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n406_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n457_), .A2(new_n462_), .A3(new_n465_), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n408_), .B(new_n445_), .C1(new_n454_), .C2(new_n456_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n409_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(new_n461_), .A3(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n469_), .A2(new_n472_), .A3(KEYINPUT27), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n468_), .A2(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(G155gat), .A2(G162gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G155gat), .A2(G162gat), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT86), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(KEYINPUT86), .A2(G155gat), .A3(G162gat), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n475_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NOR4_X1   g279(.A1(KEYINPUT87), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT87), .ZN(new_n482_));
  NOR2_X1   g281(.A1(G141gat), .A2(G148gat), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT3), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n482_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G141gat), .A2(G148gat), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n486_), .A2(KEYINPUT2), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n486_), .A2(KEYINPUT2), .ZN(new_n488_));
  OAI22_X1  g287(.A1(new_n481_), .A2(new_n485_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT88), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n480_), .B1(new_n489_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n483_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT1), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n478_), .A2(new_n495_), .A3(new_n479_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n475_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n495_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n486_), .B(new_n494_), .C1(new_n498_), .C2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n493_), .A2(new_n500_), .A3(new_n351_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n351_), .B1(new_n493_), .B2(new_n500_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G225gat), .A2(G233gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n503_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n507_), .A2(KEYINPUT4), .A3(new_n501_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT4), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n505_), .B1(new_n503_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n506_), .B1(new_n509_), .B2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G1gat), .B(G29gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT0), .ZN(new_n515_));
  INV_X1    g314(.A(G57gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(G85gat), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n513_), .A2(new_n519_), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n506_), .B(new_n518_), .C1(new_n509_), .C2(new_n512_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT29), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n523_), .B1(new_n493_), .B2(new_n500_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(G233gat), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT89), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n527_), .A2(G228gat), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(G228gat), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n526_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n453_), .A2(new_n525_), .A3(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n531_), .B1(new_n441_), .B2(new_n524_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G78gat), .B(G106gat), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n533_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n536_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(G22gat), .B(G50gat), .Z(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n493_), .A2(new_n500_), .A3(new_n523_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT28), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT28), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n493_), .A2(new_n500_), .A3(new_n545_), .A4(new_n523_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n542_), .B1(new_n544_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n544_), .A2(new_n546_), .A3(new_n542_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n550_), .B1(new_n539_), .B2(KEYINPUT95), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n540_), .A2(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n532_), .B1(new_n453_), .B2(new_n525_), .ZN(new_n553_));
  NOR3_X1   g352(.A1(new_n441_), .A2(new_n524_), .A3(new_n531_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n535_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n549_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n556_), .A2(new_n547_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT95), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n555_), .B(new_n537_), .C1(new_n557_), .C2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n522_), .B1(new_n552_), .B2(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n405_), .B1(new_n474_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n520_), .A2(new_n521_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n555_), .A2(new_n537_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n564_), .B(new_n550_), .C1(KEYINPUT95), .C2(new_n539_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n563_), .B1(new_n565_), .B2(new_n559_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n566_), .A2(KEYINPUT98), .A3(new_n468_), .A4(new_n473_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n562_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n565_), .A2(new_n559_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT33), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n521_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n508_), .A2(new_n511_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n506_), .A2(new_n518_), .A3(new_n572_), .A4(KEYINPUT33), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n508_), .B(new_n505_), .C1(KEYINPUT4), .C2(new_n507_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n504_), .A2(G225gat), .A3(G233gat), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n574_), .A2(new_n519_), .A3(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n571_), .A2(new_n573_), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT97), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n579_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n457_), .A2(new_n465_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n461_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n582_), .A2(KEYINPUT97), .A3(new_n469_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n578_), .A2(new_n580_), .A3(new_n583_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n470_), .A2(KEYINPUT32), .A3(new_n462_), .A4(new_n471_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n462_), .A2(KEYINPUT32), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n457_), .A2(new_n586_), .A3(new_n465_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n563_), .A2(new_n585_), .A3(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n569_), .B1(new_n584_), .B2(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n404_), .B1(new_n568_), .B2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n400_), .A2(new_n403_), .A3(new_n522_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT99), .ZN(new_n592_));
  AOI21_X1  g391(.A(KEYINPUT27), .B1(new_n582_), .B2(new_n469_), .ZN(new_n593_));
  AND3_X1   g392(.A1(new_n469_), .A2(new_n472_), .A3(KEYINPUT27), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n592_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n468_), .A2(KEYINPUT99), .A3(new_n473_), .ZN(new_n596_));
  AOI211_X1 g395(.A(new_n569_), .B(new_n591_), .C1(new_n595_), .C2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n590_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n348_), .A2(new_n599_), .ZN(new_n600_));
  NOR3_X1   g399(.A1(new_n600_), .A2(G1gat), .A3(new_n522_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT38), .Z(new_n602_));
  INV_X1    g401(.A(new_n588_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n466_), .A2(new_n467_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n577_), .B1(new_n604_), .B2(KEYINPUT97), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n603_), .B1(new_n605_), .B2(new_n580_), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n562_), .B(new_n567_), .C1(new_n606_), .C2(new_n569_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n597_), .B1(new_n607_), .B2(new_n404_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n345_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n330_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n608_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n305_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n241_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(G1gat), .B1(new_n615_), .B2(new_n522_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n602_), .A2(new_n616_), .ZN(G1324gat));
  INV_X1    g416(.A(KEYINPUT40), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n595_), .A2(new_n596_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n611_), .A2(new_n620_), .A3(new_n614_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(G8gat), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(KEYINPUT100), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT100), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n621_), .A2(new_n624_), .A3(G8gat), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n623_), .A2(KEYINPUT39), .A3(new_n625_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n620_), .A2(new_n215_), .ZN(new_n630_));
  OAI211_X1 g429(.A(new_n628_), .B(new_n629_), .C1(new_n600_), .C2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(KEYINPUT101), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n631_), .A2(KEYINPUT101), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n618_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n634_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n636_), .A2(KEYINPUT40), .A3(new_n632_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(G1325gat));
  OAI21_X1  g437(.A(G15gat), .B1(new_n615_), .B2(new_n404_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n639_), .A2(KEYINPUT41), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(KEYINPUT41), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n404_), .A2(G15gat), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n640_), .B(new_n641_), .C1(new_n600_), .C2(new_n642_), .ZN(G1326gat));
  INV_X1    g442(.A(new_n569_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G22gat), .B1(new_n615_), .B2(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT42), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n644_), .A2(G22gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n646_), .B1(new_n600_), .B2(new_n647_), .ZN(G1327gat));
  INV_X1    g447(.A(new_n242_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n649_), .A2(new_n305_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n650_), .A2(new_n611_), .ZN(new_n651_));
  AOI21_X1  g450(.A(G29gat), .B1(new_n651_), .B2(new_n563_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT44), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n306_), .A2(new_n307_), .ZN(new_n654_));
  OAI21_X1  g453(.A(KEYINPUT43), .B1(new_n608_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT43), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n599_), .A2(new_n656_), .A3(new_n308_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n610_), .A2(new_n609_), .ZN(new_n659_));
  AND4_X1   g458(.A1(KEYINPUT102), .A2(new_n658_), .A3(new_n659_), .A4(new_n242_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n649_), .B1(new_n655_), .B2(new_n657_), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT102), .B1(new_n661_), .B2(new_n659_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n653_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n658_), .A2(new_n659_), .A3(new_n242_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT102), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n661_), .A2(KEYINPUT102), .A3(new_n659_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n670_), .A2(KEYINPUT103), .A3(new_n653_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n665_), .A2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(KEYINPUT104), .B1(new_n666_), .B2(new_n653_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n661_), .A2(new_n674_), .A3(KEYINPUT44), .A4(new_n659_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n676_), .A2(G29gat), .A3(new_n563_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n652_), .B1(new_n672_), .B2(new_n677_), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT105), .Z(G1328gat));
  INV_X1    g478(.A(KEYINPUT46), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n680_), .A2(KEYINPUT106), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(KEYINPUT106), .ZN(new_n682_));
  INV_X1    g481(.A(G36gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n619_), .B1(new_n673_), .B2(new_n675_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n672_), .B2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n651_), .A2(new_n683_), .A3(new_n620_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT45), .Z(new_n687_));
  OAI211_X1 g486(.A(new_n681_), .B(new_n682_), .C1(new_n685_), .C2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT103), .B1(new_n670_), .B2(new_n653_), .ZN(new_n689_));
  AOI211_X1 g488(.A(new_n664_), .B(KEYINPUT44), .C1(new_n668_), .C2(new_n669_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n684_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(G36gat), .ZN(new_n692_));
  INV_X1    g491(.A(new_n687_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n692_), .A2(KEYINPUT106), .A3(new_n680_), .A4(new_n693_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n688_), .A2(new_n694_), .ZN(G1329gat));
  INV_X1    g494(.A(new_n404_), .ZN(new_n696_));
  AOI21_X1  g495(.A(G43gat), .B1(new_n651_), .B2(new_n696_), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n676_), .A2(G43gat), .A3(new_n696_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n672_), .B2(new_n698_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g499(.A(G50gat), .B1(new_n651_), .B2(new_n569_), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n676_), .A2(G50gat), .A3(new_n569_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n672_), .B2(new_n702_), .ZN(G1331gat));
  NOR2_X1   g502(.A1(new_n330_), .A2(new_n345_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  NOR4_X1   g504(.A1(new_n705_), .A2(new_n608_), .A3(new_n242_), .A4(new_n308_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G57gat), .B1(new_n706_), .B2(new_n563_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n331_), .A2(new_n608_), .A3(new_n345_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n708_), .A2(new_n305_), .A3(new_n649_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n563_), .A2(new_n710_), .A3(G57gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n711_), .B1(new_n710_), .B2(G57gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n707_), .B1(new_n709_), .B2(new_n712_), .ZN(G1332gat));
  INV_X1    g512(.A(G64gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n714_), .B1(new_n709_), .B2(new_n620_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT48), .Z(new_n716_));
  NAND3_X1  g515(.A1(new_n706_), .A2(new_n714_), .A3(new_n620_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1333gat));
  INV_X1    g517(.A(G71gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n719_), .B1(new_n709_), .B2(new_n696_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT49), .Z(new_n721_));
  NAND3_X1  g520(.A1(new_n706_), .A2(new_n719_), .A3(new_n696_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1334gat));
  INV_X1    g522(.A(G78gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n724_), .B1(new_n709_), .B2(new_n569_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT50), .Z(new_n726_));
  NAND3_X1  g525(.A1(new_n706_), .A2(new_n724_), .A3(new_n569_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1335gat));
  INV_X1    g527(.A(new_n658_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT108), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n649_), .A2(new_n705_), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n730_), .A2(new_n731_), .A3(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n731_), .B1(new_n730_), .B2(new_n732_), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(G85gat), .B1(new_n735_), .B2(new_n522_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n708_), .A2(new_n650_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n738_), .A2(new_n263_), .A3(new_n563_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n736_), .A2(new_n739_), .ZN(G1336gat));
  OAI21_X1  g539(.A(G92gat), .B1(new_n735_), .B2(new_n619_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n738_), .A2(new_n264_), .A3(new_n620_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1337gat));
  NAND3_X1  g542(.A1(new_n738_), .A2(new_n696_), .A3(new_n259_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n733_), .A2(new_n734_), .A3(new_n404_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n744_), .B1(new_n745_), .B2(new_n246_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT51), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT51), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n748_), .B(new_n744_), .C1(new_n745_), .C2(new_n246_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1338gat));
  NAND3_X1  g549(.A1(new_n738_), .A2(new_n569_), .A3(new_n260_), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT110), .Z(new_n752_));
  NOR2_X1   g551(.A1(new_n705_), .A2(new_n644_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n247_), .B1(new_n661_), .B2(new_n753_), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n754_), .A2(KEYINPUT52), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(KEYINPUT52), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n752_), .A2(new_n755_), .A3(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g557(.A(new_n344_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT113), .ZN(new_n760_));
  OR2_X1    g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n760_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n761_), .B(new_n762_), .C1(new_n334_), .C2(new_n337_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT114), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n764_), .B1(new_n343_), .B2(new_n338_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n765_), .A2(new_n326_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n316_), .B(KEYINPUT55), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n310_), .A2(new_n315_), .A3(new_n313_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n768_), .A2(new_n769_), .A3(new_n318_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n768_), .B2(new_n318_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT56), .B1(new_n772_), .B2(new_n323_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n773_), .A2(KEYINPUT115), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n772_), .A2(KEYINPUT56), .A3(new_n323_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n775_), .B1(new_n773_), .B2(KEYINPUT115), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n766_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT58), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  OAI211_X1 g578(.A(KEYINPUT58), .B(new_n766_), .C1(new_n774_), .C2(new_n776_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n308_), .A3(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n345_), .A2(new_n325_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n772_), .A2(new_n323_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT56), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n782_), .B1(new_n785_), .B2(new_n775_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n326_), .A2(new_n327_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n765_), .A2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n305_), .B1(new_n786_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT57), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT57), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n791_), .B(new_n305_), .C1(new_n786_), .C2(new_n788_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n781_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n613_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n610_), .A2(new_n345_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n309_), .A2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n796_), .B1(new_n798_), .B2(KEYINPUT54), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n309_), .A2(KEYINPUT111), .A3(new_n800_), .A4(new_n797_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n798_), .A2(KEYINPUT54), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n799_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n795_), .A2(new_n803_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n619_), .A2(new_n563_), .A3(new_n696_), .A4(new_n644_), .ZN(new_n805_));
  XOR2_X1   g604(.A(new_n805_), .B(KEYINPUT116), .Z(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(G113gat), .B1(new_n808_), .B2(new_n345_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(KEYINPUT59), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n649_), .B1(new_n781_), .B2(new_n793_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n803_), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT59), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n813_), .A2(new_n814_), .A3(new_n806_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n810_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n345_), .A2(G113gat), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(KEYINPUT117), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n809_), .B1(new_n817_), .B2(new_n819_), .ZN(G1340gat));
  INV_X1    g619(.A(KEYINPUT60), .ZN(new_n821_));
  INV_X1    g620(.A(G120gat), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n610_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n808_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT118), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n808_), .A2(KEYINPUT118), .A3(new_n824_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(G120gat), .B1(new_n816_), .B2(new_n331_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(G1341gat));
  INV_X1    g630(.A(G127gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n832_), .B1(new_n807_), .B2(new_n242_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT119), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n810_), .A2(G127gat), .A3(new_n241_), .A4(new_n815_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT119), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n836_), .B(new_n832_), .C1(new_n807_), .C2(new_n242_), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n834_), .A2(new_n835_), .A3(new_n837_), .ZN(G1342gat));
  INV_X1    g637(.A(G134gat), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n654_), .A2(new_n839_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(KEYINPUT121), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n839_), .B1(new_n807_), .B2(new_n305_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  OAI211_X1 g643(.A(KEYINPUT120), .B(new_n839_), .C1(new_n807_), .C2(new_n305_), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n817_), .A2(new_n841_), .B1(new_n844_), .B2(new_n845_), .ZN(G1343gat));
  NAND4_X1  g645(.A1(new_n619_), .A2(new_n563_), .A3(new_n404_), .A4(new_n569_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n847_), .B1(new_n795_), .B2(new_n803_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n345_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g649(.A(new_n331_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n851_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g652(.A1(new_n848_), .A2(new_n649_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(KEYINPUT61), .B(G155gat), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n854_), .B(new_n855_), .ZN(G1346gat));
  NAND3_X1  g655(.A1(new_n848_), .A2(G162gat), .A3(new_n308_), .ZN(new_n857_));
  AOI21_X1  g656(.A(G162gat), .B1(new_n848_), .B2(new_n612_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n857_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n860_), .B1(new_n859_), .B2(new_n858_), .ZN(G1347gat));
  NOR2_X1   g660(.A1(new_n619_), .A2(new_n591_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(new_n569_), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n345_), .B(new_n864_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(G169gat), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(KEYINPUT62), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT124), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT62), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n865_), .A2(KEYINPUT123), .A3(new_n869_), .A4(G169gat), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT123), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n871_), .B1(new_n866_), .B2(KEYINPUT62), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT124), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n866_), .A2(new_n873_), .A3(KEYINPUT62), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n868_), .A2(new_n870_), .A3(new_n872_), .A4(new_n874_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n813_), .A2(new_n864_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(new_n382_), .A3(new_n345_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(G1348gat));
  AOI21_X1  g677(.A(G176gat), .B1(new_n876_), .B2(new_n610_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n569_), .B1(new_n795_), .B2(new_n803_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n331_), .A2(new_n383_), .A3(new_n863_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n879_), .B1(new_n880_), .B2(new_n881_), .ZN(G1349gat));
  AOI21_X1  g681(.A(new_n613_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n880_), .A2(new_n649_), .A3(new_n862_), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n876_), .A2(new_n883_), .B1(new_n884_), .B2(new_n355_), .ZN(G1350gat));
  NAND4_X1  g684(.A1(new_n876_), .A2(new_n360_), .A3(new_n362_), .A4(new_n612_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n876_), .A2(new_n308_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n886_), .B1(new_n888_), .B2(new_n359_), .ZN(G1351gat));
  NOR3_X1   g688(.A1(new_n619_), .A2(new_n696_), .A3(new_n561_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n804_), .A2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n345_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT125), .B(G197gat), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1352gat));
  OAI21_X1  g694(.A(G204gat), .B1(new_n891_), .B2(new_n331_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT126), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n419_), .A2(new_n420_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n804_), .A2(new_n899_), .A3(new_n851_), .A4(new_n890_), .ZN(new_n900_));
  AND3_X1   g699(.A1(new_n896_), .A2(new_n897_), .A3(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n897_), .B1(new_n896_), .B2(new_n900_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1353gat));
  NAND2_X1  g702(.A1(new_n892_), .A2(new_n241_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n904_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n905_));
  XOR2_X1   g704(.A(KEYINPUT63), .B(G211gat), .Z(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n904_), .B2(new_n906_), .ZN(G1354gat));
  INV_X1    g706(.A(G218gat), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n892_), .A2(new_n908_), .A3(new_n612_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n892_), .A2(new_n308_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n909_), .B1(new_n911_), .B2(new_n908_), .ZN(G1355gat));
endmodule


