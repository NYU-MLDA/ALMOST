//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 0 0 1 0 0 0 1 0 1 0 1 1 0 1 0 1 0 1 0 0 1 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n898_, new_n900_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  AND2_X1   g001(.A1(new_n202_), .A2(KEYINPUT70), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(KEYINPUT70), .ZN(new_n204_));
  XOR2_X1   g003(.A(G43gat), .B(G50gat), .Z(new_n205_));
  OR3_X1    g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n205_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT15), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G15gat), .B(G22gat), .ZN(new_n210_));
  INV_X1    g009(.A(G1gat), .ZN(new_n211_));
  INV_X1    g010(.A(G8gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT14), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G1gat), .B(G8gat), .ZN(new_n215_));
  XOR2_X1   g014(.A(new_n214_), .B(new_n215_), .Z(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n209_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G229gat), .A2(G233gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n208_), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n218_), .B(new_n219_), .C1(new_n217_), .C2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n208_), .B(new_n216_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(KEYINPUT76), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n221_), .B1(new_n223_), .B2(new_n219_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G113gat), .B(G141gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G169gat), .B(G197gat), .ZN(new_n226_));
  XOR2_X1   g025(.A(new_n225_), .B(new_n226_), .Z(new_n227_));
  OR2_X1    g026(.A1(new_n227_), .A2(KEYINPUT77), .ZN(new_n228_));
  XOR2_X1   g027(.A(new_n224_), .B(new_n228_), .Z(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G228gat), .A2(G233gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT29), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G155gat), .A2(G162gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT1), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT1), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n236_), .A2(G155gat), .A3(G162gat), .ZN(new_n237_));
  OR2_X1    g036(.A1(G155gat), .A2(G162gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n235_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G141gat), .A2(G148gat), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(G141gat), .A2(G148gat), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n239_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT83), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n239_), .A2(KEYINPUT83), .A3(new_n243_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n238_), .A2(new_n234_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT84), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT2), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n240_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n250_), .B1(new_n240_), .B2(new_n251_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT3), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n242_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n249_), .B1(new_n254_), .B2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n233_), .B1(new_n248_), .B2(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(G211gat), .B(G218gat), .Z(new_n262_));
  NOR2_X1   g061(.A1(G197gat), .A2(G204gat), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G197gat), .A2(G204gat), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n262_), .A2(KEYINPUT21), .A3(new_n264_), .A4(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n264_), .A2(KEYINPUT21), .A3(new_n265_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT21), .ZN(new_n268_));
  AND2_X1   g067(.A1(G197gat), .A2(G204gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n268_), .B1(new_n269_), .B2(new_n263_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G211gat), .B(G218gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n267_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n266_), .A2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n232_), .B1(new_n261_), .B2(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT83), .B1(new_n239_), .B2(new_n243_), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n239_), .A2(KEYINPUT83), .A3(new_n243_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n260_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT29), .ZN(new_n278_));
  INV_X1    g077(.A(new_n273_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(new_n231_), .A3(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G78gat), .B(G106gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT85), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n274_), .A2(new_n280_), .A3(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G22gat), .B(G50gat), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NOR3_X1   g084(.A1(new_n277_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT28), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n258_), .A2(new_n257_), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n288_), .B(new_n256_), .C1(new_n253_), .C2(new_n252_), .ZN(new_n289_));
  AOI22_X1  g088(.A1(new_n246_), .A2(new_n247_), .B1(new_n289_), .B2(new_n249_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n287_), .B1(new_n290_), .B2(new_n233_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n285_), .B1(new_n286_), .B2(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT28), .B1(new_n277_), .B2(KEYINPUT29), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n290_), .A2(new_n287_), .A3(new_n233_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(new_n294_), .A3(new_n284_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n292_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT87), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n274_), .A2(new_n280_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n298_), .B1(new_n299_), .B2(new_n281_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n281_), .ZN(new_n301_));
  AOI211_X1 g100(.A(KEYINPUT87), .B(new_n301_), .C1(new_n274_), .C2(new_n280_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n283_), .B(new_n297_), .C1(new_n300_), .C2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n282_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n231_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n305_));
  AOI211_X1 g104(.A(new_n232_), .B(new_n273_), .C1(new_n277_), .C2(KEYINPUT29), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n304_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n283_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT86), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n308_), .A2(new_n309_), .A3(new_n296_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n309_), .B1(new_n308_), .B2(new_n296_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n303_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT88), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  OAI211_X1 g113(.A(KEYINPUT88), .B(new_n303_), .C1(new_n310_), .C2(new_n311_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(G8gat), .B(G36gat), .Z(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G64gat), .B(G92gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G226gat), .A2(G233gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT19), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G183gat), .A2(G190gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT23), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT23), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n327_), .A2(G183gat), .A3(G190gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  OR2_X1    g128(.A1(KEYINPUT78), .A2(G183gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(KEYINPUT78), .A2(G183gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n329_), .B1(new_n332_), .B2(G190gat), .ZN(new_n333_));
  INV_X1    g132(.A(G176gat), .ZN(new_n334_));
  INV_X1    g133(.A(G169gat), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT22), .B1(new_n335_), .B2(KEYINPUT81), .ZN(new_n336_));
  OR2_X1    g135(.A1(new_n335_), .A2(KEYINPUT22), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n334_), .B(new_n336_), .C1(new_n337_), .C2(KEYINPUT81), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G169gat), .A2(G176gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n333_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT26), .B(G190gat), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT25), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n342_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n341_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n335_), .A2(new_n334_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n346_), .A2(KEYINPUT24), .A3(new_n339_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT24), .ZN(new_n348_));
  NOR2_X1   g147(.A1(G169gat), .A2(G176gat), .ZN(new_n349_));
  AOI22_X1  g148(.A1(new_n347_), .A2(KEYINPUT79), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n339_), .A2(KEYINPUT24), .ZN(new_n351_));
  OR3_X1    g150(.A1(new_n351_), .A2(KEYINPUT79), .A3(new_n349_), .ZN(new_n352_));
  AND3_X1   g151(.A1(new_n325_), .A2(KEYINPUT80), .A3(KEYINPUT23), .ZN(new_n353_));
  AOI21_X1  g152(.A(KEYINPUT80), .B1(new_n325_), .B2(KEYINPUT23), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n328_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n345_), .A2(new_n350_), .A3(new_n352_), .A4(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n273_), .B1(new_n340_), .B2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT25), .B(G183gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n341_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n349_), .A2(new_n348_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n359_), .A2(new_n329_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT89), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n339_), .A2(new_n362_), .A3(KEYINPUT24), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n362_), .B1(new_n339_), .B2(KEYINPUT24), .ZN(new_n365_));
  NOR3_X1   g164(.A1(new_n364_), .A2(new_n365_), .A3(new_n349_), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n272_), .B(new_n266_), .C1(new_n361_), .C2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT22), .B(G169gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(new_n334_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n339_), .B(KEYINPUT91), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(G183gat), .A2(G190gat), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n371_), .B1(new_n355_), .B2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT20), .B1(new_n367_), .B2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n357_), .B1(new_n375_), .B2(KEYINPUT98), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT98), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n377_), .B(KEYINPUT20), .C1(new_n367_), .C2(new_n374_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n324_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n329_), .A2(new_n360_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n365_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(new_n346_), .A3(new_n363_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(new_n382_), .A3(new_n359_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n355_), .A2(new_n373_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n369_), .A2(new_n370_), .ZN(new_n385_));
  AOI22_X1  g184(.A1(new_n383_), .A2(KEYINPUT90), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  OR3_X1    g185(.A1(new_n361_), .A2(new_n366_), .A3(KEYINPUT90), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n273_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n356_), .A2(new_n340_), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT20), .B1(new_n389_), .B2(new_n279_), .ZN(new_n390_));
  NOR3_X1   g189(.A1(new_n388_), .A2(new_n390_), .A3(new_n323_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n321_), .B1(new_n379_), .B2(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n323_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n321_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n386_), .A2(new_n273_), .A3(new_n387_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n389_), .A2(new_n279_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n395_), .A2(KEYINPUT20), .A3(new_n324_), .A4(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n393_), .A2(new_n394_), .A3(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n392_), .A2(KEYINPUT27), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT27), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n393_), .A2(new_n394_), .A3(new_n397_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n394_), .B1(new_n393_), .B2(new_n397_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n400_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n399_), .A2(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n316_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(G1gat), .B(G29gat), .Z(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G57gat), .B(G85gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G225gat), .A2(G233gat), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(G134gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(G127gat), .ZN(new_n415_));
  INV_X1    g214(.A(G127gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(G134gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(G120gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(G113gat), .ZN(new_n420_));
  INV_X1    g219(.A(G113gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(G120gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n420_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n418_), .A2(new_n423_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n415_), .A2(new_n417_), .A3(new_n420_), .A4(new_n422_), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n424_), .A2(KEYINPUT82), .A3(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(KEYINPUT82), .B1(new_n424_), .B2(new_n425_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n277_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n413_), .B1(new_n428_), .B2(KEYINPUT4), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n424_), .A2(new_n425_), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n260_), .B(new_n430_), .C1(new_n275_), .C2(new_n276_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n426_), .A2(new_n427_), .ZN(new_n432_));
  OAI211_X1 g231(.A(KEYINPUT4), .B(new_n431_), .C1(new_n290_), .C2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT93), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT93), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n428_), .A2(new_n435_), .A3(KEYINPUT4), .A4(new_n431_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n429_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n428_), .A2(new_n431_), .A3(new_n412_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n411_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT99), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  OAI211_X1 g241(.A(KEYINPUT99), .B(new_n411_), .C1(new_n437_), .C2(new_n439_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n437_), .A2(new_n439_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n411_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n442_), .A2(new_n443_), .A3(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G227gat), .A2(G233gat), .ZN(new_n448_));
  INV_X1    g247(.A(G15gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT30), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n389_), .B(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(new_n432_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G71gat), .B(G99gat), .ZN(new_n454_));
  INV_X1    g253(.A(G43gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT31), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n453_), .B(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n447_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n406_), .A2(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n447_), .A2(new_n404_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n315_), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n274_), .A2(new_n280_), .A3(new_n282_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n282_), .B1(new_n274_), .B2(new_n280_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n296_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT86), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n308_), .A2(new_n309_), .A3(new_n296_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(KEYINPUT88), .B1(new_n469_), .B2(new_n303_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n462_), .B1(new_n463_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT100), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT100), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n316_), .A2(new_n473_), .A3(new_n462_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n463_), .A2(new_n470_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n394_), .A2(KEYINPUT32), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n393_), .A2(new_n397_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n476_), .B1(new_n477_), .B2(KEYINPUT97), .ZN(new_n478_));
  OR3_X1    g277(.A1(new_n379_), .A2(new_n391_), .A3(new_n476_), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n393_), .A2(KEYINPUT97), .A3(new_n397_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n478_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n447_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n428_), .A2(KEYINPUT95), .A3(new_n431_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(new_n413_), .ZN(new_n484_));
  AOI21_X1  g283(.A(KEYINPUT95), .B1(new_n428_), .B2(new_n431_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n411_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT96), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT96), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n488_), .B(new_n411_), .C1(new_n484_), .C2(new_n485_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n434_), .A2(new_n436_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n490_), .B(new_n412_), .C1(KEYINPUT4), .C2(new_n428_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n487_), .A2(new_n489_), .A3(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n401_), .A2(new_n402_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT33), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n494_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n495_));
  NOR4_X1   g294(.A1(new_n437_), .A2(KEYINPUT33), .A3(new_n439_), .A4(new_n411_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n492_), .B(new_n493_), .C1(new_n495_), .C2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n482_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n475_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n472_), .A2(new_n474_), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n458_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT101), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n461_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n458_), .ZN(new_n504_));
  AOI22_X1  g303(.A1(new_n471_), .A2(KEYINPUT100), .B1(new_n475_), .B2(new_n498_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n504_), .B1(new_n505_), .B2(new_n474_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT101), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n230_), .B1(new_n503_), .B2(new_n507_), .ZN(new_n508_));
  XOR2_X1   g307(.A(KEYINPUT10), .B(G99gat), .Z(new_n509_));
  INV_X1    g308(.A(G106gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(G85gat), .B(G92gat), .Z(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT9), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT9), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(G85gat), .A3(G92gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G99gat), .A2(G106gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT6), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT6), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n518_), .A2(G99gat), .A3(G106gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n511_), .A2(new_n513_), .A3(new_n515_), .A4(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT64), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT7), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n522_), .B(new_n523_), .C1(G99gat), .C2(G106gat), .ZN(new_n524_));
  INV_X1    g323(.A(G99gat), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n525_), .B(new_n510_), .C1(KEYINPUT64), .C2(KEYINPUT7), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n520_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT8), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n528_), .A2(new_n529_), .A3(new_n512_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT65), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n520_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n517_), .A2(new_n519_), .A3(KEYINPUT65), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(new_n527_), .A3(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n529_), .B1(new_n534_), .B2(new_n512_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT66), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n530_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n527_), .A2(new_n533_), .ZN(new_n538_));
  AOI21_X1  g337(.A(KEYINPUT65), .B1(new_n517_), .B2(new_n519_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n512_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT8), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n541_), .A2(KEYINPUT66), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n220_), .B(new_n521_), .C1(new_n537_), .C2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n521_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n530_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n545_), .B1(new_n541_), .B2(KEYINPUT66), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n535_), .A2(new_n536_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n544_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n543_), .B1(new_n209_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT35), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G232gat), .A2(G233gat), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT34), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n549_), .A2(KEYINPUT71), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n554_), .B1(new_n549_), .B2(KEYINPUT71), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n553_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n549_), .A2(KEYINPUT71), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(KEYINPUT34), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n549_), .A2(KEYINPUT71), .A3(new_n554_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n559_), .A2(new_n552_), .A3(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n551_), .B1(new_n557_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n557_), .A2(new_n561_), .A3(KEYINPUT35), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G190gat), .B(G218gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G134gat), .B(G162gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n567_), .A2(KEYINPUT36), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n563_), .A2(new_n564_), .A3(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n567_), .B(KEYINPUT36), .Z(new_n570_));
  AND3_X1   g369(.A1(new_n557_), .A2(new_n561_), .A3(KEYINPUT35), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n570_), .B1(new_n571_), .B2(new_n562_), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n569_), .A2(KEYINPUT37), .A3(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT72), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  OAI211_X1 g375(.A(KEYINPUT72), .B(new_n570_), .C1(new_n571_), .C2(new_n562_), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n576_), .A2(new_n577_), .A3(new_n569_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n574_), .B1(new_n578_), .B2(KEYINPUT37), .ZN(new_n579_));
  XOR2_X1   g378(.A(G57gat), .B(G64gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT67), .B(G71gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(G78gat), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT11), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n580_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n584_), .B1(new_n583_), .B2(new_n582_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n582_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n586_), .A2(KEYINPUT11), .A3(new_n580_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  AND2_X1   g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n590_), .A2(KEYINPUT73), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(KEYINPUT73), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n591_), .A2(new_n216_), .A3(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n216_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(KEYINPUT17), .B1(KEYINPUT68), .B2(KEYINPUT75), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n593_), .A2(new_n594_), .ZN(new_n598_));
  AOI21_X1  g397(.A(KEYINPUT75), .B1(new_n598_), .B2(KEYINPUT17), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT75), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT17), .ZN(new_n601_));
  OAI21_X1  g400(.A(KEYINPUT68), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n597_), .B1(new_n599_), .B2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G127gat), .B(G155gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G183gat), .B(G211gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  XOR2_X1   g405(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n603_), .A2(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(new_n601_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n595_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n579_), .A2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n521_), .B1(new_n537_), .B2(new_n542_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n588_), .B1(new_n614_), .B2(KEYINPUT12), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n614_), .A2(KEYINPUT68), .A3(KEYINPUT12), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G230gat), .A2(G233gat), .ZN(new_n618_));
  INV_X1    g417(.A(new_n588_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n617_), .B(new_n618_), .C1(new_n619_), .C2(new_n616_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n618_), .B1(new_n619_), .B2(new_n614_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n621_), .B1(new_n614_), .B2(new_n619_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(G120gat), .B(G148gat), .Z(new_n624_));
  XNOR2_X1  g423(.A(G176gat), .B(G204gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n623_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n623_), .A2(new_n629_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT13), .Z(new_n634_));
  AND3_X1   g433(.A1(new_n508_), .A2(new_n613_), .A3(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n635_), .A2(new_n211_), .A3(new_n447_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT38), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n638_), .B(KEYINPUT102), .Z(new_n639_));
  AOI211_X1 g438(.A(new_n578_), .B(new_n612_), .C1(new_n503_), .C2(new_n507_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n634_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n641_), .A2(new_n230_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n211_), .B1(new_n643_), .B2(new_n447_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n637_), .B2(new_n636_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n639_), .A2(new_n645_), .ZN(G1324gat));
  NAND3_X1  g445(.A1(new_n635_), .A2(new_n212_), .A3(new_n404_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT39), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n643_), .A2(new_n404_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n649_), .B2(G8gat), .ZN(new_n650_));
  AOI211_X1 g449(.A(KEYINPUT39), .B(new_n212_), .C1(new_n643_), .C2(new_n404_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n647_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT40), .Z(G1325gat));
  NAND2_X1  g452(.A1(new_n643_), .A2(new_n504_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(G15gat), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n655_), .A2(KEYINPUT41), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(KEYINPUT41), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n635_), .A2(new_n449_), .A3(new_n504_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT103), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n656_), .A2(new_n657_), .A3(new_n659_), .ZN(G1326gat));
  INV_X1    g459(.A(G22gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n661_), .B1(new_n643_), .B2(new_n316_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT42), .Z(new_n663_));
  NAND3_X1  g462(.A1(new_n635_), .A2(new_n661_), .A3(new_n316_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1327gat));
  NAND2_X1  g464(.A1(new_n612_), .A2(new_n578_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n666_), .A2(new_n641_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(new_n508_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n447_), .ZN(new_n669_));
  OR3_X1    g468(.A1(new_n668_), .A2(G29gat), .A3(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n576_), .A2(new_n577_), .A3(new_n569_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT37), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n573_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n503_), .B2(new_n507_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n671_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n461_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n678_), .B1(new_n506_), .B2(KEYINPUT101), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n501_), .A2(new_n502_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n579_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n681_), .A2(KEYINPUT104), .A3(KEYINPUT43), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n675_), .A2(new_n676_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n677_), .A2(new_n682_), .A3(new_n683_), .ZN(new_n684_));
  AOI22_X1  g483(.A1(new_n603_), .A2(new_n608_), .B1(new_n595_), .B2(new_n610_), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n685_), .A2(new_n641_), .A3(new_n230_), .ZN(new_n686_));
  AOI21_X1  g485(.A(KEYINPUT44), .B1(new_n684_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n684_), .A2(KEYINPUT44), .A3(new_n686_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n688_), .A2(new_n447_), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT105), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(G29gat), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n690_), .A2(KEYINPUT105), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n670_), .B1(new_n692_), .B2(new_n693_), .ZN(G1328gat));
  AND2_X1   g493(.A1(new_n667_), .A2(new_n508_), .ZN(new_n695_));
  INV_X1    g494(.A(G36gat), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n695_), .A2(KEYINPUT107), .A3(new_n696_), .A4(new_n404_), .ZN(new_n697_));
  XOR2_X1   g496(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n698_));
  INV_X1    g497(.A(KEYINPUT107), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n404_), .A2(new_n696_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n699_), .B1(new_n668_), .B2(new_n700_), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n697_), .A2(new_n698_), .A3(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n698_), .B1(new_n697_), .B2(new_n701_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n684_), .A2(KEYINPUT44), .A3(new_n686_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n404_), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n705_), .A2(new_n687_), .A3(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n704_), .B1(new_n707_), .B2(new_n696_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT46), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  OAI211_X1 g509(.A(KEYINPUT46), .B(new_n704_), .C1(new_n707_), .C2(new_n696_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1329gat));
  NOR4_X1   g511(.A1(new_n705_), .A2(new_n687_), .A3(new_n455_), .A4(new_n458_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n695_), .A2(new_n504_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n715_), .B2(new_n455_), .ZN(new_n716_));
  AOI211_X1 g515(.A(KEYINPUT108), .B(G43gat), .C1(new_n695_), .C2(new_n504_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(KEYINPUT47), .B1(new_n713_), .B2(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n705_), .A2(new_n687_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(G43gat), .A3(new_n504_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT47), .ZN(new_n722_));
  INV_X1    g521(.A(new_n718_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n721_), .A2(new_n722_), .A3(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n719_), .A2(new_n724_), .ZN(G1330gat));
  AOI21_X1  g524(.A(G50gat), .B1(new_n695_), .B2(new_n316_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n316_), .A2(G50gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n720_), .B2(new_n727_), .ZN(G1331gat));
  NAND2_X1  g527(.A1(new_n613_), .A2(new_n641_), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n729_), .A2(KEYINPUT109), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(KEYINPUT109), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n229_), .B1(new_n503_), .B2(new_n507_), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n730_), .A2(new_n731_), .A3(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(G57gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(new_n734_), .A3(new_n447_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n634_), .A2(new_n229_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n640_), .A2(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(G57gat), .B1(new_n737_), .B2(new_n669_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n735_), .A2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT110), .ZN(G1332gat));
  OAI21_X1  g539(.A(G64gat), .B1(new_n737_), .B2(new_n706_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT48), .ZN(new_n742_));
  INV_X1    g541(.A(G64gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n733_), .A2(new_n743_), .A3(new_n404_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1333gat));
  OAI21_X1  g544(.A(G71gat), .B1(new_n737_), .B2(new_n458_), .ZN(new_n746_));
  XOR2_X1   g545(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n747_));
  XNOR2_X1  g546(.A(new_n746_), .B(new_n747_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n458_), .A2(G71gat), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT112), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n733_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n748_), .A2(new_n751_), .ZN(G1334gat));
  OAI21_X1  g551(.A(G78gat), .B1(new_n737_), .B2(new_n475_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT50), .ZN(new_n754_));
  INV_X1    g553(.A(G78gat), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n733_), .A2(new_n755_), .A3(new_n316_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(G1335gat));
  NAND2_X1  g556(.A1(new_n736_), .A2(new_n612_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT113), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n684_), .A2(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n669_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n666_), .A2(new_n634_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n732_), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n669_), .A2(G85gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n761_), .B1(new_n763_), .B2(new_n764_), .ZN(G1336gat));
  OAI21_X1  g564(.A(G92gat), .B1(new_n760_), .B2(new_n706_), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n706_), .A2(G92gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n766_), .B1(new_n763_), .B2(new_n767_), .ZN(G1337gat));
  OAI21_X1  g567(.A(G99gat), .B1(new_n760_), .B2(new_n458_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n763_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n770_), .A2(new_n504_), .A3(new_n509_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n769_), .A2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n773_));
  MUX2_X1   g572(.A(KEYINPUT51), .B(new_n773_), .S(KEYINPUT115), .Z(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n775_), .B1(new_n772_), .B2(new_n773_), .ZN(G1338gat));
  NAND3_X1  g575(.A1(new_n770_), .A2(new_n510_), .A3(new_n316_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n684_), .A2(new_n759_), .A3(new_n316_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n778_), .A2(new_n779_), .A3(G106gat), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n778_), .B2(G106gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n777_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT53), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n784_), .B(new_n777_), .C1(new_n780_), .C2(new_n781_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(G1339gat));
  NOR3_X1   g585(.A1(new_n406_), .A2(new_n458_), .A3(new_n669_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT57), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n615_), .A2(new_n616_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n618_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n616_), .A2(new_n619_), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n789_), .A2(new_n790_), .A3(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n792_), .A2(KEYINPUT117), .A3(KEYINPUT55), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT117), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n794_), .B1(new_n620_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n620_), .A2(new_n795_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n790_), .B1(new_n789_), .B2(new_n791_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n793_), .A2(new_n796_), .A3(new_n797_), .A4(new_n798_), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n799_), .A2(KEYINPUT56), .A3(new_n628_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT56), .B1(new_n799_), .B2(new_n628_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n229_), .B(new_n630_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n227_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n224_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n219_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n803_), .B1(new_n223_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT118), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n219_), .B1(new_n208_), .B2(new_n216_), .ZN(new_n809_));
  AOI22_X1  g608(.A1(new_n806_), .A2(new_n807_), .B1(new_n218_), .B2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n804_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n802_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n672_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT119), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n788_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  AOI211_X1 g615(.A(KEYINPUT119), .B(KEYINPUT57), .C1(new_n813_), .C2(new_n672_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n799_), .A2(KEYINPUT56), .A3(new_n628_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT120), .ZN(new_n820_));
  INV_X1    g619(.A(new_n801_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT120), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n799_), .A2(new_n822_), .A3(KEYINPUT56), .A4(new_n628_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n820_), .A2(new_n821_), .A3(new_n823_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n811_), .A2(new_n630_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n824_), .A2(new_n825_), .A3(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n827_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n828_), .A2(new_n829_), .A3(new_n674_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n685_), .B1(new_n818_), .B2(new_n831_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n674_), .A2(new_n230_), .A3(new_n685_), .A4(new_n634_), .ZN(new_n833_));
  XOR2_X1   g632(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n834_));
  XNOR2_X1  g633(.A(new_n833_), .B(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n787_), .B1(new_n832_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n838_), .A2(new_n421_), .A3(new_n229_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n837_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n578_), .B1(new_n802_), .B2(new_n812_), .ZN(new_n842_));
  OAI21_X1  g641(.A(KEYINPUT57), .B1(new_n842_), .B2(KEYINPUT119), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n814_), .A2(new_n815_), .A3(new_n788_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n612_), .B1(new_n845_), .B2(new_n830_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n835_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n847_), .A2(KEYINPUT59), .A3(new_n787_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n230_), .B1(new_n841_), .B2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n839_), .B1(new_n849_), .B2(new_n421_), .ZN(G1340gat));
  OAI21_X1  g649(.A(new_n419_), .B1(new_n634_), .B2(KEYINPUT60), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n838_), .B(new_n851_), .C1(KEYINPUT60), .C2(new_n419_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n634_), .B1(new_n841_), .B2(new_n848_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n419_), .ZN(G1341gat));
  NAND3_X1  g653(.A1(new_n838_), .A2(new_n416_), .A3(new_n685_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n612_), .B1(new_n841_), .B2(new_n848_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(new_n416_), .ZN(G1342gat));
  NAND2_X1  g656(.A1(new_n579_), .A2(G134gat), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(KEYINPUT122), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n859_), .B1(new_n841_), .B2(new_n848_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n414_), .B1(new_n837_), .B2(new_n672_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT123), .B1(new_n860_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n859_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n848_), .ZN(new_n865_));
  AOI21_X1  g664(.A(KEYINPUT59), .B1(new_n847_), .B2(new_n787_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n864_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT123), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n867_), .A2(new_n868_), .A3(new_n861_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n863_), .A2(new_n869_), .ZN(G1343gat));
  INV_X1    g669(.A(new_n847_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n475_), .A2(new_n504_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n872_), .A2(new_n447_), .A3(new_n706_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(KEYINPUT124), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n871_), .A2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n229_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n641_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g678(.A1(new_n875_), .A2(new_n685_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(KEYINPUT61), .B(G155gat), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n880_), .B(new_n881_), .ZN(G1346gat));
  INV_X1    g681(.A(G162gat), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n875_), .A2(new_n883_), .A3(new_n578_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n871_), .A2(new_n674_), .A3(new_n874_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n883_), .B2(new_n885_), .ZN(G1347gat));
  NOR3_X1   g685(.A1(new_n316_), .A2(new_n460_), .A3(new_n706_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n847_), .A2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n229_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(G169gat), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT62), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n889_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n888_), .A2(new_n229_), .A3(new_n368_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n892_), .A2(new_n893_), .A3(new_n894_), .ZN(G1348gat));
  NAND2_X1  g694(.A1(new_n888_), .A2(new_n641_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g696(.A1(new_n888_), .A2(new_n685_), .ZN(new_n898_));
  MUX2_X1   g697(.A(new_n358_), .B(new_n332_), .S(new_n898_), .Z(G1350gat));
  NAND2_X1  g698(.A1(new_n888_), .A2(new_n579_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(G190gat), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n888_), .A2(new_n341_), .A3(new_n578_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1351gat));
  NOR2_X1   g702(.A1(new_n706_), .A2(new_n447_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n872_), .A2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n871_), .A2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n229_), .ZN(new_n907_));
  XOR2_X1   g706(.A(KEYINPUT125), .B(G197gat), .Z(new_n908_));
  XNOR2_X1  g707(.A(new_n907_), .B(new_n908_), .ZN(G1352gat));
  NAND2_X1  g708(.A1(new_n906_), .A2(new_n641_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(G204gat), .ZN(G1353gat));
  OR2_X1    g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  XNOR2_X1  g711(.A(KEYINPUT63), .B(G211gat), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n871_), .A2(new_n612_), .A3(new_n905_), .ZN(new_n914_));
  MUX2_X1   g713(.A(new_n912_), .B(new_n913_), .S(new_n914_), .Z(G1354gat));
  NAND4_X1  g714(.A1(new_n847_), .A2(new_n578_), .A3(new_n872_), .A4(new_n904_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(KEYINPUT126), .B(G218gat), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  NOR4_X1   g718(.A1(new_n871_), .A2(new_n674_), .A3(new_n905_), .A4(new_n917_), .ZN(new_n920_));
  OAI21_X1  g719(.A(KEYINPUT127), .B1(new_n919_), .B2(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n917_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n906_), .A2(new_n579_), .A3(new_n922_), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT127), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n923_), .A2(new_n924_), .A3(new_n918_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n921_), .A2(new_n925_), .ZN(G1355gat));
endmodule


