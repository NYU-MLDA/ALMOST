//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 0 0 0 0 1 0 1 1 0 1 0 1 1 0 0 0 1 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 1 0 0 0 1 1 1 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n673_, new_n674_, new_n675_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n885_, new_n886_, new_n887_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n202_));
  XOR2_X1   g001(.A(G197gat), .B(G204gat), .Z(new_n203_));
  AND2_X1   g002(.A1(KEYINPUT88), .A2(KEYINPUT21), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G211gat), .B(G218gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n203_), .A2(KEYINPUT21), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n203_), .A2(new_n204_), .A3(new_n206_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G141gat), .ZN(new_n213_));
  INV_X1    g012(.A(G148gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(KEYINPUT83), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n219_), .A2(KEYINPUT1), .ZN(new_n220_));
  INV_X1    g019(.A(G155gat), .ZN(new_n221_));
  INV_X1    g020(.A(G162gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(new_n222_), .A3(KEYINPUT82), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT82), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n224_), .B1(G155gat), .B2(G162gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n226_), .B1(new_n219_), .B2(KEYINPUT1), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n217_), .B1(new_n220_), .B2(new_n227_), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n218_), .A2(KEYINPUT83), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n218_), .A2(KEYINPUT83), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n223_), .B(new_n225_), .C1(new_n229_), .C2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT3), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n234_), .B1(G141gat), .B2(G148gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  AND3_X1   g035(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n237_));
  AOI21_X1  g036(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  AND3_X1   g038(.A1(new_n236_), .A2(new_n239_), .A3(KEYINPUT84), .ZN(new_n240_));
  AOI21_X1  g039(.A(KEYINPUT84), .B1(new_n236_), .B2(new_n239_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n232_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT85), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT85), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n244_), .B(new_n232_), .C1(new_n240_), .C2(new_n241_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n228_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT29), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n212_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT28), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n246_), .A2(new_n249_), .A3(new_n247_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n249_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n202_), .B(new_n248_), .C1(new_n251_), .C2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n248_), .A2(new_n202_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n252_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(new_n255_), .A3(new_n250_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(new_n256_), .ZN(new_n257_));
  OAI211_X1 g056(.A(KEYINPUT89), .B(new_n212_), .C1(new_n246_), .C2(new_n247_), .ZN(new_n258_));
  XOR2_X1   g057(.A(KEYINPUT87), .B(G233gat), .Z(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT86), .B(G228gat), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G78gat), .B(G106gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT90), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n258_), .A2(new_n264_), .A3(new_n261_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G22gat), .B(G50gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n266_), .A2(new_n267_), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n269_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n257_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n267_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n264_), .B1(new_n258_), .B2(new_n261_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n268_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n276_), .A2(new_n270_), .A3(new_n256_), .A4(new_n253_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n273_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G8gat), .B(G36gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G64gat), .B(G92gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(G169gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT23), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n286_), .A2(G183gat), .A3(G190gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT80), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n286_), .B1(G183gat), .B2(G190gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(KEYINPUT79), .B(G190gat), .Z(new_n291_));
  NOR2_X1   g090(.A1(new_n291_), .A2(G183gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n285_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(G169gat), .ZN(new_n296_));
  INV_X1    g095(.A(G176gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n295_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  OR3_X1    g097(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(G183gat), .ZN(new_n301_));
  INV_X1    g100(.A(G190gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT23), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n287_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n305_), .B1(new_n291_), .B2(KEYINPUT26), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n301_), .A2(KEYINPUT25), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n307_), .A2(KEYINPUT78), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(KEYINPUT78), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n301_), .A2(KEYINPUT25), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n308_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n300_), .B(new_n304_), .C1(new_n306_), .C2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n293_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n212_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n304_), .B1(G183gat), .B2(G190gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n285_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT26), .B(G190gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n317_), .A2(new_n307_), .A3(new_n310_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n316_), .B1(new_n290_), .B2(new_n319_), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n212_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n314_), .A2(new_n321_), .A3(KEYINPUT20), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G226gat), .A2(G233gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(KEYINPUT96), .B1(new_n322_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT20), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n328_), .B1(new_n212_), .B2(new_n320_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n293_), .A2(new_n312_), .A3(new_n211_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n331_), .A2(new_n326_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n327_), .A2(new_n332_), .ZN(new_n333_));
  NOR3_X1   g132(.A1(new_n331_), .A2(KEYINPUT96), .A3(new_n326_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n283_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT27), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT20), .B1(new_n212_), .B2(new_n320_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n211_), .B1(new_n293_), .B2(new_n312_), .ZN(new_n338_));
  NOR3_X1   g137(.A1(new_n337_), .A2(new_n338_), .A3(new_n326_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n325_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n283_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n336_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n340_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n314_), .A2(new_n321_), .A3(KEYINPUT20), .A4(new_n325_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n344_), .A2(new_n342_), .A3(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n283_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  AOI22_X1  g147(.A1(new_n335_), .A2(new_n343_), .B1(new_n336_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n278_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n228_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT84), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n233_), .A2(new_n235_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n238_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n353_), .B1(new_n354_), .B2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n236_), .A2(new_n239_), .A3(KEYINPUT84), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n244_), .B1(new_n360_), .B2(new_n232_), .ZN(new_n361_));
  AOI211_X1 g160(.A(KEYINPUT85), .B(new_n231_), .C1(new_n358_), .C2(new_n359_), .ZN(new_n362_));
  OAI211_X1 g161(.A(KEYINPUT93), .B(new_n352_), .C1(new_n361_), .C2(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G127gat), .B(G134gat), .Z(new_n364_));
  XOR2_X1   g163(.A(G113gat), .B(G120gat), .Z(new_n365_));
  XOR2_X1   g164(.A(new_n364_), .B(new_n365_), .Z(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n363_), .A2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n366_), .B1(new_n246_), .B2(KEYINPUT93), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT4), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G225gat), .A2(G233gat), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  OR3_X1    g171(.A1(new_n246_), .A2(KEYINPUT4), .A3(new_n367_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n370_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n371_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT95), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n363_), .A2(new_n367_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n246_), .A2(KEYINPUT93), .A3(new_n366_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n380_), .A2(KEYINPUT95), .A3(new_n371_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n374_), .A2(new_n377_), .A3(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(G1gat), .B(G29gat), .Z(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G57gat), .B(G85gat), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n385_), .B(new_n386_), .Z(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n382_), .A2(new_n388_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n374_), .A2(new_n377_), .A3(new_n387_), .A4(new_n381_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G227gat), .A2(G233gat), .ZN(new_n392_));
  INV_X1    g191(.A(G71gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(G99gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n313_), .B(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(new_n366_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G15gat), .B(G43gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT81), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT30), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT31), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n398_), .B(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n391_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n351_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT97), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n333_), .A2(new_n334_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n342_), .A2(KEYINPUT32), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  OR2_X1    g209(.A1(new_n341_), .A2(new_n409_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n370_), .A2(new_n371_), .A3(new_n373_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n387_), .B1(new_n380_), .B2(new_n372_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n348_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT33), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n388_), .A2(new_n416_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n374_), .A2(new_n377_), .A3(new_n381_), .A4(new_n417_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n415_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n390_), .A2(new_n416_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n391_), .A2(new_n412_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n407_), .B1(new_n421_), .B2(new_n278_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n391_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n423_), .A2(new_n278_), .A3(new_n349_), .ZN(new_n424_));
  NOR3_X1   g223(.A1(new_n271_), .A2(new_n272_), .A3(new_n257_), .ZN(new_n425_));
  AOI22_X1  g224(.A1(new_n276_), .A2(new_n270_), .B1(new_n256_), .B2(new_n253_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n390_), .A2(new_n416_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n415_), .A2(new_n418_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n389_), .A2(new_n390_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n431_));
  OAI211_X1 g230(.A(KEYINPUT97), .B(new_n427_), .C1(new_n430_), .C2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n422_), .A2(new_n424_), .A3(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n406_), .B1(new_n433_), .B2(new_n403_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G15gat), .B(G22gat), .ZN(new_n435_));
  INV_X1    g234(.A(G1gat), .ZN(new_n436_));
  INV_X1    g235(.A(G8gat), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT14), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n435_), .A2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G1gat), .B(G8gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G29gat), .B(G36gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G43gat), .B(G50gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  XOR2_X1   g243(.A(new_n441_), .B(new_n444_), .Z(new_n445_));
  NAND2_X1  g244(.A1(G229gat), .A2(G233gat), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n444_), .B(KEYINPUT15), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n441_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n441_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n447_), .B1(new_n450_), .B2(new_n444_), .ZN(new_n451_));
  AOI22_X1  g250(.A1(new_n445_), .A2(new_n447_), .B1(new_n449_), .B2(new_n451_), .ZN(new_n452_));
  XOR2_X1   g251(.A(G113gat), .B(G141gat), .Z(new_n453_));
  XNOR2_X1  g252(.A(G169gat), .B(G197gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  XOR2_X1   g254(.A(new_n455_), .B(KEYINPUT76), .Z(new_n456_));
  NOR3_X1   g255(.A1(new_n452_), .A2(KEYINPUT77), .A3(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n457_), .B1(new_n452_), .B2(new_n455_), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT77), .B1(new_n452_), .B2(new_n456_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n434_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT98), .ZN(new_n463_));
  XOR2_X1   g262(.A(G190gat), .B(G218gat), .Z(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT69), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G134gat), .B(G162gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  XOR2_X1   g266(.A(new_n467_), .B(KEYINPUT36), .Z(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT71), .ZN(new_n469_));
  XOR2_X1   g268(.A(G85gat), .B(G92gat), .Z(new_n470_));
  NOR2_X1   g269(.A1(G99gat), .A2(G106gat), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT7), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G99gat), .A2(G106gat), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT6), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n470_), .B1(new_n473_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT8), .ZN(new_n478_));
  OR3_X1    g277(.A1(new_n477_), .A2(KEYINPUT65), .A3(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT65), .B(KEYINPUT8), .ZN(new_n480_));
  XOR2_X1   g279(.A(KEYINPUT10), .B(G99gat), .Z(new_n481_));
  INV_X1    g280(.A(G106gat), .ZN(new_n482_));
  AOI22_X1  g281(.A1(KEYINPUT9), .A2(new_n470_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(G85gat), .ZN(new_n484_));
  INV_X1    g283(.A(G92gat), .ZN(new_n485_));
  NOR3_X1   g284(.A1(new_n484_), .A2(new_n485_), .A3(KEYINPUT9), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n476_), .A2(new_n486_), .ZN(new_n487_));
  AOI22_X1  g286(.A1(new_n477_), .A2(new_n480_), .B1(new_n483_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n479_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(new_n444_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n448_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G232gat), .A2(G233gat), .ZN(new_n493_));
  XOR2_X1   g292(.A(new_n493_), .B(KEYINPUT34), .Z(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT68), .B(KEYINPUT35), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n491_), .A2(new_n492_), .A3(new_n496_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n494_), .A2(new_n495_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n498_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n491_), .A2(new_n500_), .A3(new_n492_), .A4(new_n496_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n469_), .B1(KEYINPUT72), .B2(new_n502_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n502_), .A2(KEYINPUT72), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT73), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT37), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n467_), .A2(KEYINPUT36), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n499_), .A2(new_n501_), .A3(new_n508_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .A4(new_n509_), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n507_), .B(new_n509_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT73), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n469_), .A2(new_n502_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(KEYINPUT70), .A3(new_n509_), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT37), .B1(new_n509_), .B2(KEYINPUT70), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n513_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G57gat), .B(G64gat), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n520_), .A2(KEYINPUT11), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(KEYINPUT11), .ZN(new_n522_));
  XOR2_X1   g321(.A(G71gat), .B(G78gat), .Z(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n522_), .A2(new_n523_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  AND2_X1   g325(.A1(G231gat), .A2(G233gat), .ZN(new_n527_));
  XOR2_X1   g326(.A(new_n526_), .B(new_n527_), .Z(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT74), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(new_n441_), .ZN(new_n530_));
  XOR2_X1   g329(.A(G127gat), .B(G155gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G183gat), .B(G211gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT17), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n530_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n529_), .B(new_n450_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n535_), .A2(KEYINPUT17), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n519_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n490_), .A2(new_n526_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n526_), .B1(new_n479_), .B2(new_n488_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G230gat), .A2(G233gat), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n547_), .B(KEYINPUT64), .Z(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n546_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT66), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n544_), .A2(KEYINPUT67), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT12), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(KEYINPUT12), .B1(new_n544_), .B2(KEYINPUT67), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n554_), .A2(new_n555_), .A3(new_n548_), .A4(new_n543_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT66), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n546_), .A2(new_n557_), .A3(new_n549_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n551_), .A2(new_n556_), .A3(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G120gat), .B(G148gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT5), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G176gat), .B(G204gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n561_), .B(new_n562_), .Z(new_n563_));
  NAND2_X1  g362(.A1(new_n559_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n563_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n551_), .A2(new_n556_), .A3(new_n558_), .A4(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT13), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n564_), .A2(KEYINPUT13), .A3(new_n566_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n542_), .A2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n462_), .A2(new_n463_), .A3(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n432_), .A2(new_n424_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n391_), .A2(new_n412_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n419_), .A2(new_n420_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(KEYINPUT97), .B1(new_n577_), .B2(new_n427_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n403_), .B1(new_n574_), .B2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(new_n405_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n580_), .A2(new_n572_), .A3(new_n460_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT98), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n573_), .A2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n423_), .A2(G1gat), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n541_), .ZN(new_n586_));
  NOR3_X1   g385(.A1(new_n571_), .A2(new_n461_), .A3(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT101), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n505_), .A2(new_n509_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n580_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(G1gat), .B1(new_n590_), .B2(new_n423_), .ZN(new_n591_));
  XOR2_X1   g390(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n585_), .A2(new_n593_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n573_), .A2(new_n582_), .A3(new_n584_), .A4(new_n592_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT100), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n595_), .A2(new_n596_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n594_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT102), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(G1324gat));
  NAND4_X1  g400(.A1(new_n573_), .A2(new_n582_), .A3(new_n437_), .A4(new_n350_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT39), .ZN(new_n603_));
  INV_X1    g402(.A(new_n589_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n434_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n605_), .A2(new_n350_), .A3(new_n588_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n603_), .B1(new_n606_), .B2(G8gat), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n603_), .B(G8gat), .C1(new_n590_), .C2(new_n349_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n602_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT104), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT104), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n602_), .B(new_n612_), .C1(new_n607_), .C2(new_n609_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n611_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n614_), .B1(new_n611_), .B2(new_n613_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(G1325gat));
  OAI21_X1  g416(.A(G15gat), .B1(new_n590_), .B2(new_n403_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT41), .Z(new_n619_));
  INV_X1    g418(.A(G15gat), .ZN(new_n620_));
  INV_X1    g419(.A(new_n403_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n583_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n619_), .A2(new_n622_), .ZN(G1326gat));
  OAI21_X1  g422(.A(G22gat), .B1(new_n590_), .B2(new_n427_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT42), .ZN(new_n625_));
  INV_X1    g424(.A(G22gat), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n583_), .A2(new_n626_), .A3(new_n278_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(G1327gat));
  NOR3_X1   g427(.A1(new_n571_), .A2(new_n589_), .A3(new_n541_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n462_), .A2(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(G29gat), .B1(new_n630_), .B2(new_n391_), .ZN(new_n631_));
  OAI21_X1  g430(.A(KEYINPUT43), .B1(new_n434_), .B2(new_n519_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT43), .ZN(new_n633_));
  AOI22_X1  g432(.A1(new_n510_), .A2(new_n512_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n278_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n349_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  AOI22_X1  g436(.A1(new_n635_), .A2(KEYINPUT97), .B1(new_n637_), .B2(new_n423_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n621_), .B1(new_n638_), .B2(new_n422_), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n633_), .B(new_n634_), .C1(new_n639_), .C2(new_n406_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n632_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n571_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n642_), .A2(new_n460_), .A3(new_n586_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT105), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT44), .B1(new_n641_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT44), .ZN(new_n647_));
  AOI211_X1 g446(.A(new_n647_), .B(new_n644_), .C1(new_n632_), .C2(new_n640_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n391_), .A2(G29gat), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n631_), .B1(new_n649_), .B2(new_n650_), .ZN(G1328gat));
  INV_X1    g450(.A(G36gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n652_), .B1(new_n649_), .B2(new_n350_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n349_), .A2(G36gat), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n630_), .A2(KEYINPUT45), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT45), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n462_), .A2(new_n629_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n654_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n656_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n655_), .A2(new_n659_), .ZN(new_n660_));
  OAI211_X1 g459(.A(KEYINPUT106), .B(KEYINPUT46), .C1(new_n653_), .C2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT46), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n633_), .B1(new_n580_), .B2(new_n634_), .ZN(new_n663_));
  AOI211_X1 g462(.A(KEYINPUT43), .B(new_n519_), .C1(new_n579_), .C2(new_n405_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n645_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(new_n647_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n641_), .A2(KEYINPUT44), .A3(new_n645_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n666_), .A2(new_n350_), .A3(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n660_), .B1(new_n668_), .B2(G36gat), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT106), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n662_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n661_), .A2(new_n671_), .ZN(G1329gat));
  AOI21_X1  g471(.A(G43gat), .B1(new_n630_), .B2(new_n621_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n621_), .A2(G43gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n649_), .B2(new_n674_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT47), .Z(G1330gat));
  NOR3_X1   g475(.A1(new_n646_), .A2(new_n648_), .A3(new_n427_), .ZN(new_n677_));
  INV_X1    g476(.A(G50gat), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n278_), .A2(new_n678_), .ZN(new_n679_));
  OAI22_X1  g478(.A1(new_n677_), .A2(new_n678_), .B1(new_n657_), .B2(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT107), .ZN(G1331gat));
  NAND2_X1  g480(.A1(new_n541_), .A2(new_n461_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n642_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n605_), .A2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G57gat), .B1(new_n684_), .B2(new_n423_), .ZN(new_n685_));
  NOR4_X1   g484(.A1(new_n434_), .A2(new_n460_), .A3(new_n642_), .A4(new_n542_), .ZN(new_n686_));
  INV_X1    g485(.A(G57gat), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n686_), .A2(new_n687_), .A3(new_n391_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n685_), .A2(new_n688_), .ZN(G1332gat));
  OAI21_X1  g488(.A(G64gat), .B1(new_n684_), .B2(new_n349_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT48), .ZN(new_n691_));
  INV_X1    g490(.A(G64gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n686_), .A2(new_n692_), .A3(new_n350_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1333gat));
  NAND3_X1  g493(.A1(new_n686_), .A2(new_n393_), .A3(new_n621_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G71gat), .B1(new_n684_), .B2(new_n403_), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT109), .Z(new_n697_));
  XNOR2_X1  g496(.A(KEYINPUT108), .B(KEYINPUT49), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n697_), .A2(new_n698_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n695_), .B1(new_n699_), .B2(new_n700_), .ZN(G1334gat));
  OAI21_X1  g500(.A(G78gat), .B1(new_n684_), .B2(new_n427_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT50), .ZN(new_n703_));
  INV_X1    g502(.A(G78gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n686_), .A2(new_n704_), .A3(new_n278_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(G1335gat));
  NOR2_X1   g505(.A1(new_n434_), .A2(new_n460_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n642_), .A2(new_n589_), .A3(new_n541_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n710_), .A2(new_n484_), .A3(new_n391_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n642_), .A2(new_n460_), .A3(new_n541_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n641_), .A2(KEYINPUT110), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n641_), .A2(KEYINPUT110), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n713_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n716_), .A2(new_n391_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n711_), .B1(new_n717_), .B2(new_n484_), .ZN(G1336gat));
  NAND3_X1  g517(.A1(new_n710_), .A2(new_n485_), .A3(new_n350_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n716_), .A2(new_n350_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n720_), .B2(new_n485_), .ZN(G1337gat));
  AOI21_X1  g520(.A(new_n395_), .B1(new_n716_), .B2(new_n621_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n621_), .A2(new_n481_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n709_), .A2(new_n723_), .ZN(new_n724_));
  OAI211_X1 g523(.A(KEYINPUT111), .B(KEYINPUT51), .C1(new_n722_), .C2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n726_));
  AOI211_X1 g525(.A(new_n403_), .B(new_n713_), .C1(new_n714_), .C2(new_n715_), .ZN(new_n727_));
  OAI221_X1 g526(.A(new_n726_), .B1(new_n709_), .B2(new_n723_), .C1(new_n727_), .C2(new_n395_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n725_), .A2(new_n728_), .ZN(G1338gat));
  NAND3_X1  g528(.A1(new_n710_), .A2(new_n482_), .A3(new_n278_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n712_), .A2(new_n278_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n632_), .B2(new_n640_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT112), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT52), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n482_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n734_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n735_), .B1(new_n734_), .B2(new_n736_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n730_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT53), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT53), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n741_), .B(new_n730_), .C1(new_n737_), .C2(new_n738_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(G1339gat));
  NAND3_X1  g542(.A1(new_n351_), .A2(new_n391_), .A3(new_n621_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT113), .ZN(new_n745_));
  OR3_X1    g544(.A1(new_n571_), .A2(new_n682_), .A3(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n571_), .B2(new_n682_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n634_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n748_), .B(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n455_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n446_), .B1(new_n450_), .B2(new_n444_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n449_), .A2(new_n752_), .ZN(new_n753_));
  AOI22_X1  g552(.A1(new_n452_), .A2(new_n455_), .B1(new_n751_), .B2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n566_), .A2(new_n754_), .ZN(new_n755_));
  AOI22_X1  g554(.A1(new_n552_), .A2(new_n553_), .B1(new_n490_), .B2(new_n526_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n555_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n549_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT55), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n556_), .A2(new_n759_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n756_), .A2(KEYINPUT55), .A3(new_n548_), .A4(new_n555_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n758_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n563_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT56), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n762_), .A2(KEYINPUT56), .A3(new_n563_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n755_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT117), .ZN(new_n768_));
  OR3_X1    g567(.A1(new_n767_), .A2(new_n768_), .A3(KEYINPUT58), .ZN(new_n769_));
  OAI21_X1  g568(.A(KEYINPUT58), .B1(new_n767_), .B2(new_n768_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n770_), .A3(new_n634_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n460_), .A2(new_n566_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n763_), .A2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n772_), .B1(new_n774_), .B2(new_n764_), .ZN(new_n775_));
  AOI21_X1  g574(.A(KEYINPUT115), .B1(new_n762_), .B2(new_n563_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT56), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n567_), .A2(new_n754_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n780_), .A2(new_n589_), .A3(new_n782_), .ZN(new_n783_));
  AOI22_X1  g582(.A1(new_n775_), .A2(new_n777_), .B1(new_n567_), .B2(new_n754_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n781_), .B1(new_n784_), .B2(new_n604_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n771_), .A2(new_n783_), .A3(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n586_), .ZN(new_n787_));
  AOI211_X1 g586(.A(KEYINPUT59), .B(new_n744_), .C1(new_n750_), .C2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT118), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n786_), .A2(new_n789_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n771_), .A2(new_n783_), .A3(new_n785_), .A4(KEYINPUT118), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n586_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n750_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n744_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n788_), .B1(new_n795_), .B2(KEYINPUT59), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n460_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(G113gat), .ZN(new_n798_));
  OR2_X1    g597(.A1(new_n461_), .A2(G113gat), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n795_), .B2(new_n799_), .ZN(G1340gat));
  INV_X1    g599(.A(G120gat), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT59), .ZN(new_n802_));
  XOR2_X1   g601(.A(new_n748_), .B(new_n749_), .Z(new_n803_));
  INV_X1    g602(.A(new_n787_), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n802_), .B(new_n794_), .C1(new_n803_), .C2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n786_), .A2(new_n789_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(new_n586_), .A3(new_n791_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n744_), .B1(new_n807_), .B2(new_n750_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n805_), .B(new_n571_), .C1(new_n808_), .C2(new_n802_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT119), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n801_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n810_), .B2(new_n809_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n801_), .B1(new_n642_), .B2(KEYINPUT60), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n808_), .B(new_n813_), .C1(KEYINPUT60), .C2(new_n801_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(G1341gat));
  OAI211_X1 g614(.A(new_n805_), .B(new_n541_), .C1(new_n808_), .C2(new_n802_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n816_), .A2(G127gat), .ZN(new_n817_));
  OR2_X1    g616(.A1(new_n586_), .A2(G127gat), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n795_), .A2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(KEYINPUT120), .B1(new_n817_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n816_), .A2(G127gat), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT120), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n821_), .B(new_n822_), .C1(new_n795_), .C2(new_n818_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n820_), .A2(new_n823_), .ZN(G1342gat));
  XNOR2_X1  g623(.A(KEYINPUT121), .B(G134gat), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n519_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n796_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(G134gat), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(new_n795_), .B2(new_n589_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT122), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n827_), .A2(KEYINPUT122), .A3(new_n829_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(G1343gat));
  INV_X1    g633(.A(new_n793_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n637_), .A2(new_n391_), .A3(new_n403_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n460_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n571_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g640(.A(KEYINPUT123), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n837_), .B2(new_n541_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NOR4_X1   g643(.A1(new_n835_), .A2(KEYINPUT123), .A3(new_n586_), .A4(new_n836_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(KEYINPUT61), .B(G155gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n844_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n847_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n843_), .B2(new_n845_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n850_), .ZN(G1346gat));
  INV_X1    g650(.A(new_n837_), .ZN(new_n852_));
  OAI21_X1  g651(.A(G162gat), .B1(new_n852_), .B2(new_n519_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n837_), .A2(new_n222_), .A3(new_n604_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(G1347gat));
  INV_X1    g654(.A(KEYINPUT62), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n404_), .A2(new_n350_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n427_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n859_), .B1(new_n750_), .B2(new_n787_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(new_n461_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT22), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n856_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(G169gat), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n296_), .B1(new_n862_), .B2(new_n856_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n864_), .B2(new_n866_), .ZN(G1348gat));
  AOI21_X1  g666(.A(G176gat), .B1(new_n860_), .B2(new_n571_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n835_), .A2(new_n278_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n642_), .A2(new_n857_), .A3(new_n297_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n868_), .B1(new_n869_), .B2(new_n870_), .ZN(G1349gat));
  NAND3_X1  g670(.A1(new_n869_), .A2(new_n541_), .A3(new_n858_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n586_), .B1(new_n307_), .B2(new_n310_), .ZN(new_n873_));
  AOI22_X1  g672(.A1(new_n872_), .A2(new_n301_), .B1(new_n860_), .B2(new_n873_), .ZN(G1350gat));
  NAND3_X1  g673(.A1(new_n860_), .A2(new_n317_), .A3(new_n604_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n302_), .B1(new_n860_), .B2(new_n634_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n876_), .A2(new_n877_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n875_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(KEYINPUT125), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT125), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n882_), .B(new_n875_), .C1(new_n878_), .C2(new_n879_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n883_), .ZN(G1351gat));
  NAND4_X1  g683(.A1(new_n423_), .A2(new_n278_), .A3(new_n350_), .A4(new_n403_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n835_), .A2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n460_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n571_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g689(.A(new_n586_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n886_), .A2(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(KEYINPUT126), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n892_), .B1(KEYINPUT127), .B2(new_n894_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n894_), .B(KEYINPUT127), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n895_), .B1(new_n892_), .B2(new_n896_), .ZN(G1354gat));
  INV_X1    g696(.A(G218gat), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n886_), .A2(new_n898_), .A3(new_n604_), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n835_), .A2(new_n519_), .A3(new_n885_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(new_n898_), .ZN(G1355gat));
endmodule


