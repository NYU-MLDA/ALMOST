//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 0 0 1 0 1 1 1 1 0 0 1 0 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n650_, new_n651_, new_n652_, new_n654_, new_n655_,
    new_n656_, new_n658_, new_n659_, new_n660_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n784_, new_n785_, new_n786_, new_n787_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n803_, new_n804_, new_n805_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n815_, new_n816_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n835_, new_n837_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_;
  NOR2_X1   g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT23), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204_));
  AOI21_X1  g003(.A(new_n202_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n205_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT22), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n207_), .A2(KEYINPUT80), .ZN(new_n208_));
  OAI21_X1  g007(.A(G169gat), .B1(new_n208_), .B2(G176gat), .ZN(new_n209_));
  INV_X1    g008(.A(G169gat), .ZN(new_n210_));
  INV_X1    g009(.A(G176gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n206_), .B(new_n209_), .C1(new_n208_), .C2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT25), .B(G183gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT79), .ZN(new_n215_));
  INV_X1    g014(.A(G190gat), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n216_), .A2(KEYINPUT26), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n214_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT26), .B(G190gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n219_), .A2(KEYINPUT79), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n204_), .B(KEYINPUT23), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n212_), .A2(KEYINPUT24), .A3(new_n223_), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n222_), .B(new_n224_), .C1(KEYINPUT24), .C2(new_n212_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n213_), .B1(new_n221_), .B2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT81), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G71gat), .B(G99gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(G43gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n227_), .B(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G227gat), .A2(G233gat), .ZN(new_n231_));
  INV_X1    g030(.A(G15gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT30), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT31), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n230_), .B(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT82), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G127gat), .B(G134gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G113gat), .B(G120gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n238_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G197gat), .B(G204gat), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT21), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G211gat), .B(G218gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n243_), .A2(new_n244_), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT86), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT86), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n250_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n249_), .B1(new_n248_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G155gat), .A2(G162gat), .ZN(new_n253_));
  NOR2_X1   g052(.A1(G155gat), .A2(G162gat), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(G141gat), .A2(G148gat), .ZN(new_n256_));
  XOR2_X1   g055(.A(new_n256_), .B(KEYINPUT3), .Z(new_n257_));
  NAND2_X1  g056(.A1(G141gat), .A2(G148gat), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n258_), .B(KEYINPUT2), .Z(new_n259_));
  OAI211_X1 g058(.A(new_n253_), .B(new_n255_), .C1(new_n257_), .C2(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n253_), .A2(KEYINPUT1), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n253_), .B1(new_n254_), .B2(KEYINPUT1), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n261_), .B1(new_n262_), .B2(KEYINPUT83), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n263_), .B1(KEYINPUT83), .B2(new_n262_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n258_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n265_), .A2(new_n256_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n264_), .A2(KEYINPUT84), .A3(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT84), .B1(new_n264_), .B2(new_n266_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n260_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n252_), .B1(new_n270_), .B2(KEYINPUT29), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(G228gat), .ZN(new_n273_));
  INV_X1    g072(.A(G233gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n272_), .A2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n271_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G78gat), .B(G106gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT88), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT88), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n278_), .A2(new_n282_), .A3(new_n279_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n279_), .B(KEYINPUT87), .Z(new_n285_));
  NAND3_X1  g084(.A1(new_n276_), .A2(new_n277_), .A3(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G22gat), .B(G50gat), .ZN(new_n287_));
  OR3_X1    g086(.A1(new_n270_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT28), .B1(new_n270_), .B2(KEYINPUT29), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n287_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n288_), .A2(new_n289_), .A3(new_n287_), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n286_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n284_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n292_), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT85), .B1(new_n295_), .B2(new_n290_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT85), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n291_), .A2(new_n297_), .A3(new_n292_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n285_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n278_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n286_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n299_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n294_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G1gat), .B(G29gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(G85gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT0), .B(G57gat), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n306_), .B(new_n307_), .Z(new_n308_));
  NAND2_X1  g107(.A1(G225gat), .A2(G233gat), .ZN(new_n309_));
  INV_X1    g108(.A(new_n241_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n270_), .A2(new_n310_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n311_), .A2(KEYINPUT4), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT95), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n241_), .B(new_n260_), .C1(new_n268_), .C2(new_n269_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n311_), .A2(KEYINPUT4), .A3(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n312_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n311_), .A2(KEYINPUT95), .A3(KEYINPUT4), .A4(new_n314_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n309_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n311_), .A2(new_n314_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n309_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n308_), .B1(new_n318_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT33), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(G64gat), .B(G92gat), .Z(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT94), .ZN(new_n326_));
  XOR2_X1   g125(.A(G8gat), .B(G36gat), .Z(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT81), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n226_), .B(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n252_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G226gat), .A2(G233gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT19), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT22), .B(G169gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(new_n211_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n206_), .A2(new_n223_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(new_n212_), .A3(new_n223_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n219_), .A2(new_n214_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT90), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n222_), .B1(new_n212_), .B2(new_n342_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT91), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n341_), .B1(new_n347_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n252_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n334_), .A2(KEYINPUT20), .A3(new_n337_), .A4(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT20), .B1(new_n332_), .B2(new_n333_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT92), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n354_), .B1(new_n350_), .B2(new_n252_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n347_), .A2(new_n349_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n340_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n357_), .A2(KEYINPUT92), .A3(new_n333_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n353_), .B1(new_n355_), .B2(new_n358_), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n330_), .B(new_n352_), .C1(new_n359_), .C2(new_n337_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n358_), .A2(new_n355_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT20), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n363_), .B1(new_n227_), .B2(new_n252_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n336_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n330_), .B1(new_n366_), .B2(new_n352_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n361_), .A2(new_n367_), .ZN(new_n368_));
  OAI211_X1 g167(.A(KEYINPUT33), .B(new_n308_), .C1(new_n318_), .C2(new_n321_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n316_), .A2(new_n309_), .A3(new_n317_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n308_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n324_), .A2(new_n368_), .A3(new_n369_), .A4(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n334_), .A2(KEYINPUT20), .A3(new_n351_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(new_n336_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n362_), .A2(new_n337_), .A3(new_n364_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n366_), .A2(new_n352_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n330_), .A2(KEYINPUT32), .ZN(new_n379_));
  MUX2_X1   g178(.A(new_n377_), .B(new_n378_), .S(new_n379_), .Z(new_n380_));
  INV_X1    g179(.A(new_n322_), .ZN(new_n381_));
  NOR3_X1   g180(.A1(new_n318_), .A2(new_n308_), .A3(new_n321_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n380_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n304_), .B1(new_n373_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT27), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n385_), .B1(new_n361_), .B2(new_n367_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n360_), .B(KEYINPUT27), .C1(new_n377_), .C2(new_n330_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  AOI22_X1  g187(.A1(new_n284_), .A2(new_n293_), .B1(new_n299_), .B2(new_n302_), .ZN(new_n389_));
  OR3_X1    g188(.A1(new_n318_), .A2(new_n308_), .A3(new_n321_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n322_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n388_), .A2(new_n389_), .A3(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n242_), .B1(new_n384_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT96), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n238_), .B(new_n310_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n391_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n304_), .A2(new_n388_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n396_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  OAI211_X1 g198(.A(KEYINPUT96), .B(new_n242_), .C1(new_n384_), .C2(new_n392_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n395_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G15gat), .B(G22gat), .ZN(new_n402_));
  INV_X1    g201(.A(G1gat), .ZN(new_n403_));
  INV_X1    g202(.A(G8gat), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT14), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n402_), .B1(new_n405_), .B2(KEYINPUT75), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n405_), .A2(KEYINPUT75), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G1gat), .B(G8gat), .ZN(new_n408_));
  OR3_X1    g207(.A1(new_n406_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n408_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G29gat), .B(G36gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G43gat), .B(G50gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n411_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n409_), .A2(new_n410_), .A3(new_n414_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G229gat), .A2(G233gat), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n418_), .A2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n414_), .B(KEYINPUT15), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n411_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n423_), .A2(new_n417_), .A3(new_n419_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n421_), .A2(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(G113gat), .B(G141gat), .Z(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT78), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G169gat), .B(G197gat), .ZN(new_n428_));
  XOR2_X1   g227(.A(new_n427_), .B(new_n428_), .Z(new_n429_));
  OR2_X1    g228(.A1(new_n425_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n425_), .A2(new_n429_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G230gat), .A2(G233gat), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT8), .ZN(new_n435_));
  XOR2_X1   g234(.A(G85gat), .B(G92gat), .Z(new_n436_));
  NAND2_X1  g235(.A1(G99gat), .A2(G106gat), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT6), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT7), .ZN(new_n440_));
  INV_X1    g239(.A(G99gat), .ZN(new_n441_));
  INV_X1    g240(.A(G106gat), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n435_), .B(new_n436_), .C1(new_n439_), .C2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT67), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT66), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n443_), .A2(new_n448_), .A3(new_n444_), .ZN(new_n449_));
  AND2_X1   g248(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n450_));
  NOR2_X1   g249(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n437_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  OR2_X1    g251(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n453_));
  AND2_X1   g252(.A1(G99gat), .A2(G106gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n453_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n449_), .A2(new_n452_), .A3(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n448_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n447_), .B(new_n436_), .C1(new_n457_), .C2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT8), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n445_), .A2(KEYINPUT66), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n461_), .A2(new_n449_), .A3(new_n452_), .A4(new_n456_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n447_), .B1(new_n462_), .B2(new_n436_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n446_), .B1(new_n460_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n439_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n436_), .A2(KEYINPUT9), .ZN(new_n466_));
  XOR2_X1   g265(.A(KEYINPUT10), .B(G99gat), .Z(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(new_n442_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT64), .B(G92gat), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT9), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(new_n470_), .A3(G85gat), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n465_), .A2(new_n466_), .A3(new_n468_), .A4(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n464_), .A2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G57gat), .B(G64gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT11), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT68), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n474_), .A2(KEYINPUT11), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G71gat), .B(G78gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n476_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT68), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n475_), .B(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n477_), .A2(new_n478_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n479_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n473_), .A2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n464_), .A2(new_n484_), .A3(new_n472_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n486_), .A2(KEYINPUT12), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT12), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n473_), .A2(new_n489_), .A3(new_n485_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n434_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n486_), .A2(KEYINPUT69), .A3(new_n487_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n484_), .B1(new_n464_), .B2(new_n472_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT69), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n433_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n491_), .B1(new_n492_), .B2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G120gat), .B(G148gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT5), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G176gat), .B(G204gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT70), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n496_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n496_), .A2(new_n500_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT13), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT13), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n502_), .A2(new_n506_), .A3(new_n503_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G183gat), .B(G211gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT77), .ZN(new_n510_));
  XOR2_X1   g309(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G127gat), .B(G155gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT17), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G231gat), .A2(G233gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n411_), .B(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(new_n485_), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n515_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(KEYINPUT17), .A3(new_n514_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n473_), .A2(new_n415_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n522_), .B1(new_n422_), .B2(new_n473_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G232gat), .A2(G233gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT34), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n525_), .B(KEYINPUT35), .Z(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(KEYINPUT35), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n527_), .B(KEYINPUT73), .C1(new_n523_), .C2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT73), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n523_), .A2(new_n530_), .A3(new_n526_), .ZN(new_n531_));
  XOR2_X1   g330(.A(G190gat), .B(G218gat), .Z(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT71), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G134gat), .B(G162gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT36), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n536_), .B(KEYINPUT74), .Z(new_n537_));
  AND3_X1   g336(.A1(new_n529_), .A2(new_n531_), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n535_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n542_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n543_));
  OAI21_X1  g342(.A(KEYINPUT37), .B1(new_n538_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n529_), .A2(new_n531_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n541_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT37), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n529_), .A2(new_n531_), .A3(new_n536_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n546_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n521_), .B1(new_n544_), .B2(new_n549_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n401_), .A2(new_n432_), .A3(new_n508_), .A4(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT97), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n552_), .A2(new_n403_), .A3(new_n391_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT38), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n546_), .A2(new_n548_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n401_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n508_), .A2(new_n432_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n558_), .A2(new_n521_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(G1gat), .B1(new_n560_), .B2(new_n397_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n553_), .A2(new_n554_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n555_), .A2(new_n561_), .A3(new_n562_), .ZN(G1324gat));
  INV_X1    g362(.A(new_n552_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n388_), .A2(new_n404_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n557_), .A2(new_n388_), .A3(new_n559_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT39), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n566_), .A2(new_n567_), .A3(G8gat), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n567_), .B1(new_n566_), .B2(G8gat), .ZN(new_n569_));
  OAI22_X1  g368(.A1(new_n564_), .A2(new_n565_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT40), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(G1325gat));
  OAI21_X1  g371(.A(G15gat), .B1(new_n560_), .B2(new_n242_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT98), .B(KEYINPUT41), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n574_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n552_), .A2(new_n232_), .A3(new_n396_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .ZN(G1326gat));
  OR2_X1    g377(.A1(new_n389_), .A2(G22gat), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n557_), .A2(new_n304_), .A3(new_n559_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT42), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n580_), .A2(new_n581_), .A3(G22gat), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n581_), .B1(new_n580_), .B2(G22gat), .ZN(new_n583_));
  OAI22_X1  g382(.A1(new_n564_), .A2(new_n579_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT99), .ZN(G1327gat));
  AND2_X1   g384(.A1(new_n401_), .A2(new_n432_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n556_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(new_n521_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT102), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n589_), .A2(new_n508_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n586_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(G29gat), .B1(new_n592_), .B2(new_n391_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT44), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n544_), .A2(new_n549_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT101), .ZN(new_n596_));
  INV_X1    g395(.A(new_n330_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n337_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n352_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n597_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n372_), .A2(new_n360_), .A3(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n601_), .B1(new_n323_), .B2(new_n322_), .ZN(new_n602_));
  AOI22_X1  g401(.A1(new_n602_), .A2(new_n369_), .B1(new_n391_), .B2(new_n380_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n386_), .A2(new_n387_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(new_n304_), .ZN(new_n605_));
  OAI22_X1  g404(.A1(new_n603_), .A2(new_n304_), .B1(new_n605_), .B2(new_n391_), .ZN(new_n606_));
  AOI21_X1  g405(.A(KEYINPUT96), .B1(new_n606_), .B2(new_n242_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n400_), .A2(new_n399_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n596_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(KEYINPUT100), .B(KEYINPUT43), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n595_), .A2(KEYINPUT43), .ZN(new_n612_));
  AOI22_X1  g411(.A1(new_n609_), .A2(new_n611_), .B1(new_n401_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n521_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n558_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n594_), .B1(new_n613_), .B2(new_n616_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n401_), .A2(new_n612_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n610_), .B1(new_n401_), .B2(new_n596_), .ZN(new_n619_));
  OAI211_X1 g418(.A(KEYINPUT44), .B(new_n615_), .C1(new_n618_), .C2(new_n619_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n617_), .A2(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n391_), .A2(G29gat), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n593_), .B1(new_n621_), .B2(new_n622_), .ZN(G1328gat));
  NAND3_X1  g422(.A1(new_n617_), .A2(new_n388_), .A3(new_n620_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(G36gat), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n604_), .A2(G36gat), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n586_), .A2(new_n590_), .A3(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT45), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n625_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT46), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n625_), .A2(KEYINPUT46), .A3(new_n628_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(G1329gat));
  NAND4_X1  g432(.A1(new_n617_), .A2(G43gat), .A3(new_n396_), .A4(new_n620_), .ZN(new_n634_));
  INV_X1    g433(.A(G43gat), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n635_), .B1(new_n591_), .B2(new_n242_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g437(.A1(new_n621_), .A2(new_n304_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(G50gat), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n389_), .A2(G50gat), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT103), .Z(new_n642_));
  OAI21_X1  g441(.A(new_n640_), .B1(new_n591_), .B2(new_n642_), .ZN(G1331gat));
  NOR2_X1   g442(.A1(new_n508_), .A2(new_n432_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n401_), .A2(new_n614_), .A3(new_n556_), .A4(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(G57gat), .B1(new_n645_), .B2(new_n397_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n401_), .A2(new_n550_), .A3(new_n644_), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n397_), .A2(G57gat), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n646_), .B1(new_n647_), .B2(new_n648_), .ZN(G1332gat));
  OAI21_X1  g448(.A(G64gat), .B1(new_n645_), .B2(new_n604_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT48), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n604_), .A2(G64gat), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n651_), .B1(new_n647_), .B2(new_n652_), .ZN(G1333gat));
  OAI21_X1  g452(.A(G71gat), .B1(new_n645_), .B2(new_n242_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT49), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n242_), .A2(G71gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n655_), .B1(new_n647_), .B2(new_n656_), .ZN(G1334gat));
  OAI21_X1  g456(.A(G78gat), .B1(new_n645_), .B2(new_n389_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT50), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n389_), .A2(G78gat), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n659_), .B1(new_n647_), .B2(new_n660_), .ZN(G1335gat));
  NAND3_X1  g460(.A1(new_n401_), .A2(new_n589_), .A3(new_n644_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT104), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n401_), .A2(KEYINPUT104), .A3(new_n589_), .A4(new_n644_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(G85gat), .B1(new_n666_), .B2(new_n391_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n613_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n644_), .A2(new_n521_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT105), .Z(new_n670_));
  AND2_X1   g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n391_), .A2(G85gat), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT106), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n667_), .B1(new_n671_), .B2(new_n673_), .ZN(G1336gat));
  AOI21_X1  g473(.A(G92gat), .B1(new_n666_), .B2(new_n388_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n388_), .A2(new_n469_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT107), .Z(new_n677_));
  AOI21_X1  g476(.A(new_n675_), .B1(new_n671_), .B2(new_n677_), .ZN(G1337gat));
  NOR2_X1   g477(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n666_), .A2(new_n396_), .A3(new_n467_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n396_), .B(new_n670_), .C1(new_n618_), .C2(new_n619_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(G99gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n679_), .B1(new_n680_), .B2(new_n682_), .ZN(new_n683_));
  AND2_X1   g482(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n683_), .B(new_n684_), .ZN(G1338gat));
  OAI211_X1 g484(.A(new_n304_), .B(new_n670_), .C1(new_n618_), .C2(new_n619_), .ZN(new_n686_));
  XOR2_X1   g485(.A(KEYINPUT110), .B(KEYINPUT52), .Z(new_n687_));
  AND3_X1   g486(.A1(new_n686_), .A2(G106gat), .A3(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n686_), .B2(G106gat), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT109), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n389_), .A2(G106gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n666_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n691_), .ZN(new_n693_));
  AOI211_X1 g492(.A(KEYINPUT109), .B(new_n693_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n694_));
  OAI22_X1  g493(.A1(new_n688_), .A2(new_n689_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT53), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT53), .ZN(new_n697_));
  OAI221_X1 g496(.A(new_n697_), .B1(new_n692_), .B2(new_n694_), .C1(new_n688_), .C2(new_n689_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(G1339gat));
  NAND2_X1  g498(.A1(new_n418_), .A2(new_n419_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n423_), .A2(new_n417_), .A3(new_n420_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n700_), .A2(new_n701_), .A3(new_n429_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n430_), .A2(new_n702_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n703_), .A2(KEYINPUT113), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(KEYINPUT113), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n487_), .A2(KEYINPUT12), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n709_), .A2(new_n493_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n490_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n433_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT55), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n491_), .A2(KEYINPUT55), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n488_), .A2(new_n434_), .A3(new_n490_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(KEYINPUT111), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT111), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n488_), .A2(new_n718_), .A3(new_n434_), .A4(new_n490_), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n714_), .A2(new_n715_), .A3(new_n717_), .A4(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n501_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n720_), .A2(KEYINPUT56), .A3(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT112), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(KEYINPUT56), .B1(new_n720_), .B2(new_n721_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n720_), .A2(new_n721_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT56), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n727_), .A2(KEYINPUT112), .A3(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n503_), .A2(new_n432_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n708_), .B1(new_n726_), .B2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n556_), .A2(KEYINPUT57), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n733_), .A2(KEYINPUT115), .A3(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT57), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n727_), .A2(new_n728_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n738_), .A2(new_n723_), .A3(new_n722_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n730_), .B1(new_n725_), .B2(KEYINPUT112), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n707_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n741_), .B2(new_n587_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT115), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n743_), .B1(new_n741_), .B2(new_n734_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n736_), .A2(new_n742_), .A3(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT114), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n738_), .A2(new_n746_), .A3(new_n722_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n720_), .A2(KEYINPUT114), .A3(KEYINPUT56), .A4(new_n721_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n706_), .B1(new_n496_), .B2(new_n500_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n747_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT58), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n595_), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n747_), .A2(KEYINPUT58), .A3(new_n748_), .A4(new_n749_), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n752_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n521_), .B1(new_n745_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n432_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n550_), .A2(new_n508_), .A3(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT54), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n758_), .B(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n756_), .A2(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n396_), .A2(new_n391_), .A3(new_n398_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n762_), .A2(KEYINPUT116), .A3(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT116), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n752_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n767_), .A2(new_n736_), .A3(new_n742_), .A4(new_n744_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n760_), .B1(new_n768_), .B2(new_n521_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n766_), .B1(new_n769_), .B2(new_n763_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n765_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(G113gat), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n772_), .A3(new_n432_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT117), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n762_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n762_), .A2(new_n764_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT59), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n775_), .A2(new_n776_), .A3(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n769_), .B2(KEYINPUT117), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n769_), .A2(new_n763_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n757_), .B1(new_n778_), .B2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n773_), .B1(new_n782_), .B2(new_n772_), .ZN(G1340gat));
  INV_X1    g582(.A(G120gat), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n784_), .B1(new_n508_), .B2(KEYINPUT60), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n771_), .B(new_n785_), .C1(KEYINPUT60), .C2(new_n784_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n508_), .B1(new_n778_), .B2(new_n781_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n786_), .B1(new_n784_), .B2(new_n787_), .ZN(G1341gat));
  INV_X1    g587(.A(KEYINPUT118), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n765_), .A2(new_n614_), .A3(new_n770_), .ZN(new_n790_));
  INV_X1    g589(.A(G127gat), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n521_), .A2(new_n791_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n794_), .B1(new_n778_), .B2(new_n781_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n789_), .B1(new_n792_), .B2(new_n795_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n779_), .A2(new_n780_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n779_), .A2(new_n780_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n793_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n790_), .A2(new_n791_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(KEYINPUT118), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n796_), .A2(new_n801_), .ZN(G1342gat));
  INV_X1    g601(.A(G134gat), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n771_), .A2(new_n803_), .A3(new_n587_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n595_), .B1(new_n778_), .B2(new_n781_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(new_n803_), .ZN(G1343gat));
  INV_X1    g605(.A(KEYINPUT119), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n396_), .A2(new_n605_), .A3(new_n397_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n762_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n808_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT119), .B1(new_n769_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n432_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g613(.A(new_n508_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n812_), .A2(new_n815_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g616(.A1(new_n812_), .A2(new_n614_), .ZN(new_n818_));
  XOR2_X1   g617(.A(KEYINPUT61), .B(G155gat), .Z(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(KEYINPUT121), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(KEYINPUT120), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n818_), .B(new_n821_), .ZN(G1346gat));
  AND3_X1   g621(.A1(new_n812_), .A2(G162gat), .A3(new_n596_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n556_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n824_));
  OR3_X1    g623(.A1(new_n824_), .A2(KEYINPUT122), .A3(G162gat), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT122), .B1(new_n824_), .B2(G162gat), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n823_), .B1(new_n825_), .B2(new_n826_), .ZN(G1347gat));
  NAND4_X1  g626(.A1(new_n396_), .A2(new_n389_), .A3(new_n397_), .A4(new_n388_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n769_), .A2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n210_), .B1(new_n829_), .B2(new_n432_), .ZN(new_n830_));
  OR2_X1    g629(.A1(new_n830_), .A2(KEYINPUT62), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n829_), .A2(new_n338_), .A3(new_n432_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(KEYINPUT62), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n831_), .A2(new_n832_), .A3(new_n833_), .ZN(G1348gat));
  NAND2_X1  g633(.A1(new_n829_), .A2(new_n815_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g635(.A1(new_n829_), .A2(new_n614_), .ZN(new_n837_));
  MUX2_X1   g636(.A(new_n214_), .B(G183gat), .S(new_n837_), .Z(G1350gat));
  NAND2_X1  g637(.A1(new_n587_), .A2(new_n219_), .ZN(new_n839_));
  XOR2_X1   g638(.A(new_n839_), .B(KEYINPUT123), .Z(new_n840_));
  NAND2_X1  g639(.A1(new_n829_), .A2(new_n840_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n769_), .A2(new_n595_), .A3(new_n828_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n842_), .B2(new_n216_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(KEYINPUT124), .ZN(G1351gat));
  NOR4_X1   g643(.A1(new_n396_), .A2(new_n389_), .A3(new_n391_), .A4(new_n604_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n762_), .A2(new_n845_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n846_), .A2(new_n757_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(KEYINPUT125), .B(G197gat), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n847_), .B(new_n848_), .ZN(G1352gat));
  INV_X1    g648(.A(new_n846_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n815_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g651(.A(KEYINPUT127), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n846_), .A2(new_n521_), .ZN(new_n854_));
  OR2_X1    g653(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n853_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  OR3_X1    g655(.A1(new_n854_), .A2(new_n853_), .A3(new_n855_), .ZN(new_n857_));
  XOR2_X1   g656(.A(KEYINPUT63), .B(G211gat), .Z(new_n858_));
  NAND2_X1  g657(.A1(new_n854_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(KEYINPUT126), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT126), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n854_), .A2(new_n861_), .A3(new_n858_), .ZN(new_n862_));
  AOI22_X1  g661(.A1(new_n856_), .A2(new_n857_), .B1(new_n860_), .B2(new_n862_), .ZN(G1354gat));
  OR3_X1    g662(.A1(new_n846_), .A2(G218gat), .A3(new_n556_), .ZN(new_n864_));
  OAI21_X1  g663(.A(G218gat), .B1(new_n846_), .B2(new_n595_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(G1355gat));
endmodule


