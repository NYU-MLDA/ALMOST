//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 0 1 0 0 0 0 1 1 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n782_, new_n783_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n954_,
    new_n955_, new_n957_, new_n958_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n972_, new_n973_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT74), .ZN(new_n203_));
  XOR2_X1   g002(.A(G134gat), .B(G162gat), .Z(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT36), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT36), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G232gat), .A2(G233gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT35), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT15), .ZN(new_n213_));
  INV_X1    g012(.A(G36gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(G29gat), .ZN(new_n215_));
  INV_X1    g014(.A(G29gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(G36gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n217_), .A3(KEYINPUT73), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT73), .B1(new_n215_), .B2(new_n217_), .ZN(new_n220_));
  XOR2_X1   g019(.A(G43gat), .B(G50gat), .Z(new_n221_));
  NOR3_X1   g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G43gat), .B(G50gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n215_), .A2(new_n217_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT73), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n223_), .B1(new_n226_), .B2(new_n218_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n213_), .B1(new_n222_), .B2(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n221_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n226_), .A2(new_n218_), .A3(new_n223_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(new_n230_), .A3(KEYINPUT15), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n228_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G99gat), .A2(G106gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT6), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT6), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(G99gat), .A3(G106gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  OR2_X1    g036(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n238_));
  INV_X1    g037(.A(G106gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(G85gat), .ZN(new_n242_));
  INV_X1    g041(.A(G92gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G85gat), .A2(G92gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(KEYINPUT9), .A3(new_n245_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n245_), .A2(KEYINPUT9), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n237_), .A2(new_n241_), .A3(new_n246_), .A4(new_n247_), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n248_), .A2(KEYINPUT69), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(KEYINPUT69), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT64), .ZN(new_n252_));
  AND2_X1   g051(.A1(G85gat), .A2(G92gat), .ZN(new_n253_));
  NOR2_X1   g052(.A1(G85gat), .A2(G92gat), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n252_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n244_), .A2(KEYINPUT64), .A3(new_n245_), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT8), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT7), .ZN(new_n259_));
  INV_X1    g058(.A(G99gat), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(new_n260_), .A3(new_n239_), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n234_), .A2(new_n236_), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n257_), .B(new_n258_), .C1(new_n263_), .C2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n255_), .A2(new_n256_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT65), .ZN(new_n267_));
  AOI22_X1  g066(.A1(new_n263_), .A2(new_n267_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n261_), .A2(KEYINPUT65), .A3(new_n262_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n266_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n265_), .B1(new_n270_), .B2(new_n258_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n232_), .B1(new_n251_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n229_), .A2(new_n230_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n262_), .ZN(new_n274_));
  NOR3_X1   g073(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n267_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n276_), .A2(new_n269_), .A3(new_n237_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n258_), .B1(new_n277_), .B2(new_n257_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n264_), .A2(new_n263_), .ZN(new_n279_));
  NOR3_X1   g078(.A1(new_n279_), .A2(KEYINPUT8), .A3(new_n266_), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n273_), .B(new_n248_), .C1(new_n278_), .C2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n210_), .A2(new_n211_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n212_), .B1(new_n272_), .B2(new_n283_), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n228_), .A2(new_n231_), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n250_), .B(new_n249_), .C1(new_n278_), .C2(new_n280_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n212_), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n287_), .A2(new_n288_), .A3(new_n282_), .A4(new_n281_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n207_), .B1(new_n284_), .B2(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n206_), .B1(new_n290_), .B2(new_n205_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n284_), .A2(new_n289_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT75), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n291_), .A2(new_n294_), .ZN(new_n295_));
  OAI211_X1 g094(.A(new_n293_), .B(new_n206_), .C1(new_n290_), .C2(new_n205_), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n295_), .A2(KEYINPUT37), .A3(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT37), .B1(new_n295_), .B2(new_n296_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G127gat), .B(G155gat), .Z(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT16), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G183gat), .B(G211gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT17), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT78), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT66), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n306_), .A2(G71gat), .ZN(new_n307_));
  INV_X1    g106(.A(G71gat), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n308_), .A2(KEYINPUT66), .ZN(new_n309_));
  OAI21_X1  g108(.A(G78gat), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(KEYINPUT66), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n306_), .A2(G71gat), .ZN(new_n312_));
  INV_X1    g111(.A(G78gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n311_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(G64gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(G57gat), .ZN(new_n316_));
  INV_X1    g115(.A(G57gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(G64gat), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n316_), .A2(new_n318_), .A3(KEYINPUT11), .ZN(new_n319_));
  AOI21_X1  g118(.A(KEYINPUT11), .B1(new_n316_), .B2(new_n318_), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n310_), .B(new_n314_), .C1(new_n319_), .C2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n316_), .A2(new_n318_), .A3(KEYINPUT11), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n311_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n313_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n322_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n321_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT67), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT67), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n321_), .A2(new_n328_), .A3(new_n325_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT77), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G1gat), .B(G8gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT76), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G15gat), .B(G22gat), .ZN(new_n334_));
  INV_X1    g133(.A(G1gat), .ZN(new_n335_));
  INV_X1    g134(.A(G8gat), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT14), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n334_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n333_), .A2(new_n338_), .ZN(new_n339_));
  OR2_X1    g138(.A1(new_n332_), .A2(KEYINPUT76), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n332_), .A2(KEYINPUT76), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n340_), .A2(new_n337_), .A3(new_n334_), .A4(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n339_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G231gat), .A2(G233gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n331_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n331_), .A2(new_n345_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n305_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT17), .ZN(new_n349_));
  AND2_X1   g148(.A1(new_n345_), .A2(new_n326_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n345_), .A2(new_n326_), .ZN(new_n351_));
  OR4_X1    g150(.A1(new_n349_), .A2(new_n350_), .A3(new_n351_), .A4(new_n303_), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n348_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n299_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT79), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G211gat), .B(G218gat), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(G204gat), .ZN(new_n358_));
  OR3_X1    g157(.A1(new_n358_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n359_));
  INV_X1    g158(.A(G197gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(G204gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT88), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n358_), .A2(G197gat), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n359_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT89), .B(KEYINPUT21), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n357_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT21), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n368_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT87), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n356_), .A2(new_n368_), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n367_), .A2(new_n370_), .B1(new_n364_), .B2(new_n371_), .ZN(new_n372_));
  OR2_X1    g171(.A1(G155gat), .A2(G162gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G155gat), .A2(G162gat), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n373_), .B1(KEYINPUT1), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT86), .ZN(new_n376_));
  AND3_X1   g175(.A1(new_n374_), .A2(new_n376_), .A3(KEYINPUT1), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n376_), .B1(new_n374_), .B2(KEYINPUT1), .ZN(new_n378_));
  NOR3_X1   g177(.A1(new_n375_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G141gat), .A2(G148gat), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(G141gat), .A2(G148gat), .ZN(new_n382_));
  OR3_X1    g181(.A1(new_n379_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(KEYINPUT3), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n380_), .B(KEYINPUT2), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n383_), .A2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n372_), .B1(new_n388_), .B2(KEYINPUT29), .ZN(new_n389_));
  INV_X1    g188(.A(G228gat), .ZN(new_n390_));
  INV_X1    g189(.A(G233gat), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n389_), .B(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G78gat), .B(G106gat), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n396_), .A2(KEYINPUT90), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n394_), .A2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n389_), .B(new_n392_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n397_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n396_), .A2(KEYINPUT90), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n398_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT28), .B1(new_n388_), .B2(KEYINPUT29), .ZN(new_n404_));
  INV_X1    g203(.A(new_n387_), .ZN(new_n405_));
  NOR3_X1   g204(.A1(new_n379_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT28), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT29), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n404_), .A2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G22gat), .B(G50gat), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n404_), .A2(new_n410_), .A3(new_n412_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n396_), .A2(KEYINPUT91), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n416_), .B1(new_n399_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n394_), .A2(new_n417_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n403_), .A2(new_n416_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G127gat), .B(G134gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT85), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G113gat), .B(G120gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  OR2_X1    g225(.A1(new_n422_), .A2(KEYINPUT85), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n422_), .A2(KEYINPUT85), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n427_), .A2(new_n428_), .A3(new_n424_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n426_), .A2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n430_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n383_), .A2(new_n429_), .A3(new_n426_), .A4(new_n387_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(new_n432_), .A3(KEYINPUT4), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G225gat), .A2(G233gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT4), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n388_), .A2(new_n436_), .A3(new_n430_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n433_), .A2(new_n435_), .A3(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n431_), .A2(new_n432_), .A3(new_n434_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G1gat), .B(G29gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(KEYINPUT95), .B(G85gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT0), .B(G57gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n440_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n438_), .A2(new_n439_), .A3(new_n445_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n421_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT27), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT20), .ZN(new_n452_));
  INV_X1    g251(.A(G169gat), .ZN(new_n453_));
  INV_X1    g252(.A(G176gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n455_), .A2(KEYINPUT24), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT26), .B(G190gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT25), .B(G183gat), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n456_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G183gat), .A2(G190gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT23), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G169gat), .A2(G176gat), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n455_), .A2(KEYINPUT24), .A3(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n459_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT22), .B(G169gat), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT81), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n453_), .A2(KEYINPUT22), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n454_), .B1(new_n469_), .B2(KEYINPUT81), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n462_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT82), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n461_), .B1(G183gat), .B2(G190gat), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n465_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n452_), .B1(new_n474_), .B2(new_n372_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n458_), .B(KEYINPUT92), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(new_n457_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n461_), .A2(new_n463_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n478_), .A2(new_n456_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n462_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n480_), .B1(new_n466_), .B2(new_n454_), .ZN(new_n481_));
  AOI22_X1  g280(.A1(new_n477_), .A2(new_n479_), .B1(new_n473_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT93), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n367_), .A2(new_n370_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n364_), .A2(new_n371_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n483_), .A2(new_n484_), .A3(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT93), .B1(new_n372_), .B2(new_n482_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n475_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G226gat), .A2(G233gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT19), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n493_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n452_), .B1(new_n372_), .B2(new_n482_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n495_), .B(new_n496_), .C1(new_n474_), .C2(new_n372_), .ZN(new_n497_));
  XOR2_X1   g296(.A(G8gat), .B(G36gat), .Z(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G64gat), .B(G92gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n494_), .A2(new_n497_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n502_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n495_), .B1(new_n475_), .B2(new_n490_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n497_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n504_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n503_), .A2(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n505_), .A2(new_n506_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n451_), .B1(new_n509_), .B2(new_n502_), .ZN(new_n510_));
  OAI22_X1  g309(.A1(KEYINPUT98), .A2(new_n496_), .B1(new_n474_), .B2(new_n372_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n496_), .A2(KEYINPUT98), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n493_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n475_), .A2(new_n490_), .A3(new_n495_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n504_), .ZN(new_n517_));
  AOI22_X1  g316(.A1(new_n451_), .A2(new_n508_), .B1(new_n510_), .B2(new_n517_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n438_), .A2(KEYINPUT33), .A3(new_n439_), .A4(new_n445_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n433_), .A2(new_n434_), .A3(new_n437_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n431_), .A2(new_n432_), .A3(new_n435_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n446_), .A3(new_n521_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n519_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n503_), .A2(new_n523_), .A3(new_n507_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT96), .B(KEYINPUT33), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n448_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT97), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT97), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n448_), .A2(new_n528_), .A3(new_n525_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n502_), .A2(KEYINPUT32), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n494_), .A2(new_n497_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n449_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n531_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n534_));
  OAI22_X1  g333(.A1(new_n524_), .A2(new_n530_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  AOI22_X1  g334(.A1(new_n450_), .A2(new_n518_), .B1(new_n535_), .B2(new_n421_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n430_), .B(KEYINPUT31), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G227gat), .A2(G233gat), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n537_), .B(new_n538_), .Z(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT83), .B(G43gat), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n474_), .A2(KEYINPUT30), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n474_), .A2(KEYINPUT30), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n542_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n474_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT30), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(new_n543_), .A3(new_n541_), .ZN(new_n550_));
  XOR2_X1   g349(.A(G71gat), .B(G99gat), .Z(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT84), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(G15gat), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n546_), .A2(new_n550_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n554_), .B1(new_n546_), .B2(new_n550_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n540_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n546_), .A2(new_n550_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(new_n553_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n560_), .A2(new_n539_), .A3(new_n555_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n558_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n508_), .A2(new_n451_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n510_), .A2(new_n517_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n421_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n449_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n558_), .A2(new_n567_), .A3(new_n561_), .ZN(new_n568_));
  OAI22_X1  g367(.A1(new_n536_), .A2(new_n563_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n248_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n277_), .A2(new_n257_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT8), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n570_), .B1(new_n572_), .B2(new_n265_), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n321_), .A2(new_n328_), .A3(new_n325_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n328_), .B1(new_n321_), .B2(new_n325_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n248_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n330_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n577_), .A2(KEYINPUT68), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(G230gat), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n581_), .A2(new_n391_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n580_), .B(new_n582_), .C1(KEYINPUT68), .C2(new_n577_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT12), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n584_), .B1(new_n321_), .B2(new_n325_), .ZN(new_n585_));
  AOI22_X1  g384(.A1(new_n579_), .A2(new_n584_), .B1(new_n286_), .B2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n582_), .B1(new_n573_), .B2(new_n576_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n583_), .A2(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(G120gat), .B(G148gat), .Z(new_n590_));
  XNOR2_X1  g389(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G176gat), .B(G204gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n589_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n583_), .A2(new_n588_), .A3(new_n594_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT13), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT13), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n596_), .A2(new_n600_), .A3(new_n597_), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n599_), .A2(KEYINPUT71), .A3(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(KEYINPUT71), .B1(new_n599_), .B2(new_n601_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n343_), .A2(new_n273_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n339_), .A2(new_n230_), .A3(new_n342_), .A4(new_n229_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT80), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G229gat), .A2(G233gat), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n605_), .A2(KEYINPUT80), .A3(new_n606_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n609_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n232_), .A2(new_n343_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n614_), .A2(new_n610_), .A3(new_n605_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G113gat), .B(G141gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G169gat), .B(G197gat), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n617_), .B(new_n618_), .Z(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n616_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n613_), .A2(new_n615_), .A3(new_n619_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n604_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n355_), .A2(new_n569_), .A3(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n626_), .A2(new_n335_), .A3(new_n449_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n628_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n604_), .A2(new_n623_), .A3(new_n353_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT100), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n566_), .A2(new_n568_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n535_), .A2(new_n421_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n402_), .B1(new_n394_), .B2(new_n397_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n399_), .A2(new_n400_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n416_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n419_), .A2(new_n420_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n639_), .A2(new_n564_), .A3(new_n565_), .A4(new_n567_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n634_), .A2(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n633_), .B1(new_n641_), .B2(new_n562_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n295_), .A2(new_n296_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n632_), .B1(new_n642_), .B2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n569_), .A2(KEYINPUT100), .A3(new_n643_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n631_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n647_), .A2(new_n449_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n629_), .B(new_n630_), .C1(new_n335_), .C2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT101), .ZN(G1324gat));
  INV_X1    g449(.A(new_n518_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n626_), .A2(new_n336_), .A3(new_n651_), .ZN(new_n652_));
  AOI211_X1 g451(.A(KEYINPUT102), .B(new_n336_), .C1(new_n647_), .C2(new_n651_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n654_));
  INV_X1    g453(.A(new_n631_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n642_), .A2(new_n632_), .A3(new_n644_), .ZN(new_n656_));
  AOI21_X1  g455(.A(KEYINPUT100), .B1(new_n569_), .B2(new_n643_), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n651_), .B(new_n655_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n654_), .B1(new_n658_), .B2(G8gat), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n653_), .A2(new_n659_), .A3(KEYINPUT39), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT39), .ZN(new_n661_));
  AOI211_X1 g460(.A(new_n518_), .B(new_n631_), .C1(new_n645_), .C2(new_n646_), .ZN(new_n662_));
  OAI21_X1  g461(.A(KEYINPUT102), .B1(new_n662_), .B2(new_n336_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n658_), .A2(new_n654_), .A3(G8gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n661_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n652_), .B1(new_n660_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT40), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  OAI211_X1 g467(.A(KEYINPUT40), .B(new_n652_), .C1(new_n660_), .C2(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1325gat));
  INV_X1    g469(.A(G15gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n626_), .A2(new_n671_), .A3(new_n563_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n647_), .A2(new_n563_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n673_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(KEYINPUT41), .B1(new_n673_), .B2(G15gat), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n672_), .B1(new_n674_), .B2(new_n675_), .ZN(G1326gat));
  INV_X1    g475(.A(G22gat), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n626_), .A2(new_n677_), .A3(new_n639_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n647_), .A2(new_n639_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(G22gat), .ZN(new_n680_));
  XNOR2_X1  g479(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n680_), .A2(new_n681_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n678_), .B1(new_n682_), .B2(new_n683_), .ZN(G1327gat));
  NOR2_X1   g483(.A1(new_n353_), .A2(new_n643_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n625_), .A2(new_n569_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(G29gat), .B1(new_n687_), .B2(new_n449_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT37), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n643_), .A2(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n295_), .A2(KEYINPUT37), .A3(new_n296_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT43), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n569_), .A2(new_n692_), .A3(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n642_), .A2(new_n299_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n695_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n624_), .A2(new_n353_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n698_), .A2(new_n701_), .A3(new_n699_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n567_), .A2(new_n216_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n688_), .B1(new_n705_), .B2(new_n706_), .ZN(G1328gat));
  NAND2_X1  g506(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT46), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n214_), .B1(new_n705_), .B2(new_n651_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n651_), .A2(new_n214_), .ZN(new_n714_));
  OR3_X1    g513(.A1(new_n686_), .A2(new_n713_), .A3(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n713_), .B1(new_n686_), .B2(new_n714_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n708_), .B(new_n711_), .C1(new_n712_), .C2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n704_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n701_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n651_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(G36gat), .ZN(new_n722_));
  INV_X1    g521(.A(new_n717_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n722_), .A2(new_n709_), .A3(new_n710_), .A4(new_n723_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n718_), .A2(new_n724_), .ZN(G1329gat));
  NOR3_X1   g524(.A1(new_n686_), .A2(G43gat), .A3(new_n562_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n705_), .A2(new_n563_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n727_), .B2(G43gat), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  AOI211_X1 g529(.A(KEYINPUT47), .B(new_n726_), .C1(new_n727_), .C2(G43gat), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1330gat));
  AOI21_X1  g531(.A(new_n421_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n733_));
  INV_X1    g532(.A(G50gat), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n639_), .A2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT108), .ZN(new_n736_));
  OAI22_X1  g535(.A1(new_n733_), .A2(new_n734_), .B1(new_n686_), .B2(new_n736_), .ZN(G1331gat));
  INV_X1    g536(.A(new_n604_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n355_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT109), .ZN(new_n740_));
  OR2_X1    g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n642_), .A2(new_n623_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(new_n740_), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n741_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(G57gat), .B1(new_n744_), .B2(new_n449_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n623_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n738_), .A2(new_n746_), .A3(new_n353_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n317_), .B1(new_n449_), .B2(KEYINPUT110), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(KEYINPUT110), .B2(new_n317_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n745_), .B1(new_n748_), .B2(new_n750_), .ZN(G1332gat));
  NAND3_X1  g550(.A1(new_n744_), .A2(new_n315_), .A3(new_n651_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n748_), .A2(new_n651_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(G64gat), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n754_), .A2(KEYINPUT48), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n754_), .A2(KEYINPUT48), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n752_), .B1(new_n755_), .B2(new_n756_), .ZN(G1333gat));
  NAND3_X1  g556(.A1(new_n744_), .A2(new_n308_), .A3(new_n563_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n748_), .A2(new_n563_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(G71gat), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n760_), .A2(KEYINPUT49), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n760_), .A2(KEYINPUT49), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n758_), .B1(new_n761_), .B2(new_n762_), .ZN(G1334gat));
  NAND2_X1  g562(.A1(new_n639_), .A2(new_n313_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT111), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n744_), .A2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n748_), .A2(new_n639_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(G78gat), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n768_), .A2(KEYINPUT50), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(KEYINPUT50), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n766_), .B1(new_n769_), .B2(new_n770_), .ZN(G1335gat));
  NOR3_X1   g570(.A1(new_n604_), .A2(new_n643_), .A3(new_n353_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n742_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(G85gat), .B1(new_n774_), .B2(new_n449_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n604_), .A2(new_n623_), .A3(new_n353_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n698_), .A2(new_n776_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT112), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT113), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n567_), .A2(new_n242_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n775_), .B1(new_n779_), .B2(new_n780_), .ZN(G1336gat));
  AOI21_X1  g580(.A(G92gat), .B1(new_n774_), .B2(new_n651_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n518_), .A2(new_n243_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n779_), .B2(new_n783_), .ZN(G1337gat));
  INV_X1    g583(.A(KEYINPUT114), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT112), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n777_), .B(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n260_), .B1(new_n787_), .B2(new_n563_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n238_), .A2(new_n240_), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n773_), .A2(new_n562_), .A3(new_n789_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n785_), .B(KEYINPUT51), .C1(new_n788_), .C2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(G99gat), .B1(new_n778_), .B2(new_n562_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n785_), .A2(KEYINPUT51), .ZN(new_n793_));
  INV_X1    g592(.A(new_n790_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n792_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n791_), .A2(new_n795_), .ZN(G1338gat));
  NAND3_X1  g595(.A1(new_n774_), .A2(new_n239_), .A3(new_n639_), .ZN(new_n797_));
  OAI21_X1  g596(.A(G106gat), .B1(new_n777_), .B2(new_n421_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n798_), .A2(KEYINPUT52), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n798_), .A2(KEYINPUT52), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n797_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT53), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n803_), .B(new_n797_), .C1(new_n799_), .C2(new_n800_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(G1339gat));
  INV_X1    g604(.A(new_n353_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n623_), .A2(new_n597_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n584_), .B1(new_n573_), .B2(new_n576_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n286_), .A2(new_n585_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(new_n809_), .A3(new_n577_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n582_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n813_));
  AND4_X1   g612(.A1(new_n812_), .A2(new_n808_), .A3(new_n587_), .A4(new_n809_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n811_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT56), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n594_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  AOI22_X1  g617(.A1(new_n271_), .A2(new_n248_), .B1(new_n327_), .B2(new_n329_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n809_), .B1(new_n819_), .B2(KEYINPUT12), .ZN(new_n820_));
  OAI22_X1  g619(.A1(new_n330_), .A2(new_n578_), .B1(new_n581_), .B2(new_n391_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT55), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n808_), .A2(new_n587_), .A3(new_n812_), .A4(new_n809_), .ZN(new_n823_));
  AOI22_X1  g622(.A1(new_n822_), .A2(new_n823_), .B1(new_n582_), .B2(new_n810_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n816_), .B1(new_n824_), .B2(new_n594_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n807_), .B1(new_n818_), .B2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n609_), .A2(new_n610_), .A3(new_n612_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n610_), .B1(new_n343_), .B2(new_n273_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n619_), .B1(new_n614_), .B2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n622_), .A2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n831_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n832_));
  OAI211_X1 g631(.A(KEYINPUT57), .B(new_n643_), .C1(new_n826_), .C2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT57), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n825_), .A2(new_n818_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n807_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n832_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n836_), .B1(new_n839_), .B2(new_n644_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n835_), .B(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n842_));
  INV_X1    g641(.A(new_n817_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n824_), .B2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n815_), .A2(KEYINPUT117), .A3(new_n817_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n825_), .A2(new_n844_), .A3(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n597_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n847_), .A2(new_n831_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT118), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n852_), .A3(new_n692_), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT58), .B1(new_n846_), .B2(new_n848_), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT118), .B1(new_n854_), .B2(new_n299_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n849_), .A2(new_n850_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n853_), .A2(new_n855_), .A3(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n806_), .B1(new_n841_), .B2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n623_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n299_), .A2(new_n353_), .A3(new_n861_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n862_), .B(new_n864_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n860_), .A2(new_n865_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n566_), .A2(new_n562_), .A3(new_n567_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n866_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(G113gat), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n869_), .A2(new_n870_), .A3(new_n623_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n862_), .B(new_n863_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n840_), .A2(new_n833_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n858_), .A2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n872_), .B1(new_n875_), .B2(new_n806_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n876_), .A2(KEYINPUT59), .A3(new_n868_), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n877_), .A2(KEYINPUT119), .ZN(new_n878_));
  OAI21_X1  g677(.A(KEYINPUT59), .B1(new_n866_), .B2(new_n868_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(KEYINPUT119), .ZN(new_n880_));
  AND4_X1   g679(.A1(new_n623_), .A2(new_n878_), .A3(new_n879_), .A4(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n871_), .B1(new_n881_), .B2(new_n870_), .ZN(G1340gat));
  INV_X1    g681(.A(G120gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n604_), .B2(KEYINPUT60), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(KEYINPUT60), .B2(new_n883_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n866_), .A2(new_n868_), .A3(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n886_), .B(new_n887_), .ZN(new_n888_));
  AND4_X1   g687(.A1(new_n738_), .A2(new_n878_), .A3(new_n879_), .A4(new_n880_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(new_n883_), .ZN(G1341gat));
  INV_X1    g689(.A(G127gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n869_), .A2(new_n891_), .A3(new_n353_), .ZN(new_n892_));
  AND4_X1   g691(.A1(new_n353_), .A2(new_n878_), .A3(new_n879_), .A4(new_n880_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n891_), .ZN(G1342gat));
  INV_X1    g693(.A(G134gat), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n869_), .A2(new_n895_), .A3(new_n644_), .ZN(new_n896_));
  AND4_X1   g695(.A1(new_n692_), .A2(new_n878_), .A3(new_n879_), .A4(new_n880_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n897_), .B2(new_n895_), .ZN(G1343gat));
  NOR2_X1   g697(.A1(new_n866_), .A2(new_n563_), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n651_), .A2(new_n567_), .A3(new_n421_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n899_), .A2(new_n623_), .A3(new_n900_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g701(.A1(new_n899_), .A2(new_n738_), .A3(new_n900_), .ZN(new_n903_));
  XOR2_X1   g702(.A(KEYINPUT121), .B(G148gat), .Z(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1345gat));
  NAND3_X1  g704(.A1(new_n899_), .A2(new_n353_), .A3(new_n900_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT61), .B(G155gat), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n906_), .B(new_n907_), .ZN(G1346gat));
  INV_X1    g707(.A(G162gat), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n899_), .A2(new_n909_), .A3(new_n644_), .A4(new_n900_), .ZN(new_n910_));
  AND3_X1   g709(.A1(new_n899_), .A2(new_n692_), .A3(new_n900_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n911_), .B2(new_n909_), .ZN(G1347gat));
  NAND4_X1  g711(.A1(new_n651_), .A2(new_n563_), .A3(new_n567_), .A4(new_n421_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(new_n746_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n353_), .B1(new_n858_), .B2(new_n874_), .ZN(new_n915_));
  OAI211_X1 g714(.A(KEYINPUT122), .B(new_n914_), .C1(new_n915_), .C2(new_n872_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(G169gat), .ZN(new_n917_));
  AOI22_X1  g716(.A1(new_n849_), .A2(new_n850_), .B1(new_n691_), .B2(new_n690_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n856_), .B1(new_n918_), .B2(new_n852_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n873_), .B1(new_n919_), .B2(new_n855_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n865_), .B1(new_n920_), .B2(new_n353_), .ZN(new_n921_));
  AOI21_X1  g720(.A(KEYINPUT122), .B1(new_n921_), .B2(new_n914_), .ZN(new_n922_));
  OAI21_X1  g721(.A(KEYINPUT123), .B1(new_n917_), .B2(new_n922_), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT122), .ZN(new_n924_));
  INV_X1    g723(.A(new_n914_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n876_), .B2(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n927_));
  NAND4_X1  g726(.A1(new_n926_), .A2(new_n927_), .A3(G169gat), .A4(new_n916_), .ZN(new_n928_));
  AND3_X1   g727(.A1(new_n923_), .A2(KEYINPUT62), .A3(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n930_));
  OAI211_X1 g729(.A(KEYINPUT123), .B(new_n930_), .C1(new_n917_), .C2(new_n922_), .ZN(new_n931_));
  OAI21_X1  g730(.A(KEYINPUT124), .B1(new_n876_), .B2(new_n913_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n933_));
  INV_X1    g732(.A(new_n913_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n921_), .A2(new_n933_), .A3(new_n934_), .ZN(new_n935_));
  NAND4_X1  g734(.A1(new_n932_), .A2(new_n935_), .A3(new_n466_), .A4(new_n623_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n931_), .A2(new_n936_), .ZN(new_n937_));
  OAI21_X1  g736(.A(KEYINPUT125), .B1(new_n929_), .B2(new_n937_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n923_), .A2(KEYINPUT62), .A3(new_n928_), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT125), .ZN(new_n940_));
  NAND4_X1  g739(.A1(new_n939_), .A2(new_n940_), .A3(new_n931_), .A4(new_n936_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n938_), .A2(new_n941_), .ZN(G1348gat));
  NOR4_X1   g741(.A1(new_n866_), .A2(new_n454_), .A3(new_n604_), .A4(new_n913_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n932_), .A2(new_n935_), .ZN(new_n944_));
  INV_X1    g743(.A(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n945_), .A2(new_n738_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n943_), .B1(new_n946_), .B2(new_n454_), .ZN(G1349gat));
  NOR3_X1   g746(.A1(new_n866_), .A2(new_n806_), .A3(new_n913_), .ZN(new_n948_));
  OR2_X1    g747(.A1(new_n948_), .A2(G183gat), .ZN(new_n949_));
  OR2_X1    g748(.A1(new_n806_), .A2(new_n476_), .ZN(new_n950_));
  OR3_X1    g749(.A1(new_n944_), .A2(KEYINPUT126), .A3(new_n950_), .ZN(new_n951_));
  OAI21_X1  g750(.A(KEYINPUT126), .B1(new_n944_), .B2(new_n950_), .ZN(new_n952_));
  AND3_X1   g751(.A1(new_n949_), .A2(new_n951_), .A3(new_n952_), .ZN(G1350gat));
  OAI21_X1  g752(.A(G190gat), .B1(new_n944_), .B2(new_n299_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n644_), .A2(new_n457_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n954_), .B1(new_n944_), .B2(new_n955_), .ZN(G1351gat));
  NOR3_X1   g755(.A1(new_n518_), .A2(new_n449_), .A3(new_n421_), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n899_), .A2(new_n623_), .A3(new_n957_), .ZN(new_n958_));
  XNOR2_X1  g757(.A(new_n958_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g758(.A1(new_n899_), .A2(new_n957_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(new_n960_), .A2(new_n604_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(KEYINPUT127), .B(G204gat), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n961_), .A2(new_n962_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n964_));
  OAI21_X1  g763(.A(new_n963_), .B1(new_n961_), .B2(new_n964_), .ZN(G1353gat));
  INV_X1    g764(.A(new_n960_), .ZN(new_n966_));
  XOR2_X1   g765(.A(KEYINPUT63), .B(G211gat), .Z(new_n967_));
  NAND3_X1  g766(.A1(new_n966_), .A2(new_n353_), .A3(new_n967_), .ZN(new_n968_));
  NOR2_X1   g767(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n969_));
  OAI21_X1  g768(.A(new_n969_), .B1(new_n960_), .B2(new_n806_), .ZN(new_n970_));
  AND2_X1   g769(.A1(new_n968_), .A2(new_n970_), .ZN(G1354gat));
  OR3_X1    g770(.A1(new_n960_), .A2(G218gat), .A3(new_n643_), .ZN(new_n972_));
  OAI21_X1  g771(.A(G218gat), .B1(new_n960_), .B2(new_n299_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n972_), .A2(new_n973_), .ZN(G1355gat));
endmodule


