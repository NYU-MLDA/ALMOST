//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n854_, new_n856_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_;
  NAND2_X1  g000(.A1(KEYINPUT78), .A2(G190gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT25), .ZN(new_n203_));
  AOI22_X1  g002(.A1(new_n202_), .A2(KEYINPUT26), .B1(new_n203_), .B2(G183gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT77), .B1(new_n203_), .B2(G183gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT26), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n206_), .A2(KEYINPUT78), .A3(G190gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT77), .ZN(new_n208_));
  INV_X1    g007(.A(G183gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n208_), .A2(new_n209_), .A3(KEYINPUT25), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n204_), .A2(new_n205_), .A3(new_n207_), .A4(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G169gat), .ZN(new_n213_));
  INV_X1    g012(.A(G176gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(KEYINPUT24), .A3(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT24), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n217_), .A2(new_n220_), .A3(new_n221_), .A4(new_n223_), .ZN(new_n224_));
  AND2_X1   g023(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT79), .B(G176gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  OR2_X1    g028(.A1(G183gat), .A2(G190gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n220_), .A2(new_n230_), .A3(new_n221_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(new_n216_), .ZN(new_n232_));
  OAI22_X1  g031(.A1(new_n212_), .A2(new_n224_), .B1(new_n229_), .B2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT30), .ZN(new_n234_));
  INV_X1    g033(.A(G127gat), .ZN(new_n235_));
  INV_X1    g034(.A(G134gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(G120gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(G113gat), .ZN(new_n239_));
  INV_X1    g038(.A(G113gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(G120gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G127gat), .A2(G134gat), .ZN(new_n242_));
  AND4_X1   g041(.A1(new_n237_), .A2(new_n239_), .A3(new_n241_), .A4(new_n242_), .ZN(new_n243_));
  AOI22_X1  g042(.A1(new_n239_), .A2(new_n241_), .B1(new_n237_), .B2(new_n242_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n234_), .B(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(G71gat), .B(G99gat), .Z(new_n248_));
  NAND2_X1  g047(.A1(G227gat), .A2(G233gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n247_), .B(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G15gat), .B(G43gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n252_), .B(new_n253_), .Z(new_n254_));
  XNOR2_X1  g053(.A(new_n251_), .B(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT91), .B(KEYINPUT27), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n223_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT25), .B(G183gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT26), .B(G190gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n216_), .A2(KEYINPUT24), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT84), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT84), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n216_), .A2(new_n264_), .A3(KEYINPUT24), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n263_), .A2(new_n215_), .A3(new_n265_), .ZN(new_n266_));
  OR2_X1    g065(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(KEYINPUT85), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT85), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n270_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n228_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n272_));
  OAI22_X1  g071(.A1(new_n261_), .A2(new_n266_), .B1(new_n272_), .B2(new_n232_), .ZN(new_n273_));
  INV_X1    g072(.A(G197gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n274_), .A2(G204gat), .ZN(new_n275_));
  INV_X1    g074(.A(G204gat), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n276_), .A2(G197gat), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT21), .B1(new_n275_), .B2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(G197gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n274_), .A2(G204gat), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT21), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G211gat), .B(G218gat), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n278_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n283_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n281_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n284_), .A2(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT87), .B1(new_n273_), .B2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT20), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n290_), .B1(new_n233_), .B2(new_n288_), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n284_), .A2(new_n287_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n269_), .A2(new_n271_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n228_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n232_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT87), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n263_), .A2(new_n215_), .A3(new_n265_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n299_), .A2(new_n257_), .A3(new_n260_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n292_), .A2(new_n297_), .A3(new_n298_), .A4(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n289_), .A2(new_n291_), .A3(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G226gat), .A2(G233gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT19), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n273_), .A2(new_n288_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT86), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n224_), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n227_), .A2(new_n228_), .ZN(new_n311_));
  AOI22_X1  g110(.A1(new_n310_), .A2(new_n211_), .B1(new_n296_), .B2(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n290_), .B1(new_n312_), .B2(new_n292_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n273_), .A2(KEYINPUT86), .A3(new_n288_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n309_), .A2(new_n313_), .A3(new_n304_), .A4(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n306_), .A2(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(G64gat), .B(G92gat), .Z(new_n317_));
  XNOR2_X1  g116(.A(G8gat), .B(G36gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n316_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n321_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n306_), .A2(new_n315_), .A3(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n256_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n323_), .B1(new_n306_), .B2(new_n315_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n309_), .A2(new_n313_), .A3(new_n305_), .A4(new_n314_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT20), .B1(new_n312_), .B2(new_n292_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n273_), .A2(new_n288_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n304_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n321_), .B1(new_n327_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT27), .ZN(new_n332_));
  NOR3_X1   g131(.A1(new_n326_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n325_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT92), .ZN(new_n335_));
  XOR2_X1   g134(.A(G78gat), .B(G106gat), .Z(new_n336_));
  NOR2_X1   g135(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n337_));
  INV_X1    g136(.A(G141gat), .ZN(new_n338_));
  INV_X1    g137(.A(G148gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  OAI22_X1  g139(.A1(KEYINPUT81), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G141gat), .A2(G148gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT2), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n340_), .A2(new_n341_), .A3(new_n344_), .A4(new_n345_), .ZN(new_n346_));
  XOR2_X1   g145(.A(G155gat), .B(G162gat), .Z(new_n347_));
  INV_X1    g146(.A(G155gat), .ZN(new_n348_));
  INV_X1    g147(.A(G162gat), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT1), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT1), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(G155gat), .A3(G162gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n348_), .A2(new_n349_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n350_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(G141gat), .B(G148gat), .Z(new_n355_));
  AOI22_X1  g154(.A1(new_n346_), .A2(new_n347_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT29), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n288_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G228gat), .A2(G233gat), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT82), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n358_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n359_), .A2(new_n360_), .ZN(new_n363_));
  AND2_X1   g162(.A1(new_n358_), .A2(new_n363_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n336_), .B(new_n362_), .C1(new_n364_), .C2(new_n361_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n336_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n362_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n361_), .B1(new_n358_), .B2(new_n363_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n366_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n365_), .A2(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n362_), .B1(new_n364_), .B2(new_n361_), .ZN(new_n371_));
  AOI21_X1  g170(.A(KEYINPUT83), .B1(new_n371_), .B2(new_n366_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT28), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n373_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n356_), .A2(new_n373_), .A3(new_n357_), .ZN(new_n376_));
  XOR2_X1   g175(.A(G22gat), .B(G50gat), .Z(new_n377_));
  AND3_X1   g176(.A1(new_n375_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n377_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n379_));
  OR2_X1    g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n370_), .B1(new_n372_), .B2(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n378_), .A2(new_n379_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n382_), .A2(new_n369_), .A3(new_n365_), .A4(KEYINPUT83), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G225gat), .A2(G233gat), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n346_), .A2(new_n347_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n354_), .A2(new_n355_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n246_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n356_), .A2(new_n245_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n390_), .A2(KEYINPUT90), .A3(new_n391_), .A4(KEYINPUT4), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n245_), .A2(new_n388_), .A3(new_n387_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n237_), .A2(new_n239_), .A3(new_n241_), .A4(new_n242_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n239_), .A2(new_n241_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n237_), .A2(new_n242_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n387_), .A2(new_n388_), .B1(new_n394_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT4), .ZN(new_n399_));
  NOR3_X1   g198(.A1(new_n393_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT90), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n401_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n386_), .B(new_n392_), .C1(new_n400_), .C2(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n393_), .A2(new_n398_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(new_n385_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(G1gat), .B(G29gat), .Z(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(G85gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT0), .B(G57gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n406_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n403_), .A2(new_n410_), .A3(new_n405_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n334_), .A2(new_n335_), .A3(new_n384_), .A4(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n327_), .A2(new_n330_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(new_n323_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n322_), .A2(new_n419_), .A3(KEYINPUT27), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n306_), .A2(new_n323_), .A3(new_n315_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n421_), .A2(new_n326_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n420_), .B1(new_n422_), .B2(new_n256_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n381_), .A2(new_n412_), .A3(new_n414_), .A4(new_n383_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT92), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n417_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT33), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n414_), .A2(new_n427_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n403_), .A2(new_n405_), .A3(KEYINPUT33), .A4(new_n410_), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n385_), .B(new_n392_), .C1(new_n400_), .C2(new_n402_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n404_), .A2(new_n386_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(new_n411_), .A3(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT89), .B1(new_n322_), .B2(new_n324_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT89), .ZN(new_n435_));
  NOR3_X1   g234(.A1(new_n421_), .A2(new_n326_), .A3(new_n435_), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n430_), .B(new_n433_), .C1(new_n434_), .C2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n418_), .A2(KEYINPUT32), .A3(new_n321_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT32), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n316_), .B1(new_n439_), .B2(new_n323_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n438_), .B(new_n440_), .C1(new_n413_), .C2(new_n415_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n384_), .B1(new_n437_), .B2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n255_), .B1(new_n426_), .B2(new_n442_), .ZN(new_n443_));
  XOR2_X1   g242(.A(new_n251_), .B(new_n254_), .Z(new_n444_));
  INV_X1    g243(.A(KEYINPUT93), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n445_), .B1(new_n423_), .B2(new_n384_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n384_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(KEYINPUT93), .A3(new_n334_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n444_), .A2(new_n446_), .A3(new_n416_), .A4(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n443_), .A2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G29gat), .B(G36gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(G50gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT69), .B(G43gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(G50gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n451_), .B(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n453_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n454_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G15gat), .B(G22gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G1gat), .A2(G8gat), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT71), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n461_), .A2(new_n462_), .A3(KEYINPUT14), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n462_), .B1(new_n461_), .B2(KEYINPUT14), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n460_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G1gat), .B(G8gat), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n466_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n459_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n459_), .A2(new_n470_), .ZN(new_n473_));
  OAI211_X1 g272(.A(G229gat), .B(G233gat), .C1(new_n472_), .C2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G229gat), .A2(G233gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n475_), .B(KEYINPUT76), .Z(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n454_), .A2(new_n458_), .A3(KEYINPUT15), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT15), .B1(new_n454_), .B2(new_n458_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  OAI211_X1 g279(.A(new_n471_), .B(new_n477_), .C1(new_n480_), .C2(new_n470_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n474_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G113gat), .B(G141gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G169gat), .B(G197gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n482_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n485_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n474_), .A2(new_n481_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n450_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT94), .ZN(new_n491_));
  XOR2_X1   g290(.A(G190gat), .B(G218gat), .Z(new_n492_));
  XNOR2_X1  g291(.A(G134gat), .B(G162gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT36), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT36), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G99gat), .A2(G106gat), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT6), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT65), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n497_), .B(KEYINPUT6), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT65), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n500_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT9), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n505_), .A2(G85gat), .A3(G92gat), .ZN(new_n506_));
  XOR2_X1   g305(.A(KEYINPUT10), .B(G99gat), .Z(new_n507_));
  INV_X1    g306(.A(G106gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(G85gat), .B(G92gat), .Z(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT9), .ZN(new_n511_));
  AND4_X1   g310(.A1(new_n504_), .A2(new_n506_), .A3(new_n509_), .A4(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n499_), .A2(KEYINPUT66), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT66), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n501_), .A2(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(G99gat), .A2(G106gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT7), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n513_), .A2(new_n515_), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(new_n510_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT8), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n504_), .A2(new_n517_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT8), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n510_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n512_), .B1(new_n520_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(new_n459_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n504_), .A2(new_n506_), .A3(new_n509_), .A4(new_n511_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n522_), .B1(new_n518_), .B2(new_n510_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n523_), .B1(new_n504_), .B2(new_n517_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n528_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n531_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G232gat), .A2(G233gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT34), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT35), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n527_), .A2(new_n532_), .A3(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n535_), .A2(new_n536_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n539_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n527_), .A2(new_n532_), .A3(new_n541_), .A4(new_n537_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n496_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n495_), .B1(new_n543_), .B2(new_n494_), .ZN(new_n544_));
  AOI21_X1  g343(.A(KEYINPUT70), .B1(new_n540_), .B2(new_n542_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n545_), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n547_), .B(new_n495_), .C1(new_n543_), .C2(new_n494_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT37), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n546_), .A2(new_n548_), .A3(KEYINPUT37), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G231gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n469_), .B(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(G57gat), .B(G64gat), .Z(new_n556_));
  INV_X1    g355(.A(KEYINPUT11), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G57gat), .B(G64gat), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(KEYINPUT11), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(G71gat), .B(G78gat), .Z(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n562_), .B1(KEYINPUT11), .B2(new_n559_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n555_), .B(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT67), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G127gat), .B(G155gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT73), .ZN(new_n571_));
  XOR2_X1   g370(.A(KEYINPUT72), .B(KEYINPUT16), .Z(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G183gat), .B(G211gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(KEYINPUT17), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n575_), .A2(KEYINPUT17), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n569_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n576_), .A2(KEYINPUT74), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n576_), .A2(KEYINPUT74), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n580_), .A2(new_n567_), .A3(new_n581_), .ZN(new_n582_));
  OR3_X1    g381(.A1(new_n579_), .A2(KEYINPUT75), .A3(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT75), .B1(new_n579_), .B2(new_n582_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT13), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT12), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n566_), .A2(KEYINPUT67), .ZN(new_n588_));
  INV_X1    g387(.A(new_n562_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n589_), .B1(new_n558_), .B2(new_n560_), .ZN(new_n590_));
  NOR3_X1   g389(.A1(new_n590_), .A2(new_n564_), .A3(KEYINPUT67), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n588_), .A2(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n587_), .B1(new_n526_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G230gat), .A2(G233gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT64), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n526_), .A2(new_n593_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n531_), .A2(KEYINPUT12), .A3(new_n566_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n594_), .A2(new_n596_), .A3(new_n597_), .A4(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT68), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n568_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n601_), .A2(new_n591_), .ZN(new_n602_));
  AOI21_X1  g401(.A(KEYINPUT12), .B1(new_n531_), .B2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n531_), .A2(new_n602_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT68), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n605_), .A2(new_n606_), .A3(new_n596_), .A4(new_n598_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n600_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n596_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n526_), .A2(new_n593_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n609_), .B1(new_n610_), .B2(new_n604_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT5), .B(G176gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(G204gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G120gat), .B(G148gat), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n613_), .B(new_n614_), .Z(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n608_), .A2(new_n611_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n616_), .B1(new_n608_), .B2(new_n611_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n586_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n619_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(KEYINPUT13), .A3(new_n617_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n553_), .A2(new_n585_), .A3(new_n623_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n491_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(G1gat), .ZN(new_n626_));
  INV_X1    g425(.A(new_n416_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n625_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT38), .ZN(new_n629_));
  INV_X1    g428(.A(new_n585_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n489_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n623_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT95), .ZN(new_n634_));
  INV_X1    g433(.A(new_n450_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n549_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n634_), .A2(new_n637_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n638_), .A2(new_n627_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n629_), .B1(new_n626_), .B2(new_n639_), .ZN(G1324gat));
  INV_X1    g439(.A(G8gat), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n625_), .A2(new_n641_), .A3(new_n423_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n638_), .A2(new_n423_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(G8gat), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n644_), .A2(KEYINPUT39), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n644_), .A2(KEYINPUT39), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n642_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT40), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(G1325gat));
  INV_X1    g448(.A(G15gat), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n650_), .B1(new_n638_), .B2(new_n444_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT41), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n625_), .A2(new_n650_), .A3(new_n444_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1326gat));
  INV_X1    g453(.A(G22gat), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n384_), .A2(new_n655_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT97), .Z(new_n657_));
  NAND2_X1  g456(.A1(new_n625_), .A2(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n655_), .B1(new_n638_), .B2(new_n384_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT96), .B(KEYINPUT42), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n659_), .A2(new_n660_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n658_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT98), .Z(G1327gat));
  NAND3_X1  g463(.A1(new_n443_), .A2(KEYINPUT99), .A3(new_n449_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(new_n553_), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT99), .B1(new_n443_), .B2(new_n449_), .ZN(new_n667_));
  OAI21_X1  g466(.A(KEYINPUT43), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT100), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  OAI211_X1 g469(.A(KEYINPUT100), .B(KEYINPUT43), .C1(new_n666_), .C2(new_n667_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n450_), .A2(new_n553_), .A3(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT101), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n450_), .A2(new_n553_), .A3(KEYINPUT101), .A4(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n670_), .A2(new_n671_), .A3(new_n677_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n632_), .A2(new_n585_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT44), .ZN(new_n681_));
  AOI22_X1  g480(.A1(new_n678_), .A2(new_n679_), .B1(KEYINPUT102), .B2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n678_), .A2(KEYINPUT102), .A3(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(new_n680_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n682_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(KEYINPUT104), .B1(new_n686_), .B2(new_n416_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT104), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT44), .B1(new_n683_), .B2(new_n680_), .ZN(new_n689_));
  OAI211_X1 g488(.A(new_n688_), .B(new_n627_), .C1(new_n689_), .C2(new_n682_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n687_), .A2(G29gat), .A3(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n623_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n630_), .A2(new_n549_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n491_), .A2(new_n692_), .A3(new_n693_), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n416_), .A2(G29gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n691_), .B1(new_n694_), .B2(new_n695_), .ZN(G1328gat));
  OAI21_X1  g495(.A(G36gat), .B1(new_n686_), .B2(new_n334_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n694_), .A2(G36gat), .A3(new_n334_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT45), .Z(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT46), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n697_), .A2(KEYINPUT46), .A3(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1329gat));
  OAI211_X1 g503(.A(G43gat), .B(new_n444_), .C1(new_n689_), .C2(new_n682_), .ZN(new_n705_));
  INV_X1    g504(.A(G43gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n706_), .B1(new_n694_), .B2(new_n255_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT105), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n705_), .A2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g509(.A(G50gat), .B1(new_n686_), .B2(new_n447_), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n694_), .A2(G50gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n711_), .B1(new_n447_), .B2(new_n712_), .ZN(G1331gat));
  NOR2_X1   g512(.A1(new_n692_), .A2(new_n489_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n553_), .ZN(new_n715_));
  AND4_X1   g514(.A1(new_n450_), .A2(new_n714_), .A3(new_n630_), .A4(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(G57gat), .B1(new_n716_), .B2(new_n627_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n637_), .A2(new_n630_), .A3(new_n714_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n718_), .A2(new_n416_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n717_), .B1(G57gat), .B2(new_n719_), .ZN(G1332gat));
  OAI21_X1  g519(.A(G64gat), .B1(new_n718_), .B2(new_n334_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT48), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n334_), .A2(G64gat), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT106), .Z(new_n724_));
  NAND2_X1  g523(.A1(new_n716_), .A2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n722_), .A2(new_n725_), .ZN(G1333gat));
  OAI21_X1  g525(.A(G71gat), .B1(new_n718_), .B2(new_n255_), .ZN(new_n727_));
  XOR2_X1   g526(.A(KEYINPUT107), .B(KEYINPUT49), .Z(new_n728_));
  XNOR2_X1  g527(.A(new_n727_), .B(new_n728_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n255_), .A2(G71gat), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT108), .Z(new_n731_));
  NAND2_X1  g530(.A1(new_n716_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n729_), .A2(new_n732_), .ZN(G1334gat));
  OAI21_X1  g532(.A(G78gat), .B1(new_n718_), .B2(new_n447_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT50), .ZN(new_n735_));
  INV_X1    g534(.A(G78gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n716_), .A2(new_n736_), .A3(new_n384_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1335gat));
  AND3_X1   g537(.A1(new_n693_), .A2(new_n450_), .A3(new_n714_), .ZN(new_n739_));
  AOI21_X1  g538(.A(G85gat), .B1(new_n739_), .B2(new_n627_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n678_), .A2(new_n585_), .A3(new_n714_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n741_), .A2(new_n416_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n740_), .B1(new_n742_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g542(.A(G92gat), .B1(new_n739_), .B2(new_n423_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n741_), .A2(new_n334_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n745_), .B2(G92gat), .ZN(G1337gat));
  OAI21_X1  g545(.A(G99gat), .B1(new_n741_), .B2(new_n255_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n739_), .A2(new_n444_), .A3(new_n507_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g549(.A1(new_n739_), .A2(new_n508_), .A3(new_n384_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n678_), .A2(new_n384_), .A3(new_n585_), .A4(new_n714_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n752_), .A2(new_n753_), .A3(G106gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n752_), .B2(G106gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g556(.A(KEYINPUT55), .B1(new_n600_), .B2(new_n607_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n605_), .A2(KEYINPUT55), .A3(new_n596_), .A4(new_n598_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n605_), .A2(new_n598_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(new_n760_), .B2(new_n596_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n615_), .B1(new_n758_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT56), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n477_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n471_), .B(new_n476_), .C1(new_n480_), .C2(new_n470_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n764_), .A2(new_n765_), .A3(new_n485_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n764_), .A2(new_n765_), .A3(KEYINPUT110), .A4(new_n485_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n768_), .A2(new_n488_), .A3(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT111), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT111), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n768_), .A2(new_n772_), .A3(new_n488_), .A4(new_n769_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT56), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n775_), .B(new_n615_), .C1(new_n758_), .C2(new_n761_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n763_), .A2(new_n617_), .A3(new_n774_), .A4(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT58), .ZN(new_n778_));
  OR2_X1    g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n778_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n553_), .A3(new_n780_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(KEYINPUT112), .A2(KEYINPUT57), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n763_), .A2(new_n489_), .A3(new_n617_), .A4(new_n776_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n774_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n785_));
  AOI211_X1 g584(.A(new_n783_), .B(new_n636_), .C1(new_n784_), .C2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n785_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n782_), .B1(new_n787_), .B2(new_n549_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n781_), .B1(new_n786_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT113), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT113), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n781_), .B(new_n791_), .C1(new_n786_), .C2(new_n788_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n790_), .A2(new_n585_), .A3(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT109), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n715_), .A2(new_n630_), .A3(new_n631_), .A4(new_n692_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(KEYINPUT54), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(KEYINPUT54), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n624_), .A2(KEYINPUT109), .A3(new_n798_), .A4(new_n631_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n796_), .A2(new_n797_), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n793_), .A2(new_n800_), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n444_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n627_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT114), .B1(new_n801_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n806_));
  AOI211_X1 g605(.A(new_n806_), .B(new_n803_), .C1(new_n793_), .C2(new_n800_), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n805_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(G113gat), .B1(new_n808_), .B2(new_n489_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n801_), .A2(new_n804_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT59), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n787_), .A2(new_n549_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n783_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n787_), .A2(new_n549_), .A3(new_n782_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n777_), .B(KEYINPUT58), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n814_), .A2(new_n815_), .B1(new_n816_), .B2(new_n553_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n812_), .B1(new_n817_), .B2(new_n630_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n789_), .A2(KEYINPUT116), .A3(new_n585_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n800_), .A3(new_n819_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(KEYINPUT115), .B(KEYINPUT59), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n820_), .A2(new_n804_), .A3(new_n822_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n811_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n489_), .A2(G113gat), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(KEYINPUT117), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n809_), .B1(new_n824_), .B2(new_n826_), .ZN(G1340gat));
  XOR2_X1   g626(.A(KEYINPUT118), .B(G120gat), .Z(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n692_), .B2(KEYINPUT60), .ZN(new_n830_));
  XOR2_X1   g629(.A(new_n830_), .B(KEYINPUT119), .Z(new_n831_));
  OAI211_X1 g630(.A(new_n808_), .B(new_n831_), .C1(KEYINPUT60), .C2(new_n829_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n824_), .A2(new_n623_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n832_), .B1(new_n833_), .B2(new_n829_), .ZN(G1341gat));
  OAI21_X1  g633(.A(new_n630_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n235_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT120), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n835_), .A2(KEYINPUT120), .A3(new_n235_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n585_), .A2(new_n235_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(KEYINPUT121), .ZN(new_n841_));
  AOI22_X1  g640(.A1(new_n838_), .A2(new_n839_), .B1(new_n824_), .B2(new_n841_), .ZN(G1342gat));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n803_), .B1(new_n793_), .B2(new_n800_), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n823_), .B(new_n553_), .C1(new_n843_), .C2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(G134gat), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n236_), .B(new_n636_), .C1(new_n805_), .C2(new_n807_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT122), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n846_), .A2(new_n847_), .A3(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n848_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1343gat));
  NOR2_X1   g650(.A1(new_n444_), .A2(new_n447_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n801_), .A2(new_n627_), .A3(new_n334_), .A4(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(new_n631_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(new_n338_), .ZN(G1344gat));
  NOR2_X1   g654(.A1(new_n853_), .A2(new_n692_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(new_n339_), .ZN(G1345gat));
  OR3_X1    g656(.A1(new_n853_), .A2(KEYINPUT123), .A3(new_n585_), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT123), .B1(new_n853_), .B2(new_n585_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(KEYINPUT61), .B(G155gat), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n858_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1346gat));
  NOR3_X1   g662(.A1(new_n853_), .A2(new_n349_), .A3(new_n715_), .ZN(new_n864_));
  OR2_X1    g663(.A1(new_n853_), .A2(new_n549_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n349_), .B2(new_n865_), .ZN(G1347gat));
  NAND3_X1  g665(.A1(new_n444_), .A2(new_n416_), .A3(new_n423_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n820_), .A2(new_n447_), .A3(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n213_), .B1(new_n870_), .B2(new_n489_), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n871_), .A2(KEYINPUT62), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n870_), .A2(new_n293_), .A3(new_n489_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(KEYINPUT62), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n872_), .A2(new_n873_), .A3(new_n874_), .ZN(G1348gat));
  AOI21_X1  g674(.A(new_n228_), .B1(new_n870_), .B2(new_n623_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n384_), .B1(new_n793_), .B2(new_n800_), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n877_), .A2(G176gat), .A3(new_n623_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n876_), .B1(new_n868_), .B2(new_n878_), .ZN(G1349gat));
  NOR2_X1   g678(.A1(new_n585_), .A2(new_n867_), .ZN(new_n880_));
  AOI21_X1  g679(.A(G183gat), .B1(new_n877_), .B2(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n869_), .A2(new_n258_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n881_), .B1(new_n882_), .B2(new_n630_), .ZN(G1350gat));
  OAI21_X1  g682(.A(G190gat), .B1(new_n869_), .B2(new_n715_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n636_), .A2(new_n259_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n869_), .B2(new_n885_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(KEYINPUT124), .ZN(G1351gat));
  NOR2_X1   g686(.A1(new_n444_), .A2(new_n424_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n334_), .B1(new_n888_), .B2(KEYINPUT125), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n801_), .B(new_n889_), .C1(KEYINPUT125), .C2(new_n888_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n631_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(new_n274_), .ZN(G1352gat));
  NOR2_X1   g691(.A1(new_n890_), .A2(new_n692_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n276_), .A2(KEYINPUT126), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n893_), .B(new_n894_), .Z(G1353gat));
  NOR2_X1   g694(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n896_), .B1(new_n890_), .B2(new_n585_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT127), .ZN(new_n898_));
  OR2_X1    g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n898_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n890_), .A2(new_n585_), .ZN(new_n901_));
  XOR2_X1   g700(.A(KEYINPUT63), .B(G211gat), .Z(new_n902_));
  AOI22_X1  g701(.A1(new_n899_), .A2(new_n900_), .B1(new_n901_), .B2(new_n902_), .ZN(G1354gat));
  NOR2_X1   g702(.A1(new_n890_), .A2(new_n549_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(G218gat), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n890_), .A2(new_n715_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n905_), .B1(G218gat), .B2(new_n906_), .ZN(G1355gat));
endmodule


