//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n877_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n914_, new_n916_, new_n917_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_, new_n940_;
  XNOR2_X1  g000(.A(G22gat), .B(G50gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT89), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  XOR2_X1   g006(.A(new_n207_), .B(KEYINPUT3), .Z(new_n208_));
  NAND2_X1  g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  XOR2_X1   g008(.A(new_n209_), .B(KEYINPUT2), .Z(new_n210_));
  OAI211_X1 g009(.A(new_n205_), .B(new_n206_), .C1(new_n208_), .C2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT1), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n206_), .B(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n205_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n207_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n209_), .A3(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n211_), .A2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT28), .B1(new_n217_), .B2(KEYINPUT29), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  NOR3_X1   g018(.A1(new_n217_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n203_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n220_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(new_n218_), .A3(new_n202_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT90), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT21), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G197gat), .B(G204gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT92), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G211gat), .B(G218gat), .ZN(new_n229_));
  AOI211_X1 g028(.A(new_n226_), .B(new_n227_), .C1(new_n228_), .C2(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n230_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT91), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n227_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT21), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n227_), .A2(new_n232_), .A3(new_n226_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(new_n229_), .A3(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n225_), .B1(new_n231_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G228gat), .A2(G233gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n217_), .A2(KEYINPUT29), .ZN(new_n239_));
  AND3_X1   g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n238_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT93), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(G78gat), .B(G106gat), .Z(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n224_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n244_), .B1(new_n224_), .B2(new_n242_), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n240_), .A2(new_n241_), .ZN(new_n248_));
  OAI22_X1  g047(.A1(new_n246_), .A2(new_n247_), .B1(KEYINPUT93), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n247_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n248_), .A2(KEYINPUT93), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(new_n251_), .A3(new_n245_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n249_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G127gat), .B(G134gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G113gat), .B(G120gat), .ZN(new_n256_));
  OR2_X1    g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n256_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n211_), .A2(new_n216_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT98), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n257_), .A2(KEYINPUT88), .A3(new_n258_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT88), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n255_), .A2(new_n256_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n217_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G225gat), .A2(G233gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT98), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n211_), .A2(new_n216_), .A3(new_n268_), .A4(new_n259_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n261_), .A2(new_n266_), .A3(new_n267_), .A4(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT101), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(new_n267_), .B(KEYINPUT99), .Z(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n266_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n274_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n261_), .A2(new_n266_), .A3(KEYINPUT4), .A4(new_n269_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT100), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT100), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n277_), .A2(new_n281_), .A3(new_n278_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n272_), .A2(new_n280_), .A3(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G1gat), .B(G29gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(G85gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT0), .B(G57gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n283_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n287_), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n272_), .A2(new_n280_), .A3(new_n289_), .A4(new_n282_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G227gat), .A2(G233gat), .ZN(new_n292_));
  INV_X1    g091(.A(G15gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT30), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT31), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G183gat), .A2(G190gat), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n298_), .A2(KEYINPUT23), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT86), .B(KEYINPUT23), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n299_), .B1(new_n300_), .B2(new_n298_), .ZN(new_n301_));
  INV_X1    g100(.A(G169gat), .ZN(new_n302_));
  INV_X1    g101(.A(G176gat), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT24), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n304_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n303_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n306_), .A2(KEYINPUT24), .ZN(new_n307_));
  NOR3_X1   g106(.A1(new_n301_), .A2(new_n305_), .A3(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(G190gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT26), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT85), .ZN(new_n311_));
  NAND2_X1  g110(.A1(KEYINPUT84), .A2(G183gat), .ZN(new_n312_));
  AOI22_X1  g111(.A1(new_n310_), .A2(new_n311_), .B1(KEYINPUT25), .B2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n313_), .B1(new_n311_), .B2(new_n310_), .ZN(new_n314_));
  OAI22_X1  g113(.A1(new_n312_), .A2(KEYINPUT25), .B1(new_n309_), .B2(KEYINPUT26), .ZN(new_n315_));
  OR2_X1    g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  OR3_X1    g115(.A1(new_n300_), .A2(KEYINPUT87), .A3(new_n298_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(G183gat), .A2(G190gat), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n298_), .A2(KEYINPUT23), .ZN(new_n320_));
  OAI211_X1 g119(.A(KEYINPUT87), .B(new_n320_), .C1(new_n300_), .C2(new_n298_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n317_), .A2(new_n319_), .A3(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(G169gat), .ZN(new_n324_));
  AOI22_X1  g123(.A1(new_n308_), .A2(new_n316_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G71gat), .B(G99gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(G43gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n325_), .B(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n265_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n328_), .A2(new_n329_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n297_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n332_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n334_), .A2(new_n296_), .A3(new_n330_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n291_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT20), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n231_), .A2(new_n236_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n339_), .B1(new_n340_), .B2(new_n325_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n231_), .A2(new_n236_), .ZN(new_n342_));
  AOI22_X1  g141(.A1(new_n304_), .A2(KEYINPUT95), .B1(new_n302_), .B2(new_n303_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n343_), .B1(KEYINPUT95), .B2(new_n304_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT26), .B(G190gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT25), .B(G183gat), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n307_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n344_), .A2(new_n321_), .A3(new_n317_), .A4(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n324_), .B1(new_n301_), .B2(new_n318_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n342_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT96), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT96), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n342_), .A2(new_n350_), .A3(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n341_), .A2(new_n352_), .A3(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G226gat), .A2(G233gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n355_), .A2(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n340_), .A2(new_n325_), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT20), .B1(new_n342_), .B2(new_n350_), .ZN(new_n362_));
  OR3_X1    g161(.A1(new_n361_), .A2(new_n362_), .A3(new_n359_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n360_), .A2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G8gat), .B(G36gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT18), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G64gat), .B(G92gat), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n366_), .B(new_n367_), .Z(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n364_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n360_), .A2(new_n363_), .A3(new_n368_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(KEYINPUT97), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT97), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n360_), .A2(new_n363_), .A3(new_n373_), .A4(new_n368_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT103), .B(KEYINPUT27), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n372_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n359_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n377_), .B1(new_n355_), .B2(new_n359_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(new_n369_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(KEYINPUT27), .A3(new_n371_), .ZN(new_n380_));
  AND4_X1   g179(.A1(new_n254_), .A2(new_n338_), .A3(new_n376_), .A4(new_n380_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n288_), .A2(new_n290_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n376_), .A2(new_n253_), .A3(new_n382_), .A4(new_n380_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n368_), .A2(KEYINPUT32), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n378_), .A2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n360_), .A2(new_n363_), .A3(new_n384_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n388_), .B1(new_n290_), .B2(new_n288_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT33), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n290_), .A2(new_n390_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n277_), .A2(new_n281_), .A3(new_n278_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n281_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n394_), .A2(KEYINPUT33), .A3(new_n289_), .A4(new_n272_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n261_), .A2(new_n266_), .A3(new_n269_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n287_), .B1(new_n396_), .B2(new_n274_), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n397_), .A2(KEYINPUT102), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n275_), .A2(new_n276_), .B1(G225gat), .B2(G233gat), .ZN(new_n399_));
  AOI22_X1  g198(.A1(new_n397_), .A2(KEYINPUT102), .B1(new_n399_), .B2(new_n278_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n391_), .A2(new_n395_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n372_), .A2(new_n374_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n389_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n383_), .B1(new_n404_), .B2(new_n253_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n381_), .B1(new_n405_), .B2(new_n337_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G113gat), .B(G141gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G169gat), .B(G197gat), .ZN(new_n408_));
  XOR2_X1   g207(.A(new_n407_), .B(new_n408_), .Z(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT71), .B(KEYINPUT15), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G29gat), .B(G36gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT69), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT69), .ZN(new_n415_));
  INV_X1    g214(.A(G29gat), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n416_), .A2(G36gat), .ZN(new_n417_));
  INV_X1    g216(.A(G36gat), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n418_), .A2(G29gat), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n415_), .B1(new_n417_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n414_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(G43gat), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n422_), .A2(G50gat), .ZN(new_n423_));
  INV_X1    g222(.A(G50gat), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n424_), .A2(G43gat), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT70), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(G43gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n422_), .A2(G50gat), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT70), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n426_), .A2(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n421_), .A2(new_n431_), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n414_), .A2(new_n420_), .B1(new_n426_), .B2(new_n430_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n412_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n421_), .A2(new_n431_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n414_), .A2(new_n420_), .A3(new_n426_), .A4(new_n430_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n435_), .A2(new_n436_), .A3(new_n411_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n434_), .A2(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(G1gat), .B(G8gat), .Z(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G15gat), .B(G22gat), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT77), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G1gat), .A2(G8gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT14), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n441_), .A2(new_n442_), .A3(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n442_), .B1(new_n441_), .B2(new_n444_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n440_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n447_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(new_n439_), .A3(new_n445_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n438_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n435_), .A2(new_n436_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G229gat), .A2(G233gat), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n452_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n457_), .A2(KEYINPUT82), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT82), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n452_), .A2(new_n455_), .A3(new_n459_), .A4(new_n456_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n456_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n451_), .A2(new_n453_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n461_), .B1(new_n462_), .B2(new_n454_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n460_), .A2(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n410_), .B1(new_n458_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT83), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n457_), .A2(KEYINPUT82), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n467_), .A2(new_n463_), .A3(new_n460_), .A4(new_n409_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n465_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n469_));
  OAI211_X1 g268(.A(KEYINPUT83), .B(new_n410_), .C1(new_n458_), .C2(new_n464_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n406_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT66), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT66), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT6), .ZN(new_n476_));
  AND2_X1   g275(.A1(G99gat), .A2(G106gat), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n474_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n477_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT65), .B(G85gat), .ZN(new_n481_));
  INV_X1    g280(.A(G92gat), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n482_), .A2(KEYINPUT9), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  OR2_X1    g283(.A1(G85gat), .A2(G92gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G85gat), .A2(G92gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(KEYINPUT9), .A3(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT64), .B(G106gat), .ZN(new_n488_));
  OR2_X1    g287(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n488_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n480_), .A2(new_n484_), .A3(new_n487_), .A4(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n475_), .A2(KEYINPUT6), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n473_), .A2(KEYINPUT66), .ZN(new_n494_));
  INV_X1    g293(.A(G99gat), .ZN(new_n495_));
  INV_X1    g294(.A(G106gat), .ZN(new_n496_));
  OAI22_X1  g295(.A1(new_n493_), .A2(new_n494_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NOR3_X1   g298(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n474_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n497_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT8), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n485_), .A2(new_n486_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n503_), .A2(new_n504_), .A3(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n504_), .B1(new_n503_), .B2(new_n506_), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n453_), .B(new_n492_), .C1(new_n507_), .C2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n491_), .A2(new_n484_), .A3(new_n487_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n497_), .A2(new_n502_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT7), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n513_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(new_n498_), .ZN(new_n515_));
  NOR3_X1   g314(.A1(new_n478_), .A2(new_n479_), .A3(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT8), .B1(new_n516_), .B2(new_n505_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n503_), .A2(new_n504_), .A3(new_n506_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n512_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n509_), .B1(new_n438_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT72), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT35), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n509_), .B(new_n523_), .C1(new_n438_), .C2(new_n519_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G232gat), .A2(G233gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n522_), .A2(new_n524_), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n527_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n520_), .A2(new_n521_), .A3(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(G190gat), .B(G218gat), .Z(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT73), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G134gat), .B(G162gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT36), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n531_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT36), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n535_), .A2(new_n538_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n537_), .B(KEYINPUT74), .C1(new_n531_), .C2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT37), .ZN(new_n541_));
  INV_X1    g340(.A(new_n536_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n542_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT74), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n541_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n540_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT75), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n531_), .A2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n528_), .A2(KEYINPUT75), .A3(new_n530_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n548_), .A2(new_n536_), .A3(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n531_), .A2(new_n539_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n550_), .A2(new_n541_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT76), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n542_), .B1(new_n531_), .B2(new_n547_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n551_), .B1(new_n555_), .B2(new_n549_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT76), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n556_), .A2(new_n557_), .A3(new_n541_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n546_), .B1(new_n554_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT81), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G57gat), .B(G64gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT11), .ZN(new_n563_));
  XOR2_X1   g362(.A(G71gat), .B(G78gat), .Z(new_n564_));
  OR2_X1    g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n562_), .A2(KEYINPUT11), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n564_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n565_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n568_), .B(new_n569_), .Z(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(new_n451_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n568_), .B(new_n569_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n572_), .A2(new_n450_), .A3(new_n448_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n561_), .B1(new_n571_), .B2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT80), .ZN(new_n576_));
  XOR2_X1   g375(.A(G127gat), .B(G155gat), .Z(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G183gat), .B(G211gat), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n579_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n580_), .A2(KEYINPUT17), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(KEYINPUT17), .B1(new_n580_), .B2(new_n581_), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n574_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n571_), .A2(new_n561_), .A3(new_n573_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n571_), .A2(new_n573_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT78), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n582_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n571_), .A2(KEYINPUT78), .A3(new_n573_), .ZN(new_n590_));
  AOI22_X1  g389(.A1(new_n585_), .A2(new_n586_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n560_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT13), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G230gat), .A2(G233gat), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  OAI211_X1 g394(.A(new_n568_), .B(new_n492_), .C1(new_n507_), .C2(new_n508_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT67), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n517_), .A2(new_n518_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n599_), .A2(KEYINPUT67), .A3(new_n568_), .A4(new_n492_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n519_), .A2(new_n568_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n595_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n595_), .B1(new_n519_), .B2(new_n568_), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n519_), .A2(KEYINPUT12), .A3(new_n568_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT12), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n492_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n568_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n606_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n604_), .B1(new_n605_), .B2(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(G120gat), .B(G148gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT5), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G176gat), .B(G204gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT68), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n603_), .A2(new_n610_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n615_), .B1(new_n603_), .B2(new_n610_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n593_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n618_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(KEYINPUT13), .A3(new_n616_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n592_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n472_), .A2(new_n624_), .ZN(new_n625_));
  OR3_X1    g424(.A1(new_n625_), .A2(G1gat), .A3(new_n382_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT38), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n406_), .A2(new_n556_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n591_), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n623_), .A2(new_n471_), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n629_), .A2(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G1gat), .B1(new_n632_), .B2(new_n382_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n626_), .A2(new_n627_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n628_), .A2(new_n633_), .A3(new_n634_), .ZN(G1324gat));
  NAND2_X1  g434(.A1(new_n376_), .A2(new_n380_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n625_), .A2(G8gat), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT104), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n639_), .B1(new_n632_), .B2(new_n637_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n629_), .A2(KEYINPUT104), .A3(new_n636_), .A4(new_n631_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(G8gat), .A3(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT39), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT39), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n640_), .A2(new_n644_), .A3(G8gat), .A4(new_n641_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n638_), .B1(new_n643_), .B2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n647_), .ZN(new_n649_));
  AOI211_X1 g448(.A(new_n638_), .B(new_n649_), .C1(new_n643_), .C2(new_n645_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n648_), .A2(new_n650_), .ZN(G1325gat));
  INV_X1    g450(.A(new_n632_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n293_), .B1(new_n652_), .B2(new_n336_), .ZN(new_n653_));
  XOR2_X1   g452(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n654_));
  OR2_X1    g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n654_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n336_), .A2(new_n293_), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n655_), .B(new_n656_), .C1(new_n625_), .C2(new_n657_), .ZN(G1326gat));
  OAI21_X1  g457(.A(G22gat), .B1(new_n632_), .B2(new_n254_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT42), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n254_), .A2(G22gat), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT107), .Z(new_n662_));
  OAI21_X1  g461(.A(new_n660_), .B1(new_n625_), .B2(new_n662_), .ZN(G1327gat));
  NAND2_X1  g462(.A1(new_n622_), .A2(new_n630_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n556_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n472_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(G29gat), .B1(new_n668_), .B2(new_n291_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n664_), .A2(new_n471_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT108), .Z(new_n671_));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n672_));
  AOI22_X1  g471(.A1(new_n290_), .A2(new_n390_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n403_), .A2(new_n395_), .A3(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n389_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n253_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n383_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n337_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n381_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n672_), .B1(new_n680_), .B2(new_n559_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n406_), .A2(KEYINPUT43), .A3(new_n560_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n671_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n680_), .A2(new_n672_), .A3(new_n559_), .ZN(new_n686_));
  OAI21_X1  g485(.A(KEYINPUT43), .B1(new_n406_), .B2(new_n560_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n688_), .A2(KEYINPUT44), .A3(new_n671_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n685_), .A2(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n382_), .A2(new_n416_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n669_), .B1(new_n690_), .B2(new_n691_), .ZN(G1328gat));
  NAND2_X1  g491(.A1(new_n636_), .A2(new_n418_), .ZN(new_n693_));
  OR3_X1    g492(.A1(new_n667_), .A2(KEYINPUT45), .A3(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(KEYINPUT45), .B1(new_n667_), .B2(new_n693_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n685_), .A2(new_n636_), .A3(new_n689_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n696_), .B1(new_n697_), .B2(new_n418_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT46), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  OAI211_X1 g499(.A(KEYINPUT46), .B(new_n696_), .C1(new_n697_), .C2(new_n418_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1329gat));
  NOR2_X1   g501(.A1(new_n337_), .A2(new_n422_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n685_), .A2(new_n689_), .A3(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT109), .ZN(new_n705_));
  XNOR2_X1  g504(.A(KEYINPUT110), .B(G43gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n706_), .B1(new_n667_), .B2(new_n337_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT111), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n707_), .B(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT109), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n685_), .A2(new_n710_), .A3(new_n689_), .A4(new_n703_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n705_), .A2(new_n709_), .A3(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT47), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT47), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n705_), .A2(new_n709_), .A3(new_n714_), .A4(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1330gat));
  AOI21_X1  g515(.A(G50gat), .B1(new_n668_), .B2(new_n253_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n254_), .A2(new_n424_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n690_), .B2(new_n718_), .ZN(G1331gat));
  NAND2_X1  g518(.A1(new_n680_), .A2(new_n471_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n720_), .A2(new_n622_), .A3(new_n592_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT112), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(G57gat), .B1(new_n723_), .B2(new_n291_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n471_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n622_), .A2(new_n725_), .A3(new_n630_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n629_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(G57gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n729_), .B1(new_n291_), .B2(KEYINPUT113), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n730_), .B1(KEYINPUT113), .B2(new_n729_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n724_), .B1(new_n728_), .B2(new_n731_), .ZN(G1332gat));
  OAI21_X1  g531(.A(G64gat), .B1(new_n727_), .B2(new_n637_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT48), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n637_), .A2(G64gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n722_), .B2(new_n735_), .ZN(G1333gat));
  OAI21_X1  g535(.A(G71gat), .B1(new_n727_), .B2(new_n337_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT49), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n337_), .A2(G71gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n722_), .B2(new_n739_), .ZN(G1334gat));
  OAI21_X1  g539(.A(G78gat), .B1(new_n727_), .B2(new_n254_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT50), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n254_), .A2(G78gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n742_), .B1(new_n722_), .B2(new_n743_), .ZN(G1335gat));
  NOR4_X1   g543(.A1(new_n720_), .A2(new_n622_), .A3(new_n591_), .A4(new_n665_), .ZN(new_n745_));
  AOI21_X1  g544(.A(G85gat), .B1(new_n745_), .B2(new_n291_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n622_), .A2(new_n725_), .A3(new_n591_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n688_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT114), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n688_), .A2(KEYINPUT114), .A3(new_n747_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n291_), .A2(new_n481_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT115), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n746_), .B1(new_n752_), .B2(new_n754_), .ZN(G1336gat));
  NAND3_X1  g554(.A1(new_n745_), .A2(new_n482_), .A3(new_n636_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n637_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n757_), .B2(new_n482_), .ZN(G1337gat));
  NAND4_X1  g557(.A1(new_n745_), .A2(new_n336_), .A3(new_n489_), .A4(new_n490_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n337_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(new_n760_), .B2(new_n495_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT51), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n763_), .B(new_n759_), .C1(new_n760_), .C2(new_n495_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(G1338gat));
  XNOR2_X1  g564(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n766_));
  OAI21_X1  g565(.A(G106gat), .B1(new_n748_), .B2(new_n254_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT52), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n769_), .B(G106gat), .C1(new_n748_), .C2(new_n254_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n745_), .A2(new_n253_), .A3(new_n488_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n766_), .B1(new_n771_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n766_), .ZN(new_n775_));
  AOI211_X1 g574(.A(new_n772_), .B(new_n775_), .C1(new_n768_), .C2(new_n770_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1339gat));
  INV_X1    g576(.A(G113gat), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n603_), .A2(new_n610_), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n779_), .A2(new_n614_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n469_), .A2(new_n780_), .A3(new_n470_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n610_), .A2(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(KEYINPUT12), .B1(new_n519_), .B2(new_n568_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n607_), .A2(new_n606_), .A3(new_n608_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n786_), .A2(KEYINPUT55), .A3(new_n604_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n598_), .A2(new_n600_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n594_), .B1(new_n788_), .B2(new_n786_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT118), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n783_), .B(new_n787_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n605_), .A2(new_n609_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n595_), .B1(new_n792_), .B2(new_n601_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n793_), .A2(KEYINPUT118), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n614_), .B1(new_n791_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT56), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  OAI211_X1 g596(.A(KEYINPUT56), .B(new_n614_), .C1(new_n791_), .C2(new_n794_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n781_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n452_), .A2(new_n461_), .A3(new_n455_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n456_), .B1(new_n462_), .B2(new_n454_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n800_), .A2(new_n410_), .A3(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n468_), .A2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n803_), .B1(new_n620_), .B2(new_n616_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n665_), .B1(new_n799_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT57), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n780_), .A2(new_n468_), .A3(new_n802_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n798_), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n786_), .A2(KEYINPUT55), .A3(new_n604_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT55), .B1(new_n786_), .B2(new_n604_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n793_), .A2(KEYINPUT118), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n789_), .A2(new_n790_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n812_), .A2(new_n813_), .A3(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT56), .B1(new_n815_), .B2(new_n614_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n808_), .B1(new_n809_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT58), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(KEYINPUT58), .B(new_n808_), .C1(new_n809_), .C2(new_n816_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n559_), .A3(new_n820_), .ZN(new_n821_));
  OAI211_X1 g620(.A(KEYINPUT57), .B(new_n665_), .C1(new_n799_), .C2(new_n804_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n807_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n630_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n471_), .A2(new_n619_), .A3(new_n591_), .A4(new_n621_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n825_), .B(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT54), .B1(new_n827_), .B2(new_n559_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n825_), .B(KEYINPUT117), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n560_), .A3(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n828_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n824_), .A2(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n636_), .A2(new_n253_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n834_), .A2(new_n291_), .A3(new_n336_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n833_), .A2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n778_), .B1(new_n837_), .B2(new_n471_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT119), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n838_), .B(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n833_), .A2(KEYINPUT59), .A3(new_n836_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT59), .ZN(new_n842_));
  AOI22_X1  g641(.A1(new_n823_), .A2(new_n630_), .B1(new_n828_), .B2(new_n831_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n835_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n841_), .A2(new_n844_), .A3(KEYINPUT120), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT120), .B1(new_n841_), .B2(new_n844_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n471_), .A2(new_n778_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n840_), .B1(new_n848_), .B2(new_n849_), .ZN(G1340gat));
  AOI21_X1  g649(.A(new_n622_), .B1(new_n841_), .B2(new_n844_), .ZN(new_n851_));
  INV_X1    g650(.A(G120gat), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n852_), .B1(new_n622_), .B2(KEYINPUT60), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(KEYINPUT60), .B2(new_n852_), .ZN(new_n854_));
  OAI22_X1  g653(.A1(new_n851_), .A2(new_n852_), .B1(new_n837_), .B2(new_n854_), .ZN(G1341gat));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n856_));
  AOI21_X1  g655(.A(KEYINPUT59), .B1(new_n833_), .B2(new_n836_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n843_), .A2(new_n842_), .A3(new_n835_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n856_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(G127gat), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n630_), .A2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n859_), .A2(new_n845_), .A3(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n860_), .B1(new_n837_), .B2(new_n630_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(KEYINPUT121), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n862_), .A2(new_n866_), .A3(new_n863_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n867_), .ZN(G1342gat));
  NOR3_X1   g667(.A1(new_n846_), .A2(new_n847_), .A3(new_n560_), .ZN(new_n869_));
  INV_X1    g668(.A(G134gat), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n556_), .A2(new_n870_), .ZN(new_n871_));
  OAI22_X1  g670(.A1(new_n869_), .A2(new_n870_), .B1(new_n837_), .B2(new_n871_), .ZN(G1343gat));
  NAND3_X1  g671(.A1(new_n253_), .A2(new_n291_), .A3(new_n337_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n843_), .A2(new_n636_), .A3(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n725_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n623_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g677(.A1(new_n874_), .A2(new_n591_), .ZN(new_n879_));
  XOR2_X1   g678(.A(KEYINPUT61), .B(G155gat), .Z(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n879_), .B(new_n881_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT122), .B(KEYINPUT123), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n879_), .B(new_n880_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n883_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n884_), .A2(new_n887_), .ZN(G1346gat));
  INV_X1    g687(.A(G162gat), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n874_), .A2(new_n889_), .A3(new_n556_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n874_), .A2(new_n559_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n889_), .ZN(G1347gat));
  INV_X1    g691(.A(KEYINPUT125), .ZN(new_n893_));
  XOR2_X1   g692(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n254_), .A2(new_n338_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n833_), .A2(new_n636_), .A3(new_n725_), .A4(new_n897_), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n302_), .B(new_n895_), .C1(new_n898_), .C2(KEYINPUT22), .ZN(new_n899_));
  NOR4_X1   g698(.A1(new_n843_), .A2(new_n637_), .A3(new_n471_), .A4(new_n896_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT22), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n894_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(G169gat), .B1(new_n898_), .B2(new_n895_), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n893_), .B(new_n899_), .C1(new_n902_), .C2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n895_), .B1(new_n898_), .B2(KEYINPUT22), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n900_), .A2(new_n894_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n906_), .A2(G169gat), .A3(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n893_), .B1(new_n908_), .B2(new_n899_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n905_), .A2(new_n909_), .ZN(G1348gat));
  NOR3_X1   g709(.A1(new_n843_), .A2(new_n637_), .A3(new_n896_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n623_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g712(.A1(new_n911_), .A2(new_n591_), .ZN(new_n914_));
  MUX2_X1   g713(.A(new_n346_), .B(G183gat), .S(new_n914_), .Z(G1350gat));
  NAND3_X1  g714(.A1(new_n911_), .A2(new_n345_), .A3(new_n556_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n911_), .A2(new_n559_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(new_n309_), .ZN(G1351gat));
  NOR3_X1   g717(.A1(new_n254_), .A2(new_n291_), .A3(new_n336_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n833_), .A2(new_n636_), .A3(new_n919_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(KEYINPUT126), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n921_), .A2(G197gat), .A3(new_n725_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(G197gat), .B1(new_n921_), .B2(new_n725_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1352gat));
  NAND2_X1  g724(.A1(new_n921_), .A2(new_n623_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(G204gat), .ZN(new_n927_));
  INV_X1    g726(.A(G204gat), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n921_), .A2(new_n928_), .A3(new_n623_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n929_), .ZN(G1353gat));
  NOR2_X1   g729(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(KEYINPUT127), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n630_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n921_), .A2(new_n932_), .A3(new_n933_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n932_), .B1(new_n921_), .B2(new_n933_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n935_), .A2(new_n936_), .ZN(G1354gat));
  INV_X1    g736(.A(G218gat), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n921_), .A2(new_n938_), .A3(new_n556_), .ZN(new_n939_));
  AND2_X1   g738(.A1(new_n921_), .A2(new_n559_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n940_), .B2(new_n938_), .ZN(G1355gat));
endmodule


