//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n600_, new_n601_, new_n602_, new_n604_, new_n605_, new_n606_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n789_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n803_, new_n804_, new_n805_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n822_, new_n823_, new_n824_, new_n826_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_;
  XOR2_X1   g000(.A(G127gat), .B(G155gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT16), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G183gat), .B(G211gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT17), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT74), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G15gat), .B(G22gat), .ZN(new_n208_));
  INV_X1    g007(.A(G1gat), .ZN(new_n209_));
  INV_X1    g008(.A(G8gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT14), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n208_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G1gat), .B(G8gat), .ZN(new_n213_));
  XOR2_X1   g012(.A(new_n212_), .B(new_n213_), .Z(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n207_), .B(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G231gat), .A2(G233gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n216_), .B(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G57gat), .B(G64gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT11), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT67), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT67), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n219_), .A2(new_n222_), .A3(KEYINPUT11), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n219_), .A2(KEYINPUT11), .ZN(new_n225_));
  XOR2_X1   g024(.A(G71gat), .B(G78gat), .Z(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n224_), .A2(new_n227_), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n221_), .A2(new_n225_), .A3(new_n226_), .A4(new_n223_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n218_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n218_), .A2(new_n230_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n205_), .A2(new_n206_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G232gat), .A2(G233gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT34), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n237_), .A2(KEYINPUT35), .ZN(new_n238_));
  XOR2_X1   g037(.A(G85gat), .B(G92gat), .Z(new_n239_));
  NOR2_X1   g038(.A1(G99gat), .A2(G106gat), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT7), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G99gat), .A2(G106gat), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT6), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n239_), .B1(new_n242_), .B2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT8), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(KEYINPUT66), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n243_), .B(KEYINPUT6), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n242_), .B1(new_n248_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT8), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n239_), .A2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n247_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n248_), .A2(new_n251_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT10), .B(G99gat), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n257_), .A2(G106gat), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n258_), .A2(KEYINPUT65), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(KEYINPUT65), .ZN(new_n260_));
  INV_X1    g059(.A(G85gat), .ZN(new_n261_));
  INV_X1    g060(.A(G92gat), .ZN(new_n262_));
  NOR3_X1   g061(.A1(new_n261_), .A2(new_n262_), .A3(KEYINPUT9), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n263_), .B1(new_n239_), .B2(KEYINPUT9), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n256_), .A2(new_n259_), .A3(new_n260_), .A4(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n255_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G29gat), .B(G36gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G43gat), .B(G50gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  XOR2_X1   g068(.A(KEYINPUT71), .B(KEYINPUT15), .Z(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n266_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n255_), .A2(new_n265_), .A3(new_n269_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n272_), .B1(new_n273_), .B2(KEYINPUT72), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n273_), .A2(KEYINPUT72), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n238_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n276_), .A2(KEYINPUT73), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(KEYINPUT73), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n274_), .A2(new_n275_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n237_), .A2(KEYINPUT35), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n238_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n277_), .A2(new_n278_), .A3(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(G134gat), .B(G162gat), .Z(new_n284_));
  XNOR2_X1  g083(.A(G190gat), .B(G218gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT36), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n286_), .A2(new_n287_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n283_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n278_), .A2(new_n282_), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n291_), .A2(new_n287_), .A3(new_n286_), .A4(new_n277_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT37), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT37), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n293_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G71gat), .B(G99gat), .ZN(new_n299_));
  INV_X1    g098(.A(G43gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G227gat), .A2(G233gat), .ZN(new_n302_));
  INV_X1    g101(.A(G15gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n301_), .B(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(G169gat), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT22), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n308_), .B1(new_n309_), .B2(KEYINPUT76), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT76), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n311_), .A2(KEYINPUT77), .A3(KEYINPUT22), .A4(G169gat), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n310_), .B(new_n312_), .C1(KEYINPUT77), .C2(KEYINPUT22), .ZN(new_n313_));
  INV_X1    g112(.A(G176gat), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n307_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT78), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G183gat), .A2(G190gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT23), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n318_), .B1(G183gat), .B2(G190gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n315_), .A2(KEYINPUT78), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT25), .B(G183gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT75), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT26), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n323_), .B1(new_n324_), .B2(G190gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n322_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT26), .B(G190gat), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n326_), .B1(KEYINPUT75), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n308_), .A2(new_n314_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n330_), .A2(KEYINPUT24), .A3(new_n306_), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n318_), .B(new_n331_), .C1(KEYINPUT24), .C2(new_n330_), .ZN(new_n332_));
  OAI22_X1  g131(.A1(new_n320_), .A2(new_n321_), .B1(new_n329_), .B2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT79), .B(KEYINPUT30), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n333_), .B(new_n334_), .Z(new_n335_));
  AOI21_X1  g134(.A(new_n305_), .B1(new_n335_), .B2(KEYINPUT80), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n335_), .A2(KEYINPUT80), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n336_), .B(new_n337_), .Z(new_n338_));
  XNOR2_X1  g137(.A(G127gat), .B(G134gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G113gat), .B(G120gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT82), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n339_), .A2(new_n340_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n339_), .A2(new_n340_), .A3(KEYINPUT82), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  OR2_X1    g146(.A1(new_n347_), .A2(KEYINPUT31), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(KEYINPUT31), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(KEYINPUT81), .A3(new_n349_), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n338_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n338_), .A2(new_n350_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT86), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT3), .ZN(new_n356_));
  NOR2_X1   g155(.A1(G141gat), .A2(G148gat), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n356_), .B1(new_n357_), .B2(KEYINPUT85), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT85), .ZN(new_n359_));
  NOR3_X1   g158(.A1(new_n359_), .A2(G141gat), .A3(G148gat), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n355_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n357_), .A2(KEYINPUT85), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n359_), .B1(G141gat), .B2(G148gat), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n362_), .A2(KEYINPUT86), .A3(new_n363_), .A4(new_n356_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT87), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n365_), .B1(new_n357_), .B2(new_n356_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G141gat), .A2(G148gat), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT2), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  OAI211_X1 g168(.A(KEYINPUT87), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n370_));
  NAND3_X1  g169(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n361_), .A2(new_n364_), .A3(new_n366_), .A4(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(G155gat), .A2(G162gat), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT83), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G155gat), .A2(G162gat), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT84), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n376_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n373_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n381_), .A2(KEYINPUT1), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT1), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n379_), .A2(new_n385_), .A3(new_n380_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n384_), .A2(new_n376_), .A3(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n357_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n388_), .A2(new_n367_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n383_), .A2(new_n390_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n391_), .A2(KEYINPUT29), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G211gat), .B(G218gat), .ZN(new_n393_));
  INV_X1    g192(.A(G197gat), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT89), .B1(new_n394_), .B2(G204gat), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n393_), .A2(KEYINPUT21), .A3(new_n395_), .ZN(new_n396_));
  XOR2_X1   g195(.A(G197gat), .B(G204gat), .Z(new_n397_));
  OR2_X1    g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n396_), .B(new_n397_), .C1(KEYINPUT21), .C2(new_n393_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT90), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n398_), .A2(new_n399_), .A3(KEYINPUT90), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  AND2_X1   g203(.A1(G228gat), .A2(G233gat), .ZN(new_n405_));
  OR3_X1    g204(.A1(new_n392_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n400_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n405_), .B1(new_n392_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(G78gat), .B(G106gat), .Z(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n409_), .B(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n391_), .A2(KEYINPUT29), .ZN(new_n413_));
  XOR2_X1   g212(.A(G22gat), .B(G50gat), .Z(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n416_));
  XOR2_X1   g215(.A(new_n415_), .B(new_n416_), .Z(new_n417_));
  XNOR2_X1  g216(.A(new_n412_), .B(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  XOR2_X1   g218(.A(KEYINPUT97), .B(KEYINPUT0), .Z(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT98), .ZN(new_n421_));
  XOR2_X1   g220(.A(G1gat), .B(G29gat), .Z(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G57gat), .B(G85gat), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n423_), .B(new_n424_), .Z(new_n425_));
  NAND2_X1  g224(.A1(G225gat), .A2(G233gat), .ZN(new_n426_));
  AOI22_X1  g225(.A1(new_n373_), .A2(new_n382_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n427_));
  NOR3_X1   g226(.A1(new_n427_), .A2(KEYINPUT4), .A3(new_n346_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT95), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n391_), .A2(new_n429_), .A3(new_n347_), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT95), .B1(new_n427_), .B2(new_n346_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n344_), .A2(new_n341_), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n383_), .A2(new_n390_), .A3(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n430_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT4), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n428_), .B1(new_n435_), .B2(KEYINPUT96), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT4), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n383_), .A2(new_n390_), .A3(new_n432_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n438_), .B(KEYINPUT95), .C1(new_n427_), .C2(new_n346_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n437_), .B1(new_n439_), .B2(new_n430_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT96), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n426_), .B1(new_n436_), .B2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n439_), .A2(new_n426_), .A3(new_n430_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n425_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT99), .ZN(new_n447_));
  INV_X1    g246(.A(new_n426_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n428_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n449_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n435_), .A2(KEYINPUT96), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n448_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n425_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n452_), .A2(new_n453_), .A3(new_n444_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n446_), .A2(new_n447_), .A3(new_n454_), .ZN(new_n455_));
  OAI211_X1 g254(.A(KEYINPUT99), .B(new_n425_), .C1(new_n443_), .C2(new_n445_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G226gat), .A2(G233gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT19), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT91), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  AND2_X1   g259(.A1(KEYINPUT92), .A2(KEYINPUT24), .ZN(new_n461_));
  NOR2_X1   g260(.A1(KEYINPUT92), .A2(KEYINPUT24), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n306_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n330_), .A2(KEYINPUT93), .ZN(new_n464_));
  XOR2_X1   g263(.A(new_n463_), .B(new_n464_), .Z(new_n465_));
  NAND2_X1  g264(.A1(new_n327_), .A2(new_n322_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n318_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT22), .B(G169gat), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n307_), .B1(new_n469_), .B2(new_n314_), .ZN(new_n470_));
  AOI22_X1  g269(.A1(new_n465_), .A2(new_n468_), .B1(new_n319_), .B2(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT20), .B1(new_n471_), .B2(new_n407_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n329_), .A2(new_n332_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n320_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n321_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n473_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n472_), .B1(new_n476_), .B2(new_n404_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT20), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n478_), .B1(new_n471_), .B2(new_n407_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n479_), .B1(new_n476_), .B2(new_n404_), .ZN(new_n480_));
  AOI22_X1  g279(.A1(new_n460_), .A2(new_n477_), .B1(new_n480_), .B2(new_n458_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n319_), .A2(new_n470_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n463_), .B(new_n464_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n482_), .B1(new_n483_), .B2(new_n467_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n478_), .B1(new_n484_), .B2(new_n400_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n402_), .A2(new_n403_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n485_), .B1(new_n486_), .B2(new_n333_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(new_n459_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n458_), .ZN(new_n489_));
  OAI211_X1 g288(.A(new_n489_), .B(new_n479_), .C1(new_n476_), .C2(new_n404_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  XOR2_X1   g290(.A(G8gat), .B(G36gat), .Z(new_n492_));
  XNOR2_X1  g291(.A(G64gat), .B(G92gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n494_), .B(new_n495_), .Z(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT32), .ZN(new_n497_));
  MUX2_X1   g296(.A(new_n481_), .B(new_n491_), .S(new_n497_), .Z(new_n498_));
  NAND3_X1  g297(.A1(new_n455_), .A2(new_n456_), .A3(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n453_), .B1(new_n452_), .B2(new_n444_), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n500_), .A2(KEYINPUT33), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n490_), .B(new_n496_), .C1(new_n477_), .C2(new_n460_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n496_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n435_), .A2(KEYINPUT96), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n506_), .A2(new_n442_), .A3(new_n426_), .A4(new_n449_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n425_), .B1(new_n448_), .B2(new_n434_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n505_), .A2(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n510_), .B1(KEYINPUT33), .B2(new_n500_), .ZN(new_n511_));
  AOI22_X1  g310(.A1(new_n499_), .A2(KEYINPUT100), .B1(new_n501_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT100), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n455_), .A2(new_n456_), .A3(new_n513_), .A4(new_n498_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n419_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n455_), .A2(new_n456_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT27), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n517_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n518_));
  OAI211_X1 g317(.A(KEYINPUT27), .B(new_n502_), .C1(new_n481_), .C2(new_n496_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n516_), .A2(new_n418_), .A3(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n354_), .B1(new_n515_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT101), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n518_), .A2(new_n523_), .A3(new_n519_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n523_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n528_), .A2(KEYINPUT102), .A3(new_n418_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT102), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n530_), .B1(new_n419_), .B2(new_n527_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n516_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n529_), .A2(new_n531_), .A3(new_n532_), .A4(new_n353_), .ZN(new_n533_));
  AOI211_X1 g332(.A(new_n235_), .B(new_n298_), .C1(new_n522_), .C2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT12), .ZN(new_n535_));
  INV_X1    g334(.A(new_n230_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n266_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n255_), .A2(new_n230_), .A3(new_n265_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n535_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT12), .B1(new_n266_), .B2(new_n536_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G230gat), .A2(G233gat), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n542_), .B(KEYINPUT64), .Z(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n541_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n537_), .A2(new_n538_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n543_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(G120gat), .B(G148gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(G176gat), .B(G204gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  XOR2_X1   g350(.A(KEYINPUT68), .B(KEYINPUT5), .Z(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n548_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(KEYINPUT69), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n548_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n557_), .A2(KEYINPUT13), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(KEYINPUT13), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT70), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n271_), .A2(new_n215_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n214_), .A2(new_n269_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G229gat), .A2(G233gat), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n214_), .B(new_n269_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n568_), .A2(G229gat), .A3(G233gat), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G113gat), .B(G141gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G169gat), .B(G197gat), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n571_), .B(new_n572_), .Z(new_n573_));
  OR2_X1    g372(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n570_), .A2(new_n573_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n562_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n534_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n580_), .A2(new_n209_), .A3(new_n516_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT38), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n499_), .A2(KEYINPUT100), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n511_), .A2(new_n501_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n583_), .A2(new_n514_), .A3(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n521_), .B1(new_n585_), .B2(new_n418_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n533_), .B1(new_n586_), .B2(new_n353_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n577_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n235_), .A2(new_n294_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(G1gat), .B1(new_n591_), .B2(new_n532_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n582_), .A2(new_n592_), .ZN(G1324gat));
  OAI21_X1  g392(.A(G8gat), .B1(new_n591_), .B2(new_n528_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT39), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n580_), .A2(new_n210_), .A3(new_n527_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT40), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(G1325gat));
  OAI21_X1  g398(.A(G15gat), .B1(new_n591_), .B2(new_n354_), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n600_), .B(KEYINPUT41), .Z(new_n601_));
  NAND3_X1  g400(.A1(new_n580_), .A2(new_n303_), .A3(new_n353_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(G1326gat));
  OAI21_X1  g402(.A(G22gat), .B1(new_n591_), .B2(new_n418_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT42), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n418_), .A2(G22gat), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n605_), .B1(new_n579_), .B2(new_n606_), .ZN(G1327gat));
  AND2_X1   g406(.A1(new_n588_), .A2(new_n235_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n293_), .B(KEYINPUT37), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT43), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT103), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n610_), .B1(new_n298_), .B2(new_n611_), .ZN(new_n612_));
  AOI211_X1 g411(.A(new_n609_), .B(new_n612_), .C1(new_n522_), .C2(new_n533_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n612_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n614_), .B1(new_n587_), .B2(new_n298_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n608_), .B1(new_n613_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT44), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  OAI211_X1 g417(.A(KEYINPUT44), .B(new_n608_), .C1(new_n613_), .C2(new_n615_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n618_), .A2(new_n516_), .A3(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(G29gat), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n234_), .A2(new_n293_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n589_), .A2(new_n622_), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n532_), .A2(G29gat), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n621_), .B1(new_n623_), .B2(new_n624_), .ZN(G1328gat));
  NAND3_X1  g424(.A1(new_n618_), .A2(new_n527_), .A3(new_n619_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(KEYINPUT104), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT104), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n618_), .A2(new_n628_), .A3(new_n527_), .A4(new_n619_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT107), .ZN(new_n630_));
  INV_X1    g429(.A(G36gat), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n627_), .A2(new_n629_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT46), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n589_), .A2(new_n631_), .A3(new_n527_), .A4(new_n622_), .ZN(new_n635_));
  XOR2_X1   g434(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT106), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n630_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n638_), .B1(new_n637_), .B2(new_n635_), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n633_), .A2(new_n634_), .A3(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n634_), .B1(new_n633_), .B2(new_n639_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1329gat));
  NAND4_X1  g441(.A1(new_n618_), .A2(G43gat), .A3(new_n353_), .A4(new_n619_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n300_), .B1(new_n623_), .B2(new_n354_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g445(.A1(new_n623_), .A2(G50gat), .A3(new_n418_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n618_), .A2(new_n419_), .A3(new_n619_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT108), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n648_), .A2(new_n649_), .A3(G50gat), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n648_), .B2(G50gat), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n647_), .B1(new_n650_), .B2(new_n651_), .ZN(G1331gat));
  AND4_X1   g451(.A1(new_n577_), .A2(new_n534_), .A3(new_n559_), .A4(new_n558_), .ZN(new_n653_));
  INV_X1    g452(.A(G57gat), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n653_), .A2(new_n654_), .A3(new_n516_), .ZN(new_n655_));
  AOI211_X1 g454(.A(new_n576_), .B(new_n561_), .C1(new_n522_), .C2(new_n533_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(new_n590_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G57gat), .B1(new_n657_), .B2(new_n532_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n655_), .A2(new_n658_), .ZN(G1332gat));
  OAI21_X1  g458(.A(G64gat), .B1(new_n657_), .B2(new_n528_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT48), .ZN(new_n661_));
  INV_X1    g460(.A(G64gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n653_), .A2(new_n662_), .A3(new_n527_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(G1333gat));
  OAI21_X1  g463(.A(G71gat), .B1(new_n657_), .B2(new_n354_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT49), .ZN(new_n666_));
  INV_X1    g465(.A(G71gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n653_), .A2(new_n667_), .A3(new_n353_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(G1334gat));
  OAI21_X1  g468(.A(G78gat), .B1(new_n657_), .B2(new_n418_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT50), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n418_), .A2(G78gat), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT109), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n653_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n671_), .A2(new_n674_), .ZN(G1335gat));
  NOR2_X1   g474(.A1(new_n613_), .A2(new_n615_), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n676_), .A2(KEYINPUT110), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(KEYINPUT110), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n560_), .A2(new_n234_), .A3(new_n576_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n677_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G85gat), .B1(new_n680_), .B2(new_n532_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n656_), .A2(new_n622_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n682_), .A2(new_n261_), .A3(new_n516_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(G1336gat));
  AOI21_X1  g483(.A(G92gat), .B1(new_n682_), .B2(new_n527_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT111), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n528_), .A2(new_n262_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n686_), .B1(new_n680_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT112), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n686_), .B(KEYINPUT112), .C1(new_n680_), .C2(new_n688_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1337gat));
  NAND2_X1  g492(.A1(new_n656_), .A2(new_n622_), .ZN(new_n694_));
  OR3_X1    g493(.A1(new_n694_), .A2(new_n257_), .A3(new_n354_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n680_), .A2(new_n354_), .ZN(new_n696_));
  INV_X1    g495(.A(G99gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n695_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT51), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT51), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n700_), .B(new_n695_), .C1(new_n696_), .C2(new_n697_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(G1338gat));
  NOR3_X1   g501(.A1(new_n694_), .A2(G106gat), .A3(new_n418_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT113), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n703_), .B(new_n704_), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n419_), .B(new_n679_), .C1(new_n613_), .C2(new_n615_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n706_), .A2(G106gat), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n707_), .A2(KEYINPUT52), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(KEYINPUT52), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n705_), .A2(new_n708_), .A3(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT53), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT53), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n705_), .A2(new_n708_), .A3(new_n712_), .A4(new_n709_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1339gat));
  INV_X1    g513(.A(KEYINPUT117), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n529_), .A2(new_n353_), .A3(new_n531_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT57), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n539_), .A2(new_n543_), .A3(new_n540_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n543_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(KEYINPUT55), .B2(new_n720_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n541_), .A2(KEYINPUT55), .A3(new_n544_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n555_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT56), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT56), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n725_), .B(new_n555_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n724_), .A2(new_n576_), .A3(new_n554_), .A4(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT114), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n548_), .A2(new_n553_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n729_), .B1(new_n723_), .B2(KEYINPUT56), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT114), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n730_), .A2(new_n731_), .A3(new_n576_), .A4(new_n726_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n573_), .B1(new_n568_), .B2(new_n566_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n565_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n734_), .B2(new_n566_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n575_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n557_), .A2(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n728_), .A2(new_n732_), .A3(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n293_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n730_), .A2(KEYINPUT58), .A3(new_n726_), .A4(new_n737_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT116), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n730_), .A2(new_n726_), .A3(new_n737_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(KEYINPUT115), .B(KEYINPUT58), .ZN(new_n744_));
  AOI22_X1  g543(.A1(new_n295_), .A2(new_n297_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  AOI22_X1  g544(.A1(new_n718_), .A2(new_n740_), .B1(new_n742_), .B2(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n739_), .A2(KEYINPUT57), .A3(new_n293_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n234_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n609_), .A2(new_n234_), .A3(new_n577_), .A4(new_n560_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT54), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n749_), .B(new_n750_), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n516_), .B(new_n717_), .C1(new_n748_), .C2(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n715_), .B1(new_n752_), .B2(KEYINPUT59), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n752_), .A2(new_n715_), .A3(KEYINPUT59), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT118), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n757_), .B1(new_n752_), .B2(KEYINPUT59), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n740_), .A2(new_n718_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n742_), .A2(new_n745_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n747_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n235_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n751_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n532_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT59), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n765_), .A2(KEYINPUT118), .A3(new_n766_), .A4(new_n717_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n758_), .A2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n756_), .A2(new_n576_), .A3(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(G113gat), .ZN(new_n770_));
  OR2_X1    g569(.A1(new_n577_), .A2(G113gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n752_), .B2(new_n771_), .ZN(G1340gat));
  INV_X1    g571(.A(new_n755_), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n768_), .B(new_n562_), .C1(new_n753_), .C2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT119), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n756_), .A2(KEYINPUT119), .A3(new_n562_), .A4(new_n768_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(G120gat), .A3(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n752_), .ZN(new_n779_));
  INV_X1    g578(.A(G120gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n780_), .B1(new_n560_), .B2(KEYINPUT60), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n779_), .B(new_n781_), .C1(KEYINPUT60), .C2(new_n780_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n778_), .A2(new_n782_), .ZN(G1341gat));
  AOI21_X1  g582(.A(G127gat), .B1(new_n779_), .B2(new_n234_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n756_), .A2(new_n768_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n234_), .A2(G127gat), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n786_), .B(KEYINPUT120), .Z(new_n787_));
  AOI21_X1  g586(.A(new_n784_), .B1(new_n785_), .B2(new_n787_), .ZN(G1342gat));
  NAND3_X1  g587(.A1(new_n756_), .A2(new_n298_), .A3(new_n768_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(G134gat), .ZN(new_n790_));
  OR2_X1    g589(.A1(new_n293_), .A2(G134gat), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n790_), .B1(new_n752_), .B2(new_n791_), .ZN(G1343gat));
  NOR2_X1   g591(.A1(new_n353_), .A2(new_n418_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n765_), .A2(new_n528_), .A3(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n794_), .A2(new_n577_), .ZN(new_n795_));
  XOR2_X1   g594(.A(new_n795_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g595(.A1(new_n794_), .A2(new_n561_), .ZN(new_n797_));
  XOR2_X1   g596(.A(KEYINPUT121), .B(G148gat), .Z(new_n798_));
  XNOR2_X1  g597(.A(new_n797_), .B(new_n798_), .ZN(G1345gat));
  NOR2_X1   g598(.A1(new_n794_), .A2(new_n235_), .ZN(new_n800_));
  XOR2_X1   g599(.A(KEYINPUT61), .B(G155gat), .Z(new_n801_));
  XNOR2_X1  g600(.A(new_n800_), .B(new_n801_), .ZN(G1346gat));
  OAI21_X1  g601(.A(G162gat), .B1(new_n794_), .B2(new_n609_), .ZN(new_n803_));
  OR2_X1    g602(.A1(new_n293_), .A2(G162gat), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n803_), .B1(new_n794_), .B2(new_n804_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(KEYINPUT122), .ZN(G1347gat));
  NAND2_X1  g605(.A1(new_n763_), .A2(new_n764_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n418_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n354_), .A2(new_n516_), .A3(new_n528_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n809_), .A2(new_n469_), .A3(new_n576_), .A4(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n576_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(KEYINPUT123), .ZN(new_n813_));
  OAI21_X1  g612(.A(G169gat), .B1(new_n808_), .B2(new_n813_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n814_), .A2(KEYINPUT62), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n814_), .A2(KEYINPUT62), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n811_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT124), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(KEYINPUT124), .B(new_n811_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(G1348gat));
  NAND2_X1  g620(.A1(new_n809_), .A2(new_n810_), .ZN(new_n822_));
  OAI21_X1  g621(.A(G176gat), .B1(new_n822_), .B2(new_n561_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n558_), .A2(new_n314_), .A3(new_n559_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n823_), .B1(new_n822_), .B2(new_n824_), .ZN(G1349gat));
  NOR2_X1   g624(.A1(new_n822_), .A2(new_n235_), .ZN(new_n826_));
  MUX2_X1   g625(.A(G183gat), .B(new_n322_), .S(new_n826_), .Z(G1350gat));
  NAND3_X1  g626(.A1(new_n809_), .A2(new_n298_), .A3(new_n810_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n828_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT125), .B1(new_n828_), .B2(G190gat), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n294_), .A2(new_n327_), .ZN(new_n832_));
  OAI22_X1  g631(.A1(new_n830_), .A2(new_n831_), .B1(new_n822_), .B2(new_n832_), .ZN(G1351gat));
  AND4_X1   g632(.A1(new_n532_), .A2(new_n807_), .A3(new_n527_), .A4(new_n793_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n576_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n562_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(KEYINPUT126), .B(G204gat), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n837_), .B(new_n838_), .ZN(G1353gat));
  AOI21_X1  g638(.A(new_n235_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n834_), .A2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n842_));
  XOR2_X1   g641(.A(new_n841_), .B(new_n842_), .Z(G1354gat));
  INV_X1    g642(.A(G218gat), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n834_), .A2(new_n844_), .A3(new_n294_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n834_), .A2(new_n298_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(new_n844_), .ZN(G1355gat));
endmodule


