//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 0 0 0 1 1 1 0 0 0 1 0 0 0 0 0 0 1 0 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n786_, new_n787_, new_n788_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n796_,
    new_n797_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n943_, new_n944_, new_n945_, new_n947_, new_n948_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n960_, new_n961_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n968_, new_n969_, new_n970_,
    new_n971_;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT34), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT35), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G29gat), .B(G36gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G43gat), .B(G50gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT9), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(G85gat), .A3(G92gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  AND2_X1   g011(.A1(G85gat), .A2(G92gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n212_), .B1(KEYINPUT9), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n217_));
  OR2_X1    g016(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n218_));
  INV_X1    g017(.A(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT64), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n218_), .A2(new_n223_), .A3(new_n219_), .A4(new_n220_), .ZN(new_n224_));
  AOI22_X1  g023(.A1(new_n216_), .A2(new_n217_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G85gat), .B(G92gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n211_), .B1(new_n226_), .B2(new_n210_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G99gat), .A2(G106gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT6), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT6), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(G99gat), .A3(G106gat), .ZN(new_n231_));
  AOI22_X1  g030(.A1(new_n227_), .A2(KEYINPUT65), .B1(new_n229_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n225_), .A2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NOR3_X1   g034(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT68), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT7), .ZN(new_n238_));
  INV_X1    g037(.A(G99gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(new_n239_), .A3(new_n219_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(new_n241_), .A3(new_n234_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n229_), .A2(new_n231_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n237_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(new_n215_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(new_n246_), .A3(KEYINPUT8), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n243_), .A2(new_n240_), .A3(new_n234_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT66), .B(KEYINPUT8), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n226_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n248_), .A2(new_n250_), .A3(KEYINPUT67), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n247_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT8), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n257_), .B1(new_n244_), .B2(new_n215_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n258_), .A2(new_n246_), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n209_), .B(new_n233_), .C1(new_n256_), .C2(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n203_), .A2(KEYINPUT35), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  XOR2_X1   g062(.A(new_n207_), .B(new_n208_), .Z(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT15), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT15), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n209_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  AOI22_X1  g067(.A1(new_n258_), .A2(new_n246_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n245_), .A2(KEYINPUT8), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT69), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT70), .ZN(new_n273_));
  AND3_X1   g072(.A1(new_n225_), .A2(new_n273_), .A3(new_n232_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n273_), .B1(new_n225_), .B2(new_n232_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n268_), .B1(new_n272_), .B2(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n206_), .B1(new_n263_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n233_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n279_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n261_), .B1(new_n280_), .B2(new_n209_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n268_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n256_), .A2(new_n259_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n275_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n225_), .A2(new_n273_), .A3(new_n232_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n282_), .B1(new_n283_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n206_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n281_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G190gat), .B(G218gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G134gat), .B(G162gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n292_), .A2(KEYINPUT36), .ZN(new_n293_));
  AND3_X1   g092(.A1(new_n278_), .A2(new_n289_), .A3(new_n293_), .ZN(new_n294_));
  XOR2_X1   g093(.A(new_n292_), .B(KEYINPUT36), .Z(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n296_), .B1(new_n278_), .B2(new_n289_), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT37), .B1(new_n294_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT72), .ZN(new_n299_));
  NOR3_X1   g098(.A1(new_n263_), .A2(new_n277_), .A3(new_n206_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n288_), .B1(new_n281_), .B2(new_n287_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n295_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n278_), .A2(new_n289_), .A3(new_n293_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT72), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(new_n305_), .A3(KEYINPUT37), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n299_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT73), .ZN(new_n308_));
  AND3_X1   g107(.A1(new_n278_), .A2(new_n289_), .A3(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n308_), .B1(new_n278_), .B2(new_n289_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n295_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT74), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT37), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n303_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n311_), .A2(new_n312_), .A3(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT73), .B1(new_n300_), .B2(new_n301_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n278_), .A2(new_n289_), .A3(new_n308_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n296_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT74), .B1(new_n319_), .B2(new_n314_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n307_), .A2(new_n316_), .A3(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G57gat), .B(G64gat), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n322_), .A2(KEYINPUT11), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(KEYINPUT11), .ZN(new_n324_));
  XOR2_X1   g123(.A(G71gat), .B(G78gat), .Z(new_n325_));
  NAND3_X1  g124(.A1(new_n323_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  OR2_X1    g125(.A1(new_n324_), .A2(new_n325_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G15gat), .B(G22gat), .ZN(new_n329_));
  INV_X1    g128(.A(G1gat), .ZN(new_n330_));
  INV_X1    g129(.A(G8gat), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT14), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n329_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G1gat), .B(G8gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n328_), .B(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G231gat), .A2(G233gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT17), .ZN(new_n339_));
  XOR2_X1   g138(.A(G127gat), .B(G155gat), .Z(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT16), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G183gat), .B(G211gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  OR3_X1    g142(.A1(new_n338_), .A2(new_n339_), .A3(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(KEYINPUT17), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n338_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n321_), .A2(new_n348_), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n349_), .B(KEYINPUT75), .Z(new_n350_));
  INV_X1    g149(.A(G183gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT25), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT25), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(G183gat), .ZN(new_n354_));
  INV_X1    g153(.A(G190gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT26), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT26), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(G190gat), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n352_), .A2(new_n354_), .A3(new_n356_), .A4(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  OR3_X1    g162(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n364_));
  OR2_X1    g163(.A1(G169gat), .A2(G176gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G169gat), .A2(G176gat), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(KEYINPUT24), .A3(new_n366_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n359_), .A2(new_n363_), .A3(new_n364_), .A4(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(G169gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G183gat), .A2(G190gat), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT23), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n373_), .B(new_n360_), .C1(G183gat), .C2(G190gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n370_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT80), .ZN(new_n376_));
  AND3_X1   g175(.A1(new_n368_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n376_), .B1(new_n368_), .B2(new_n375_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G227gat), .A2(G233gat), .ZN(new_n380_));
  INV_X1    g179(.A(G15gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT30), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n379_), .B(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(KEYINPUT81), .B(G43gat), .Z(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT82), .ZN(new_n387_));
  INV_X1    g186(.A(G127gat), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n388_), .A2(G134gat), .ZN(new_n389_));
  INV_X1    g188(.A(G134gat), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n390_), .A2(G127gat), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n387_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(G127gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n388_), .A2(G134gat), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n393_), .A2(new_n394_), .A3(KEYINPUT82), .ZN(new_n395_));
  INV_X1    g194(.A(G120gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(G113gat), .ZN(new_n397_));
  INV_X1    g196(.A(G113gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(G120gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n392_), .A2(new_n395_), .A3(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT84), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT84), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n392_), .A2(new_n403_), .A3(new_n395_), .A4(new_n400_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n392_), .A2(new_n395_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n400_), .ZN(new_n406_));
  AOI21_X1  g205(.A(KEYINPUT83), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT83), .ZN(new_n408_));
  AOI211_X1 g207(.A(new_n408_), .B(new_n400_), .C1(new_n392_), .C2(new_n395_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n402_), .B(new_n404_), .C1(new_n407_), .C2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT31), .ZN(new_n411_));
  XOR2_X1   g210(.A(G71gat), .B(G99gat), .Z(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n386_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n386_), .A2(new_n413_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  XOR2_X1   g215(.A(G78gat), .B(G106gat), .Z(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT91), .ZN(new_n418_));
  AND2_X1   g217(.A1(G228gat), .A2(G233gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  XOR2_X1   g219(.A(G22gat), .B(G50gat), .Z(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(G218gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(G211gat), .ZN(new_n424_));
  INV_X1    g223(.A(G211gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(G218gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT90), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT90), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n424_), .A2(new_n426_), .A3(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(G197gat), .A2(G204gat), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G197gat), .A2(G204gat), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(KEYINPUT21), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT21), .ZN(new_n435_));
  INV_X1    g234(.A(new_n433_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n435_), .B1(new_n436_), .B2(new_n431_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n428_), .A2(new_n430_), .A3(new_n434_), .A4(new_n437_), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n436_), .A2(new_n431_), .A3(new_n435_), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n424_), .A2(new_n426_), .A3(new_n429_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n429_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n439_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n438_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G141gat), .A2(G148gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT2), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT2), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n446_), .A2(G141gat), .A3(G148gat), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT3), .ZN(new_n448_));
  NOR2_X1   g247(.A1(G141gat), .A2(G148gat), .ZN(new_n449_));
  AOI22_X1  g248(.A1(new_n445_), .A2(new_n447_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT88), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT88), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n453_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n450_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT89), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n450_), .A2(new_n455_), .A3(KEYINPUT89), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G155gat), .A2(G162gat), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT86), .ZN(new_n462_));
  NOR3_X1   g261(.A1(new_n462_), .A2(G155gat), .A3(G162gat), .ZN(new_n463_));
  INV_X1    g262(.A(G155gat), .ZN(new_n464_));
  INV_X1    g263(.A(G162gat), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT86), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n461_), .B1(new_n463_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n461_), .A2(KEYINPUT1), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n464_), .A2(new_n465_), .A3(KEYINPUT86), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n462_), .B1(G155gat), .B2(G162gat), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n470_), .A2(new_n471_), .B1(KEYINPUT1), .B2(new_n461_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT87), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n469_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n461_), .A2(KEYINPUT1), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n475_), .B1(new_n463_), .B2(new_n466_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT87), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n474_), .A2(new_n477_), .ZN(new_n478_));
  OR2_X1    g277(.A1(new_n449_), .A2(KEYINPUT85), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n449_), .A2(KEYINPUT85), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n479_), .A2(new_n444_), .A3(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  AOI22_X1  g281(.A1(new_n460_), .A2(new_n468_), .B1(new_n478_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT29), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n443_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  AND3_X1   g284(.A1(new_n450_), .A2(new_n455_), .A3(KEYINPUT89), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT89), .B1(new_n450_), .B2(new_n455_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n468_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n473_), .B(new_n475_), .C1(new_n463_), .C2(new_n466_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n469_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n472_), .A2(new_n473_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n482_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n488_), .A2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT28), .B1(new_n494_), .B2(KEYINPUT29), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT28), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n483_), .A2(new_n496_), .A3(new_n484_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n485_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n485_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n422_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n422_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n497_), .A2(new_n495_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n438_), .A2(new_n442_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n504_), .B1(new_n494_), .B2(KEYINPUT29), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n502_), .A2(new_n506_), .A3(new_n498_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n501_), .A2(new_n507_), .ZN(new_n508_));
  XOR2_X1   g307(.A(KEYINPUT95), .B(KEYINPUT0), .Z(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT96), .ZN(new_n510_));
  XOR2_X1   g309(.A(G1gat), .B(G29gat), .Z(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G57gat), .B(G85gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n395_), .ZN(new_n515_));
  AOI21_X1  g314(.A(KEYINPUT82), .B1(new_n393_), .B2(new_n394_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n406_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(new_n401_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n488_), .A2(new_n493_), .A3(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n519_), .B1(new_n483_), .B2(new_n410_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT4), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G225gat), .A2(G233gat), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n402_), .A2(new_n404_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n517_), .A2(new_n408_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n405_), .A2(KEYINPUT83), .A3(new_n406_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n467_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n481_), .B1(new_n474_), .B2(new_n477_), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n524_), .B(new_n527_), .C1(new_n528_), .C2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT4), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n521_), .A2(new_n523_), .A3(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n520_), .A2(new_n522_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n514_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT33), .B1(new_n535_), .B2(KEYINPUT97), .ZN(new_n536_));
  INV_X1    g335(.A(new_n514_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n531_), .B1(new_n530_), .B2(new_n519_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n410_), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT4), .B1(new_n539_), .B2(new_n494_), .ZN(new_n540_));
  NOR3_X1   g339(.A1(new_n538_), .A2(new_n540_), .A3(new_n522_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n534_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n537_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT97), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT33), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G8gat), .B(G36gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G64gat), .B(G92gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n443_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G226gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT20), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n438_), .A2(new_n442_), .A3(new_n368_), .A4(new_n375_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n556_), .B1(new_n557_), .B2(KEYINPUT93), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n368_), .A2(new_n375_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT93), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n504_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n552_), .A2(new_n558_), .A3(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n378_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n368_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n563_), .A2(new_n504_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT20), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n368_), .A2(new_n375_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n566_), .B1(new_n443_), .B2(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n555_), .B1(new_n565_), .B2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n551_), .B1(new_n562_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n555_), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n377_), .A2(new_n378_), .A3(new_n443_), .ZN(new_n572_));
  OAI21_X1  g371(.A(KEYINPUT20), .B1(new_n504_), .B2(new_n559_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n571_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n551_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n552_), .A2(new_n558_), .A3(new_n561_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n574_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n570_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n520_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n537_), .B1(new_n579_), .B2(new_n523_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n522_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n578_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n536_), .A2(new_n546_), .A3(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n533_), .A2(new_n514_), .A3(new_n534_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n543_), .A2(new_n584_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n575_), .A2(KEYINPUT32), .ZN(new_n586_));
  NOR3_X1   g385(.A1(new_n586_), .A2(new_n562_), .A3(new_n569_), .ZN(new_n587_));
  NOR3_X1   g386(.A1(new_n572_), .A2(new_n573_), .A3(new_n571_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n566_), .B1(new_n504_), .B2(new_n559_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n555_), .B1(new_n552_), .B2(new_n589_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n587_), .B1(new_n591_), .B2(new_n586_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n585_), .A2(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n508_), .B1(new_n583_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT98), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n543_), .A2(new_n507_), .A3(new_n501_), .A4(new_n584_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT27), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n578_), .A2(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n551_), .B1(new_n588_), .B2(new_n590_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n599_), .A2(KEYINPUT27), .A3(new_n577_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n595_), .B1(new_n596_), .B2(new_n601_), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n541_), .A2(new_n542_), .A3(new_n537_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n603_), .A2(new_n535_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n577_), .A2(KEYINPUT27), .ZN(new_n605_));
  AOI22_X1  g404(.A1(new_n599_), .A2(new_n605_), .B1(new_n578_), .B2(new_n597_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n604_), .A2(new_n508_), .A3(new_n606_), .A4(KEYINPUT98), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n602_), .A2(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n416_), .B1(new_n594_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n508_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(new_n606_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n611_), .A2(new_n585_), .A3(new_n416_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n609_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n328_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n616_), .B1(new_n283_), .B2(new_n279_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT12), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G230gat), .A2(G233gat), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n280_), .A2(new_n328_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n616_), .A2(KEYINPUT12), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n623_), .B1(new_n283_), .B2(new_n286_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n619_), .A2(new_n620_), .A3(new_n621_), .A4(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n617_), .A2(new_n621_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n626_), .A2(G230gat), .A3(G233gat), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G120gat), .B(G148gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT5), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G176gat), .B(G204gat), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n630_), .B(new_n631_), .Z(new_n632_));
  NAND2_X1  g431(.A1(new_n628_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n632_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n625_), .A2(new_n627_), .A3(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT13), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n637_), .A2(KEYINPUT71), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(KEYINPUT71), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n636_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n633_), .B(new_n635_), .C1(KEYINPUT71), .C2(new_n637_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n335_), .A2(new_n264_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n335_), .A2(new_n264_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(KEYINPUT76), .A3(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(G229gat), .A2(G233gat), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT76), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n335_), .A2(new_n648_), .A3(new_n264_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n645_), .A2(new_n647_), .A3(new_n649_), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n650_), .A2(KEYINPUT77), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n265_), .A2(new_n335_), .A3(new_n267_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT78), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT78), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n265_), .A2(new_n654_), .A3(new_n335_), .A4(new_n267_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n653_), .A2(new_n643_), .A3(new_n655_), .ZN(new_n656_));
  OAI211_X1 g455(.A(KEYINPUT77), .B(new_n650_), .C1(new_n656_), .C2(new_n647_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n651_), .A2(new_n657_), .A3(KEYINPUT79), .ZN(new_n658_));
  XNOR2_X1  g457(.A(G113gat), .B(G141gat), .ZN(new_n659_));
  XNOR2_X1  g458(.A(G169gat), .B(G197gat), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n659_), .B(new_n660_), .Z(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n658_), .A2(new_n662_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n651_), .A2(new_n657_), .A3(KEYINPUT79), .A4(new_n661_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n642_), .A2(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n615_), .A2(new_n666_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n350_), .A2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n668_), .A2(new_n330_), .A3(new_n585_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT99), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT38), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n671_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n319_), .A2(new_n294_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n615_), .A2(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n666_), .A2(new_n347_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(G1gat), .B1(new_n677_), .B2(new_n604_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n672_), .A2(new_n673_), .A3(new_n678_), .ZN(G1324gat));
  INV_X1    g478(.A(KEYINPUT39), .ZN(new_n680_));
  INV_X1    g479(.A(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(new_n601_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n680_), .B1(new_n682_), .B2(G8gat), .ZN(new_n683_));
  AOI211_X1 g482(.A(KEYINPUT39), .B(new_n331_), .C1(new_n681_), .C2(new_n601_), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n668_), .A2(new_n331_), .A3(new_n601_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(G1325gat));
  OAI21_X1  g488(.A(G15gat), .B1(new_n677_), .B2(new_n416_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT41), .Z(new_n691_));
  INV_X1    g490(.A(new_n416_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n668_), .A2(new_n381_), .A3(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1326gat));
  OAI21_X1  g493(.A(G22gat), .B1(new_n677_), .B2(new_n610_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT42), .ZN(new_n696_));
  INV_X1    g495(.A(G22gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n668_), .A2(new_n697_), .A3(new_n508_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(G1327gat));
  INV_X1    g498(.A(new_n674_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n700_), .A2(new_n348_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n667_), .A2(new_n701_), .ZN(new_n702_));
  OR3_X1    g501(.A1(new_n702_), .A2(G29gat), .A3(new_n604_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT103), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n666_), .A2(new_n348_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(KEYINPUT101), .B(KEYINPUT43), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT102), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n320_), .A2(new_n316_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n305_), .B1(new_n304_), .B2(KEYINPUT37), .ZN(new_n709_));
  AOI211_X1 g508(.A(KEYINPUT72), .B(new_n313_), .C1(new_n302_), .C2(new_n303_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n708_), .B2(new_n711_), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n307_), .A2(KEYINPUT102), .A3(new_n316_), .A4(new_n320_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n706_), .B1(new_n714_), .B2(new_n614_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n307_), .A2(new_n716_), .A3(new_n316_), .A4(new_n320_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n717_), .B1(new_n613_), .B2(new_n609_), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n704_), .B(new_n705_), .C1(new_n715_), .C2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n583_), .A2(new_n593_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(new_n610_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n602_), .A2(new_n607_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n692_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n712_), .B(new_n713_), .C1(new_n723_), .C2(new_n612_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n706_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n718_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n705_), .ZN(new_n727_));
  OAI21_X1  g526(.A(KEYINPUT103), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n719_), .A2(new_n728_), .A3(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n724_), .A2(new_n725_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n718_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n727_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT44), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n730_), .A2(new_n585_), .A3(new_n734_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n735_), .A2(KEYINPUT104), .ZN(new_n736_));
  OAI21_X1  g535(.A(G29gat), .B1(new_n735_), .B2(KEYINPUT104), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n703_), .B1(new_n736_), .B2(new_n737_), .ZN(G1328gat));
  NOR3_X1   g537(.A1(new_n702_), .A2(G36gat), .A3(new_n606_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT45), .Z(new_n740_));
  AOI21_X1  g539(.A(new_n606_), .B1(new_n733_), .B2(KEYINPUT44), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n730_), .A2(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(KEYINPUT105), .B1(new_n742_), .B2(G36gat), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT105), .ZN(new_n744_));
  INV_X1    g543(.A(G36gat), .ZN(new_n745_));
  AOI211_X1 g544(.A(new_n744_), .B(new_n745_), .C1(new_n730_), .C2(new_n741_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n740_), .B1(new_n743_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT46), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  OAI211_X1 g548(.A(KEYINPUT46), .B(new_n740_), .C1(new_n743_), .C2(new_n746_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1329gat));
  NAND4_X1  g550(.A1(new_n730_), .A2(G43gat), .A3(new_n692_), .A4(new_n734_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n702_), .A2(new_n416_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n752_), .B1(G43gat), .B2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g554(.A1(new_n730_), .A2(new_n508_), .A3(new_n734_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT106), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n756_), .A2(new_n757_), .A3(G50gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n756_), .B2(G50gat), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n610_), .A2(G50gat), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT107), .Z(new_n761_));
  OAI22_X1  g560(.A1(new_n758_), .A2(new_n759_), .B1(new_n702_), .B2(new_n761_), .ZN(G1331gat));
  NAND2_X1  g561(.A1(new_n663_), .A2(new_n664_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n348_), .A2(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n642_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n675_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(G57gat), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n766_), .A2(new_n767_), .A3(new_n604_), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT109), .Z(new_n769_));
  NAND2_X1  g568(.A1(new_n614_), .A2(new_n763_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n770_), .B(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n642_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(new_n350_), .A3(new_n585_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n769_), .B1(new_n775_), .B2(new_n767_), .ZN(G1332gat));
  OAI21_X1  g575(.A(G64gat), .B1(new_n766_), .B2(new_n606_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT48), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n774_), .A2(new_n350_), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n606_), .A2(G64gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n778_), .B1(new_n779_), .B2(new_n780_), .ZN(G1333gat));
  OAI21_X1  g580(.A(G71gat), .B1(new_n766_), .B2(new_n416_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT49), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n416_), .A2(G71gat), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n783_), .B1(new_n779_), .B2(new_n784_), .ZN(G1334gat));
  OAI21_X1  g584(.A(G78gat), .B1(new_n766_), .B2(new_n610_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT50), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n610_), .A2(G78gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n779_), .B2(new_n788_), .ZN(G1335gat));
  NOR3_X1   g588(.A1(new_n642_), .A2(new_n348_), .A3(new_n665_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n790_), .B1(new_n715_), .B2(new_n718_), .ZN(new_n791_));
  OAI21_X1  g590(.A(G85gat), .B1(new_n791_), .B2(new_n604_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n772_), .A2(new_n773_), .A3(new_n701_), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n604_), .A2(G85gat), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n792_), .B1(new_n793_), .B2(new_n794_), .ZN(G1336gat));
  OAI21_X1  g594(.A(G92gat), .B1(new_n791_), .B2(new_n606_), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n606_), .A2(G92gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n793_), .B2(new_n797_), .ZN(G1337gat));
  OAI21_X1  g597(.A(G99gat), .B1(new_n791_), .B2(new_n416_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n692_), .A2(new_n218_), .A3(new_n220_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n799_), .B1(new_n793_), .B2(new_n800_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g601(.A(G106gat), .B1(new_n791_), .B2(new_n610_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804_));
  OR2_X1    g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n804_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n793_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n610_), .A2(G106gat), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT110), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT110), .ZN(new_n810_));
  NOR4_X1   g609(.A1(new_n793_), .A2(new_n810_), .A3(G106gat), .A4(new_n610_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n805_), .B(new_n806_), .C1(new_n809_), .C2(new_n811_), .ZN(new_n812_));
  XOR2_X1   g611(.A(KEYINPUT111), .B(KEYINPUT53), .Z(new_n813_));
  XNOR2_X1  g612(.A(new_n812_), .B(new_n813_), .ZN(G1339gat));
  NAND3_X1  g613(.A1(new_n645_), .A2(new_n646_), .A3(new_n649_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n662_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT115), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n646_), .B1(new_n656_), .B2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n819_), .B1(new_n818_), .B2(new_n656_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n817_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n651_), .A2(new_n657_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n661_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n635_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n625_), .A2(new_n827_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n624_), .A2(new_n621_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n829_), .A2(KEYINPUT55), .A3(new_n619_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n620_), .A2(KEYINPUT114), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n828_), .A2(new_n830_), .A3(new_n832_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n829_), .A2(KEYINPUT55), .A3(new_n619_), .A4(new_n831_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n834_), .A2(new_n632_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n833_), .A2(new_n835_), .A3(KEYINPUT56), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(KEYINPUT56), .B1(new_n833_), .B2(new_n835_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n826_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT58), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n321_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT117), .B1(new_n839_), .B2(new_n840_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n833_), .A2(new_n835_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT56), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n836_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n846_), .A2(new_n847_), .A3(KEYINPUT58), .A4(new_n826_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n841_), .A2(new_n842_), .A3(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n824_), .B1(new_n633_), .B2(new_n635_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n665_), .A2(KEYINPUT113), .A3(new_n635_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(new_n763_), .B2(new_n825_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n852_), .A2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n851_), .B1(new_n855_), .B2(new_n846_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n850_), .B1(new_n856_), .B2(new_n674_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n854_), .B(new_n852_), .C1(new_n837_), .C2(new_n838_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n851_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n860_), .A2(KEYINPUT57), .A3(new_n700_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n849_), .A2(new_n857_), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n347_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n764_), .ZN(new_n864_));
  AOI21_X1  g663(.A(KEYINPUT112), .B1(new_n642_), .B2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT112), .ZN(new_n866_));
  AOI211_X1 g665(.A(new_n866_), .B(new_n764_), .C1(new_n640_), .C2(new_n641_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n321_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(KEYINPUT54), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT54), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n870_), .B(new_n321_), .C1(new_n865_), .C2(new_n867_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n863_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT59), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n611_), .A2(new_n604_), .A3(new_n416_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n873_), .A2(new_n874_), .A3(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n875_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT118), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n873_), .A2(new_n878_), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n862_), .A2(new_n347_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(KEYINPUT118), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n877_), .B1(new_n879_), .B2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n876_), .B1(new_n882_), .B2(new_n874_), .ZN(new_n883_));
  OAI21_X1  g682(.A(G113gat), .B1(new_n883_), .B2(new_n763_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n882_), .A2(new_n398_), .A3(new_n665_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1340gat));
  XOR2_X1   g685(.A(KEYINPUT119), .B(G120gat), .Z(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n888_), .B1(new_n883_), .B2(new_n642_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n887_), .B1(new_n642_), .B2(KEYINPUT60), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n882_), .B(new_n890_), .C1(KEYINPUT60), .C2(new_n887_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n891_), .ZN(G1341gat));
  OAI21_X1  g691(.A(G127gat), .B1(new_n883_), .B2(new_n347_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n882_), .A2(new_n388_), .A3(new_n348_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1342gat));
  OAI21_X1  g694(.A(G134gat), .B1(new_n883_), .B2(new_n321_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n882_), .A2(new_n390_), .A3(new_n674_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1343gat));
  NAND2_X1  g697(.A1(new_n879_), .A2(new_n881_), .ZN(new_n899_));
  NOR4_X1   g698(.A1(new_n692_), .A2(new_n610_), .A3(new_n601_), .A4(new_n604_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n899_), .A2(new_n665_), .A3(new_n900_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g701(.A1(new_n899_), .A2(new_n773_), .A3(new_n900_), .ZN(new_n903_));
  XOR2_X1   g702(.A(KEYINPUT120), .B(G148gat), .Z(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1345gat));
  NAND3_X1  g704(.A1(new_n899_), .A2(new_n348_), .A3(new_n900_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT61), .B(G155gat), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n906_), .B(new_n907_), .ZN(G1346gat));
  AND2_X1   g707(.A1(new_n899_), .A2(new_n900_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(new_n674_), .ZN(new_n910_));
  AND2_X1   g709(.A1(new_n714_), .A2(G162gat), .ZN(new_n911_));
  AOI22_X1  g710(.A1(new_n910_), .A2(new_n465_), .B1(new_n909_), .B2(new_n911_), .ZN(G1347gat));
  XOR2_X1   g711(.A(KEYINPUT22), .B(G169gat), .Z(new_n913_));
  NOR2_X1   g712(.A1(new_n763_), .A2(new_n913_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n416_), .A2(new_n606_), .A3(new_n585_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n610_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(KEYINPUT121), .B1(new_n873_), .B2(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT121), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n880_), .A2(new_n919_), .A3(new_n916_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n914_), .B1(new_n918_), .B2(new_n920_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n873_), .A2(new_n665_), .A3(new_n917_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n923_));
  AND3_X1   g722(.A1(new_n922_), .A2(new_n923_), .A3(G169gat), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n923_), .B1(new_n922_), .B2(G169gat), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n921_), .B1(new_n924_), .B2(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(KEYINPUT122), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT122), .ZN(new_n928_));
  OAI211_X1 g727(.A(new_n921_), .B(new_n928_), .C1(new_n924_), .C2(new_n925_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n929_), .ZN(G1348gat));
  AND3_X1   g729(.A1(new_n863_), .A2(KEYINPUT118), .A3(new_n872_), .ZN(new_n931_));
  AOI21_X1  g730(.A(KEYINPUT118), .B1(new_n863_), .B2(new_n872_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n610_), .B1(new_n931_), .B2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(KEYINPUT123), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n935_));
  OAI211_X1 g734(.A(new_n935_), .B(new_n610_), .C1(new_n931_), .C2(new_n932_), .ZN(new_n936_));
  INV_X1    g735(.A(G176gat), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n642_), .A2(new_n937_), .ZN(new_n938_));
  NAND4_X1  g737(.A1(new_n934_), .A2(new_n915_), .A3(new_n936_), .A4(new_n938_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n918_), .A2(new_n920_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n937_), .B1(new_n940_), .B2(new_n642_), .ZN(new_n941_));
  AND2_X1   g740(.A1(new_n939_), .A2(new_n941_), .ZN(G1349gat));
  NAND4_X1  g741(.A1(new_n934_), .A2(new_n348_), .A3(new_n915_), .A4(new_n936_), .ZN(new_n943_));
  INV_X1    g742(.A(new_n940_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n347_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n945_));
  AOI22_X1  g744(.A1(new_n943_), .A2(new_n351_), .B1(new_n944_), .B2(new_n945_), .ZN(G1350gat));
  OAI21_X1  g745(.A(G190gat), .B1(new_n940_), .B2(new_n321_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n674_), .A2(new_n356_), .A3(new_n358_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n940_), .B2(new_n948_), .ZN(G1351gat));
  NOR2_X1   g748(.A1(new_n692_), .A2(new_n596_), .ZN(new_n950_));
  AND2_X1   g749(.A1(new_n950_), .A2(KEYINPUT124), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n950_), .A2(KEYINPUT124), .ZN(new_n952_));
  NOR3_X1   g751(.A1(new_n951_), .A2(new_n952_), .A3(new_n606_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n899_), .A2(new_n665_), .A3(new_n953_), .ZN(new_n954_));
  INV_X1    g753(.A(G197gat), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n954_), .B1(KEYINPUT125), .B2(new_n955_), .ZN(new_n956_));
  XOR2_X1   g755(.A(KEYINPUT125), .B(G197gat), .Z(new_n957_));
  AND2_X1   g756(.A1(new_n954_), .A2(new_n957_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n956_), .A2(new_n958_), .ZN(G1352gat));
  NAND3_X1  g758(.A1(new_n899_), .A2(new_n773_), .A3(new_n953_), .ZN(new_n960_));
  XOR2_X1   g759(.A(KEYINPUT126), .B(G204gat), .Z(new_n961_));
  XNOR2_X1  g760(.A(new_n960_), .B(new_n961_), .ZN(G1353gat));
  NAND3_X1  g761(.A1(new_n899_), .A2(new_n348_), .A3(new_n953_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(KEYINPUT63), .B(G211gat), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n963_), .A2(new_n964_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n966_));
  AOI21_X1  g765(.A(new_n965_), .B1(new_n963_), .B2(new_n966_), .ZN(G1354gat));
  AND2_X1   g766(.A1(new_n899_), .A2(new_n953_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n968_), .A2(new_n674_), .ZN(new_n969_));
  XOR2_X1   g768(.A(KEYINPUT127), .B(G218gat), .Z(new_n970_));
  NOR2_X1   g769(.A1(new_n321_), .A2(new_n970_), .ZN(new_n971_));
  AOI22_X1  g770(.A1(new_n969_), .A2(new_n970_), .B1(new_n968_), .B2(new_n971_), .ZN(G1355gat));
endmodule


