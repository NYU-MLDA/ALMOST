//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n839_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n847_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n853_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_;
  XNOR2_X1  g000(.A(G71gat), .B(G99gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G15gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT80), .B(G43gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G227gat), .A2(G233gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT77), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT77), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n210_), .B1(G169gat), .B2(G176gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT24), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n212_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G183gat), .ZN(new_n218_));
  INV_X1    g017(.A(G190gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT23), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G183gat), .A3(G190gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT26), .B(G190gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT25), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n225_), .A2(KEYINPUT76), .A3(G183gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT76), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT25), .B1(new_n227_), .B2(new_n218_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n224_), .A2(new_n226_), .A3(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n209_), .A2(new_n211_), .A3(new_n215_), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n217_), .A2(new_n223_), .A3(new_n229_), .A4(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n222_), .A2(KEYINPUT79), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT79), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n233_), .A2(new_n221_), .A3(G183gat), .A4(G190gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  AOI22_X1  g034(.A1(new_n235_), .A2(new_n220_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n236_));
  INV_X1    g035(.A(G176gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT22), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(G169gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT78), .ZN(new_n240_));
  INV_X1    g039(.A(G169gat), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n240_), .B1(KEYINPUT22), .B2(new_n241_), .ZN(new_n242_));
  NOR3_X1   g041(.A1(new_n238_), .A2(KEYINPUT78), .A3(G169gat), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n237_), .B(new_n239_), .C1(new_n242_), .C2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(new_n213_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n231_), .B1(new_n236_), .B2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT30), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT81), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n247_), .A2(new_n248_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n207_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n251_), .B1(new_n249_), .B2(new_n207_), .ZN(new_n252_));
  AND2_X1   g051(.A1(G113gat), .A2(G120gat), .ZN(new_n253_));
  NOR2_X1   g052(.A1(G113gat), .A2(G120gat), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT82), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(G113gat), .ZN(new_n256_));
  INV_X1    g055(.A(G120gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT82), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G113gat), .A2(G120gat), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n258_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  AND2_X1   g060(.A1(G127gat), .A2(G134gat), .ZN(new_n262_));
  NOR2_X1   g061(.A1(G127gat), .A2(G134gat), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n255_), .A2(new_n261_), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT84), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT84), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n255_), .A2(new_n261_), .A3(new_n267_), .A4(new_n264_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n255_), .A2(new_n261_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n264_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT83), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n269_), .A2(new_n274_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n266_), .A2(new_n272_), .A3(new_n273_), .A4(new_n268_), .ZN(new_n276_));
  AND2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(KEYINPUT85), .B(KEYINPUT31), .Z(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n252_), .A2(new_n280_), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n251_), .B(new_n279_), .C1(new_n249_), .C2(new_n207_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G78gat), .B(G106gat), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(G141gat), .A2(G148gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT3), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT2), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(G155gat), .ZN(new_n292_));
  INV_X1    g091(.A(G162gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n292_), .A2(new_n293_), .A3(KEYINPUT87), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT87), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n295_), .B1(G155gat), .B2(G162gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n294_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT1), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n297_), .B(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n300_), .A2(new_n294_), .A3(new_n296_), .ZN(new_n301_));
  XOR2_X1   g100(.A(G141gat), .B(G148gat), .Z(new_n302_));
  AOI22_X1  g101(.A1(new_n291_), .A2(new_n298_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT29), .ZN(new_n304_));
  INV_X1    g103(.A(G233gat), .ZN(new_n305_));
  NOR2_X1   g104(.A1(KEYINPUT89), .A2(G228gat), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(KEYINPUT89), .A2(G228gat), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n305_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n303_), .A2(new_n304_), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n310_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n286_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n313_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n315_), .A2(new_n285_), .A3(new_n311_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G22gat), .B(G50gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G197gat), .B(G204gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT90), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT21), .ZN(new_n322_));
  INV_X1    g121(.A(G204gat), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n323_), .A2(G197gat), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT90), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n322_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(G211gat), .A2(G218gat), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT92), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G211gat), .A2(G218gat), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n328_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  AND2_X1   g130(.A1(G211gat), .A2(G218gat), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT92), .B1(new_n332_), .B2(new_n327_), .ZN(new_n333_));
  AOI22_X1  g132(.A1(new_n321_), .A2(new_n326_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(G197gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(G204gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n323_), .A2(G197gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(new_n337_), .A3(new_n322_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT91), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT91), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n320_), .A2(new_n340_), .A3(new_n322_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n334_), .A2(new_n342_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n331_), .A2(new_n333_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n320_), .A2(new_n322_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n343_), .A2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n347_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n318_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n314_), .A2(new_n316_), .A3(new_n352_), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n319_), .A2(new_n351_), .A3(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n351_), .B1(new_n319_), .B2(new_n353_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n284_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G1gat), .B(G29gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(G85gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT0), .B(G57gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n291_), .A2(new_n298_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n301_), .A2(new_n302_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n275_), .A2(new_n276_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n272_), .A2(new_n265_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n303_), .A2(new_n367_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n366_), .A2(KEYINPUT96), .A3(KEYINPUT4), .A4(new_n368_), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n366_), .A2(KEYINPUT4), .A3(new_n368_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT4), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n275_), .A2(new_n365_), .A3(new_n371_), .A4(new_n276_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT96), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n369_), .B1(new_n370_), .B2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G225gat), .A2(G233gat), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n366_), .A2(new_n368_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n379_), .A2(new_n377_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n362_), .B1(new_n378_), .B2(new_n381_), .ZN(new_n382_));
  AOI211_X1 g181(.A(new_n380_), .B(new_n361_), .C1(new_n375_), .C2(new_n377_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT27), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT20), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n219_), .A2(KEYINPUT26), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT26), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(G190gat), .ZN(new_n389_));
  AND2_X1   g188(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n390_));
  NOR2_X1   g189(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n387_), .B(new_n389_), .C1(new_n390_), .C2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n208_), .A2(new_n215_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n213_), .A2(KEYINPUT24), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n395_), .B1(new_n209_), .B2(new_n211_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n235_), .A2(new_n220_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n223_), .B1(G183gat), .B2(G190gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT22), .B(G169gat), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n214_), .B1(new_n400_), .B2(new_n237_), .ZN(new_n401_));
  AOI22_X1  g200(.A1(new_n397_), .A2(new_n398_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n402_));
  AOI22_X1  g201(.A1(new_n334_), .A2(new_n342_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n386_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G226gat), .A2(G233gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT19), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n347_), .A2(new_n246_), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n404_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT20), .B1(new_n347_), .B2(new_n246_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT93), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  OAI211_X1 g211(.A(KEYINPUT93), .B(KEYINPUT20), .C1(new_n347_), .C2(new_n246_), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n402_), .A2(new_n403_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n412_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n409_), .B1(new_n415_), .B2(new_n406_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G8gat), .B(G36gat), .ZN(new_n417_));
  XOR2_X1   g216(.A(new_n417_), .B(KEYINPUT95), .Z(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT94), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n417_), .B(KEYINPUT95), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT94), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  XOR2_X1   g221(.A(G64gat), .B(G92gat), .Z(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT18), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n419_), .A2(new_n422_), .A3(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n424_), .B1(new_n419_), .B2(new_n422_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n416_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n427_), .ZN(new_n429_));
  AOI211_X1 g228(.A(new_n409_), .B(new_n429_), .C1(new_n415_), .C2(new_n406_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n385_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n416_), .A2(new_n427_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT99), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n408_), .B1(new_n404_), .B2(new_n433_), .ZN(new_n434_));
  AOI211_X1 g233(.A(KEYINPUT99), .B(new_n386_), .C1(new_n402_), .C2(new_n403_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n406_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n412_), .A2(new_n407_), .A3(new_n413_), .A4(new_n414_), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n432_), .B(KEYINPUT27), .C1(new_n427_), .C2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n431_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n357_), .A2(new_n384_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n384_), .A2(new_n356_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n443_), .A2(new_n440_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT32), .ZN(new_n445_));
  NOR3_X1   g244(.A1(new_n425_), .A2(new_n426_), .A3(new_n445_), .ZN(new_n446_));
  AOI211_X1 g245(.A(new_n446_), .B(new_n409_), .C1(new_n415_), .C2(new_n406_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n446_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n448_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n450_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT100), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n378_), .A2(new_n381_), .A3(new_n362_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT33), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n361_), .B1(new_n379_), .B2(new_n376_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT97), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT98), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n366_), .A2(KEYINPUT4), .A3(new_n368_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(new_n373_), .A3(new_n372_), .ZN(new_n462_));
  AOI211_X1 g261(.A(new_n460_), .B(new_n377_), .C1(new_n462_), .C2(new_n369_), .ZN(new_n463_));
  AOI21_X1  g262(.A(KEYINPUT98), .B1(new_n375_), .B2(new_n376_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n459_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n428_), .A2(new_n430_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n378_), .A2(KEYINPUT33), .A3(new_n381_), .A4(new_n362_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n456_), .A2(new_n465_), .A3(new_n466_), .A4(new_n467_), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n450_), .B(KEYINPUT100), .C1(new_n382_), .C2(new_n383_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n453_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n356_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n444_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n284_), .A2(KEYINPUT86), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT86), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n283_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n442_), .B1(new_n472_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT7), .ZN(new_n478_));
  INV_X1    g277(.A(G99gat), .ZN(new_n479_));
  INV_X1    g278(.A(G106gat), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G99gat), .A2(G106gat), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT6), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n481_), .A2(new_n484_), .A3(new_n485_), .A4(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G85gat), .B(G92gat), .Z(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT65), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT8), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT10), .B(G99gat), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n493_), .A2(G106gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n488_), .A2(KEYINPUT9), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n484_), .A2(new_n485_), .ZN(new_n496_));
  INV_X1    g295(.A(G92gat), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n497_), .A2(KEYINPUT9), .ZN(new_n498_));
  OR2_X1    g297(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n498_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .A4(new_n501_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n492_), .A2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT65), .B1(new_n487_), .B2(new_n488_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n487_), .A2(KEYINPUT65), .A3(new_n488_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(KEYINPUT8), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n503_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G29gat), .B(G36gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G43gat), .B(G50gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT15), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n508_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n506_), .A2(KEYINPUT8), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n514_), .A2(new_n504_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n492_), .A2(new_n502_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(new_n511_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G232gat), .A2(G233gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT34), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n520_), .A2(KEYINPUT35), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(KEYINPUT35), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n513_), .A2(new_n518_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n513_), .A2(KEYINPUT67), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT67), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n508_), .A2(new_n526_), .A3(new_n512_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(new_n527_), .A3(new_n518_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n524_), .B1(new_n528_), .B2(new_n521_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G190gat), .B(G218gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(new_n293_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT68), .B(G134gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n531_), .B(new_n532_), .Z(new_n533_));
  NAND2_X1  g332(.A1(KEYINPUT69), .A2(KEYINPUT36), .ZN(new_n534_));
  OR2_X1    g333(.A1(KEYINPUT69), .A2(KEYINPUT36), .ZN(new_n535_));
  AND3_X1   g334(.A1(new_n533_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n529_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT70), .B(KEYINPUT36), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n533_), .B(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n537_), .B1(new_n529_), .B2(new_n539_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n477_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT66), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT12), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G57gat), .B(G64gat), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n545_), .A2(KEYINPUT11), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(KEYINPUT11), .ZN(new_n547_));
  XOR2_X1   g346(.A(G71gat), .B(G78gat), .Z(new_n548_));
  NAND3_X1  g347(.A1(new_n546_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n547_), .A2(new_n548_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n544_), .B1(new_n508_), .B2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n503_), .A2(new_n507_), .A3(new_n551_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n542_), .A2(new_n543_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G230gat), .A2(G233gat), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n508_), .A2(new_n552_), .A3(new_n544_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n557_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n552_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n554_), .A2(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n560_), .B1(new_n558_), .B2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G120gat), .B(G148gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(new_n323_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT5), .B(G176gat), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n565_), .B(new_n566_), .Z(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n563_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT13), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n563_), .A2(new_n568_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n563_), .A2(new_n568_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n573_), .A2(KEYINPUT13), .A3(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n571_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(G1gat), .ZN(new_n578_));
  INV_X1    g377(.A(G8gat), .ZN(new_n579_));
  OAI21_X1  g378(.A(KEYINPUT14), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT72), .B(G15gat), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(G22gat), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n580_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(G1gat), .B(G8gat), .Z(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n581_), .A2(G22gat), .ZN(new_n587_));
  OR3_X1    g386(.A1(new_n584_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n586_), .B1(new_n584_), .B2(new_n587_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(new_n512_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G229gat), .A2(G233gat), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n588_), .A2(new_n511_), .A3(new_n589_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n591_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n590_), .B(new_n511_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n594_), .B1(new_n595_), .B2(new_n592_), .ZN(new_n596_));
  XOR2_X1   g395(.A(G169gat), .B(G197gat), .Z(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT74), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G113gat), .B(G141gat), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n598_), .B(new_n599_), .Z(new_n600_));
  XNOR2_X1  g399(.A(new_n596_), .B(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n577_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G231gat), .A2(G233gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT73), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n590_), .B(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(new_n552_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G127gat), .B(G155gat), .ZN(new_n608_));
  INV_X1    g407(.A(G211gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(KEYINPUT16), .B(G183gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n612_), .A2(KEYINPUT17), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(KEYINPUT17), .ZN(new_n614_));
  OR3_X1    g413(.A1(new_n607_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n607_), .A2(new_n613_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n603_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n541_), .A2(new_n618_), .ZN(new_n619_));
  OAI21_X1  g418(.A(G1gat), .B1(new_n619_), .B2(new_n384_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT102), .Z(new_n621_));
  XNOR2_X1  g420(.A(new_n601_), .B(KEYINPUT75), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n576_), .A2(new_n622_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n477_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT37), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT71), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n625_), .B1(new_n537_), .B2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n540_), .ZN(new_n628_));
  OAI221_X1 g427(.A(new_n537_), .B1(new_n626_), .B2(new_n625_), .C1(new_n529_), .C2(new_n539_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n631_), .A2(new_n617_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n624_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n384_), .B(KEYINPUT101), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n634_), .A2(new_n578_), .A3(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(KEYINPUT103), .A2(KEYINPUT38), .ZN(new_n638_));
  AND2_X1   g437(.A1(KEYINPUT103), .A2(KEYINPUT38), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n637_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n621_), .B(new_n640_), .C1(new_n638_), .C2(new_n637_), .ZN(G1324gat));
  NAND3_X1  g440(.A1(new_n634_), .A2(new_n579_), .A3(new_n440_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT105), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n618_), .A2(new_n477_), .A3(new_n540_), .A4(new_n440_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(G8gat), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n645_), .A2(KEYINPUT104), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(KEYINPUT104), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n643_), .B(KEYINPUT39), .C1(new_n646_), .C2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n645_), .B(KEYINPUT104), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n648_), .B1(KEYINPUT39), .B2(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n643_), .B1(new_n649_), .B2(KEYINPUT39), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n642_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT40), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  OAI211_X1 g453(.A(KEYINPUT40), .B(new_n642_), .C1(new_n650_), .C2(new_n651_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1325gat));
  INV_X1    g455(.A(new_n476_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G15gat), .B1(new_n619_), .B2(new_n657_), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n658_), .A2(KEYINPUT41), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(KEYINPUT41), .ZN(new_n660_));
  OR3_X1    g459(.A1(new_n633_), .A2(G15gat), .A3(new_n657_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n659_), .A2(new_n660_), .A3(new_n661_), .ZN(G1326gat));
  OAI21_X1  g461(.A(G22gat), .B1(new_n619_), .B2(new_n471_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT42), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n634_), .A2(new_n583_), .A3(new_n356_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1327gat));
  INV_X1    g465(.A(new_n617_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n603_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT43), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n477_), .A2(new_n669_), .A3(new_n631_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n669_), .B1(new_n477_), .B2(new_n631_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n668_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  OAI211_X1 g473(.A(KEYINPUT44), .B(new_n668_), .C1(new_n670_), .C2(new_n671_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G29gat), .B1(new_n676_), .B2(new_n635_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n667_), .A2(new_n540_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n624_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT106), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n624_), .A2(KEYINPUT106), .A3(new_n678_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n384_), .A2(G29gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n677_), .B1(new_n683_), .B2(new_n684_), .ZN(G1328gat));
  NOR2_X1   g484(.A1(new_n441_), .A2(G36gat), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n681_), .A2(new_n682_), .A3(new_n686_), .ZN(new_n687_));
  XOR2_X1   g486(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n674_), .A2(new_n440_), .A3(new_n675_), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n690_), .A2(KEYINPUT107), .A3(G36gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT107), .B1(new_n690_), .B2(G36gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n689_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  OAI221_X1 g494(.A(new_n689_), .B1(KEYINPUT109), .B2(KEYINPUT46), .C1(new_n691_), .C2(new_n692_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1329gat));
  OAI21_X1  g496(.A(G43gat), .B1(new_n676_), .B2(new_n284_), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n657_), .A2(G43gat), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n698_), .B1(new_n683_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT47), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n700_), .B(new_n701_), .ZN(G1330gat));
  OAI21_X1  g501(.A(G50gat), .B1(new_n676_), .B2(new_n471_), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n471_), .A2(G50gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n683_), .B2(new_n704_), .ZN(G1331gat));
  AND3_X1   g504(.A1(new_n576_), .A2(new_n667_), .A3(new_n622_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n541_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(G57gat), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n707_), .A2(new_n708_), .A3(new_n384_), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n477_), .A2(new_n576_), .A3(new_n601_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(new_n632_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n635_), .B1(new_n711_), .B2(KEYINPUT110), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n712_), .B1(KEYINPUT110), .B2(new_n711_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n709_), .B1(new_n713_), .B2(new_n708_), .ZN(G1332gat));
  OAI21_X1  g513(.A(G64gat), .B1(new_n707_), .B2(new_n441_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n715_), .A2(KEYINPUT48), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n715_), .A2(KEYINPUT48), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n441_), .A2(G64gat), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT111), .ZN(new_n719_));
  OAI22_X1  g518(.A1(new_n716_), .A2(new_n717_), .B1(new_n711_), .B2(new_n719_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT112), .Z(G1333gat));
  OAI21_X1  g520(.A(G71gat), .B1(new_n707_), .B2(new_n657_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT49), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n657_), .A2(G71gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n723_), .B1(new_n711_), .B2(new_n724_), .ZN(G1334gat));
  OAI21_X1  g524(.A(G78gat), .B1(new_n707_), .B2(new_n471_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT50), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n471_), .A2(G78gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(new_n711_), .B2(new_n728_), .ZN(G1335gat));
  NAND2_X1  g528(.A1(new_n710_), .A2(new_n678_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(G85gat), .B1(new_n731_), .B2(new_n636_), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n670_), .A2(new_n671_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n577_), .A2(new_n667_), .A3(new_n602_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT113), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n499_), .B(new_n500_), .C1(new_n382_), .C2(new_n383_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT114), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n732_), .B1(new_n736_), .B2(new_n738_), .ZN(G1336gat));
  OAI21_X1  g538(.A(new_n497_), .B1(new_n730_), .B2(new_n441_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT115), .Z(new_n741_));
  NOR2_X1   g540(.A1(new_n441_), .A2(new_n497_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n736_), .B2(new_n742_), .ZN(G1337gat));
  OAI21_X1  g542(.A(G99gat), .B1(new_n735_), .B2(new_n657_), .ZN(new_n744_));
  OR3_X1    g543(.A1(new_n730_), .A2(new_n493_), .A3(new_n284_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g546(.A1(new_n731_), .A2(new_n480_), .A3(new_n356_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n733_), .A2(new_n356_), .A3(new_n734_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n749_), .A2(new_n750_), .A3(G106gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n749_), .B2(G106gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n753_), .B(new_n755_), .ZN(G1339gat));
  NAND3_X1  g555(.A1(new_n632_), .A2(new_n577_), .A3(new_n622_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT54), .ZN(new_n758_));
  AOI22_X1  g557(.A1(new_n517_), .A2(new_n551_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n544_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n561_), .A2(new_n760_), .ZN(new_n761_));
  AND4_X1   g560(.A1(new_n558_), .A2(new_n759_), .A3(new_n559_), .A4(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n759_), .A2(new_n559_), .A3(new_n761_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n558_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n762_), .B1(KEYINPUT55), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT55), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n763_), .A2(new_n767_), .A3(new_n764_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n568_), .B1(new_n766_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT56), .ZN(new_n770_));
  INV_X1    g569(.A(new_n600_), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n596_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n592_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n591_), .A2(new_n773_), .A3(new_n593_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n771_), .B(new_n774_), .C1(new_n595_), .C2(new_n773_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n772_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT56), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n777_), .B(new_n568_), .C1(new_n766_), .C2(new_n768_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n770_), .A2(new_n573_), .A3(new_n776_), .A4(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT58), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n630_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n572_), .B1(new_n769_), .B2(KEYINPUT56), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n782_), .A2(KEYINPUT58), .A3(new_n776_), .A4(new_n778_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n540_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n601_), .B1(new_n769_), .B2(KEYINPUT117), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n558_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n560_), .B1(new_n787_), .B2(new_n767_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n768_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n790_), .A2(new_n791_), .A3(new_n777_), .A4(new_n568_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n782_), .A2(new_n786_), .A3(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n569_), .A2(new_n776_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n785_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n784_), .B1(new_n795_), .B2(KEYINPUT57), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT57), .ZN(new_n797_));
  AOI211_X1 g596(.A(new_n797_), .B(new_n785_), .C1(new_n793_), .C2(new_n794_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n617_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n758_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n357_), .A2(new_n441_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n801_), .A2(KEYINPUT59), .A3(new_n635_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n622_), .A2(new_n256_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n801_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n806_), .B1(new_n781_), .B2(new_n783_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n567_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n573_), .B1(new_n808_), .B2(new_n777_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n778_), .A2(new_n776_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n780_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  AND4_X1   g610(.A1(new_n806_), .A2(new_n811_), .A3(new_n631_), .A4(new_n783_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n807_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n793_), .A2(new_n794_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT57), .B1(new_n814_), .B2(new_n540_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n815_), .A2(new_n798_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n667_), .B1(new_n813_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n757_), .B(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n805_), .B(new_n636_), .C1(new_n817_), .C2(new_n819_), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n820_), .A2(KEYINPUT119), .A3(KEYINPUT59), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT119), .B1(new_n820_), .B2(KEYINPUT59), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n803_), .B(new_n804_), .C1(new_n821_), .C2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n256_), .B1(new_n820_), .B2(new_n601_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT120), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n823_), .A2(KEYINPUT120), .A3(new_n824_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(G1340gat));
  INV_X1    g628(.A(new_n820_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT60), .ZN(new_n831_));
  XOR2_X1   g630(.A(KEYINPUT121), .B(G120gat), .Z(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n577_), .B2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n577_), .B1(new_n830_), .B2(new_n833_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n834_), .B(new_n803_), .C1(new_n822_), .C2(new_n821_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n832_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n830_), .A2(new_n831_), .A3(new_n833_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(G1341gat));
  AOI21_X1  g637(.A(G127gat), .B1(new_n830_), .B2(new_n667_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n821_), .A2(new_n822_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n840_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n667_), .A2(G127gat), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n839_), .B1(new_n841_), .B2(new_n842_), .ZN(G1342gat));
  AOI21_X1  g642(.A(G134gat), .B1(new_n830_), .B2(new_n785_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n631_), .A2(G134gat), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n844_), .B1(new_n841_), .B2(new_n845_), .ZN(G1343gat));
  OR2_X1    g645(.A1(new_n817_), .A2(new_n819_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n476_), .A2(new_n471_), .A3(new_n440_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(new_n636_), .A3(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n849_), .A2(new_n601_), .ZN(new_n850_));
  XOR2_X1   g649(.A(new_n850_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g650(.A1(new_n849_), .A2(new_n577_), .ZN(new_n852_));
  XOR2_X1   g651(.A(KEYINPUT122), .B(G148gat), .Z(new_n853_));
  XNOR2_X1  g652(.A(new_n852_), .B(new_n853_), .ZN(G1345gat));
  NOR2_X1   g653(.A1(new_n849_), .A2(new_n617_), .ZN(new_n855_));
  XOR2_X1   g654(.A(KEYINPUT61), .B(G155gat), .Z(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1346gat));
  AND4_X1   g656(.A1(new_n785_), .A2(new_n847_), .A3(new_n636_), .A4(new_n848_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n631_), .A2(G162gat), .ZN(new_n859_));
  OAI22_X1  g658(.A1(new_n858_), .A2(G162gat), .B1(new_n849_), .B2(new_n859_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(KEYINPUT123), .ZN(G1347gat));
  AOI21_X1  g660(.A(new_n356_), .B1(new_n758_), .B2(new_n799_), .ZN(new_n862_));
  NOR3_X1   g661(.A1(new_n657_), .A2(new_n441_), .A3(new_n636_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n602_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(KEYINPUT124), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n241_), .B1(new_n862_), .B2(new_n865_), .ZN(new_n866_));
  XOR2_X1   g665(.A(new_n866_), .B(KEYINPUT62), .Z(new_n867_));
  NAND2_X1  g666(.A1(new_n862_), .A2(new_n863_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n869_), .A2(new_n400_), .A3(new_n602_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n867_), .A2(new_n870_), .ZN(G1348gat));
  AOI21_X1  g670(.A(G176gat), .B1(new_n869_), .B2(new_n576_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n817_), .A2(new_n819_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n356_), .ZN(new_n874_));
  AND3_X1   g673(.A1(new_n863_), .A2(G176gat), .A3(new_n576_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n872_), .B1(new_n874_), .B2(new_n875_), .ZN(G1349gat));
  NOR2_X1   g675(.A1(new_n390_), .A2(new_n391_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n869_), .A2(new_n877_), .A3(new_n667_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT125), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n878_), .A2(new_n879_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n863_), .A2(new_n667_), .ZN(new_n882_));
  AOI21_X1  g681(.A(G183gat), .B1(new_n874_), .B2(new_n882_), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n880_), .A2(new_n881_), .A3(new_n883_), .ZN(G1350gat));
  OAI21_X1  g683(.A(G190gat), .B1(new_n868_), .B2(new_n630_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n785_), .A2(new_n224_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n868_), .B2(new_n886_), .ZN(G1351gat));
  NOR4_X1   g686(.A1(new_n873_), .A2(new_n443_), .A3(new_n441_), .A4(new_n476_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n602_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n576_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g691(.A(KEYINPUT63), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n667_), .B1(new_n893_), .B2(new_n609_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(KEYINPUT126), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n888_), .A2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n893_), .A2(new_n609_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n896_), .B(new_n897_), .ZN(G1354gat));
  AND3_X1   g697(.A1(new_n888_), .A2(G218gat), .A3(new_n631_), .ZN(new_n899_));
  AOI21_X1  g698(.A(KEYINPUT127), .B1(new_n888_), .B2(new_n785_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n900_), .A2(G218gat), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n888_), .A2(KEYINPUT127), .A3(new_n785_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n899_), .B1(new_n901_), .B2(new_n902_), .ZN(G1355gat));
endmodule


