//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n898_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n923_,
    new_n924_, new_n926_, new_n927_, new_n928_, new_n930_, new_n931_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_, new_n950_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT74), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G232gat), .A2(G233gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT34), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT70), .B(KEYINPUT35), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n203_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G43gat), .B(G50gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G36gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G29gat), .ZN(new_n212_));
  INV_X1    g011(.A(G29gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(G36gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(new_n214_), .A3(KEYINPUT71), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(KEYINPUT71), .B1(new_n212_), .B2(new_n214_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n210_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n212_), .A2(new_n214_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT71), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(new_n215_), .A3(new_n209_), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n218_), .A2(new_n222_), .A3(KEYINPUT15), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT15), .B1(new_n218_), .B2(new_n222_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G99gat), .A2(G106gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT6), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT10), .B(G99gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G106gat), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n230_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n235_));
  INV_X1    g034(.A(G85gat), .ZN(new_n236_));
  OR2_X1    g035(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n236_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n235_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n234_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT8), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NOR3_X1   g045(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n228_), .A2(KEYINPUT65), .A3(new_n229_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n250_));
  AND3_X1   g049(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n251_));
  AOI21_X1  g050(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n250_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n248_), .A2(new_n249_), .A3(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(G85gat), .B(G92gat), .Z(new_n255_));
  AOI21_X1  g054(.A(new_n244_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n244_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n230_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n257_), .B1(new_n258_), .B2(new_n248_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n243_), .B1(new_n256_), .B2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n208_), .B1(new_n225_), .B2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n218_), .A2(new_n222_), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n262_), .B(new_n243_), .C1(new_n256_), .C2(new_n259_), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n263_), .A2(KEYINPUT72), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n263_), .A2(KEYINPUT72), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n261_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n205_), .A2(new_n207_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n261_), .B(new_n267_), .C1(new_n264_), .C2(new_n265_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n269_), .A2(KEYINPUT73), .A3(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G190gat), .B(G218gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G134gat), .B(G162gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n274_), .A2(KEYINPUT36), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n271_), .A2(new_n276_), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n269_), .A2(KEYINPUT73), .A3(new_n270_), .A4(new_n275_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n274_), .A2(KEYINPUT36), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n280_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n202_), .B1(new_n279_), .B2(new_n282_), .ZN(new_n283_));
  AOI211_X1 g082(.A(KEYINPUT37), .B(new_n281_), .C1(new_n277_), .C2(new_n278_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  AND2_X1   g084(.A1(G230gat), .A2(G233gat), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n234_), .A2(new_n242_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n254_), .A2(new_n255_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT8), .ZN(new_n289_));
  INV_X1    g088(.A(new_n259_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n287_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT11), .ZN(new_n292_));
  NAND2_X1  g091(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n295_));
  NOR3_X1   g094(.A1(new_n294_), .A2(new_n295_), .A3(G78gat), .ZN(new_n296_));
  INV_X1    g095(.A(G78gat), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT66), .ZN(new_n298_));
  INV_X1    g097(.A(G71gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n297_), .B1(new_n300_), .B2(new_n293_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n292_), .B1(new_n296_), .B2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G57gat), .B(G64gat), .ZN(new_n303_));
  OAI21_X1  g102(.A(G78gat), .B1(new_n294_), .B2(new_n295_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n300_), .A2(new_n297_), .A3(new_n293_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(new_n305_), .A3(KEYINPUT11), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n302_), .A2(new_n303_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n303_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n308_), .A2(new_n304_), .A3(new_n305_), .A4(KEYINPUT11), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n286_), .B1(new_n291_), .B2(new_n310_), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n307_), .A2(new_n309_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT12), .ZN(new_n313_));
  AND3_X1   g112(.A1(new_n260_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n313_), .B1(new_n260_), .B2(new_n312_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n311_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n291_), .A2(new_n310_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n260_), .A2(new_n312_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n286_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G176gat), .B(G204gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT69), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G120gat), .B(G148gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT67), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n320_), .B(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n329_), .B(KEYINPUT13), .Z(new_n330_));
  NAND2_X1  g129(.A1(G231gat), .A2(G233gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n310_), .B(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G1gat), .B(G8gat), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G15gat), .B(G22gat), .ZN(new_n335_));
  INV_X1    g134(.A(G8gat), .ZN(new_n336_));
  INV_X1    g135(.A(G1gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT75), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT75), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(G1gat), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n336_), .B1(new_n338_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT14), .ZN(new_n342_));
  OAI211_X1 g141(.A(KEYINPUT76), .B(new_n335_), .C1(new_n341_), .C2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT75), .B(G1gat), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT14), .B1(new_n345_), .B2(new_n336_), .ZN(new_n346_));
  AOI21_X1  g145(.A(KEYINPUT76), .B1(new_n346_), .B2(new_n335_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n334_), .B1(new_n344_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n341_), .A2(new_n342_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n335_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n349_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n352_), .A2(new_n343_), .A3(new_n333_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n348_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n332_), .B(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G127gat), .B(G155gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT16), .ZN(new_n357_));
  XOR2_X1   g156(.A(G183gat), .B(G211gat), .Z(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NOR3_X1   g159(.A1(new_n355_), .A2(KEYINPUT17), .A3(new_n360_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n355_), .A2(KEYINPUT77), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(KEYINPUT17), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n362_), .A2(new_n364_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n361_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n285_), .A2(new_n330_), .A3(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT101), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT2), .ZN(new_n372_));
  INV_X1    g171(.A(G141gat), .ZN(new_n373_));
  INV_X1    g172(.A(G148gat), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n372_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(G141gat), .A2(G148gat), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT3), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n375_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT88), .B1(new_n376_), .B2(new_n377_), .ZN(new_n381_));
  OR3_X1    g180(.A1(new_n376_), .A2(KEYINPUT88), .A3(new_n377_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n380_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(G155gat), .A2(G162gat), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT87), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G155gat), .A2(G162gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n383_), .A2(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n373_), .A2(new_n374_), .ZN(new_n390_));
  XOR2_X1   g189(.A(new_n387_), .B(KEYINPUT1), .Z(new_n391_));
  AOI211_X1 g190(.A(new_n376_), .B(new_n390_), .C1(new_n391_), .C2(new_n386_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n389_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  XOR2_X1   g193(.A(G127gat), .B(G134gat), .Z(new_n395_));
  XOR2_X1   g194(.A(G113gat), .B(G120gat), .Z(new_n396_));
  XOR2_X1   g195(.A(new_n395_), .B(new_n396_), .Z(new_n397_));
  NAND2_X1  g196(.A1(new_n394_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n397_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n393_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n398_), .A2(KEYINPUT4), .A3(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G225gat), .A2(G233gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT97), .ZN(new_n403_));
  OR3_X1    g202(.A1(new_n393_), .A2(KEYINPUT4), .A3(new_n399_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n401_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT98), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G1gat), .B(G29gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(G85gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT0), .B(G57gat), .ZN(new_n410_));
  XOR2_X1   g209(.A(new_n409_), .B(new_n410_), .Z(new_n411_));
  NAND4_X1  g210(.A1(new_n401_), .A2(KEYINPUT98), .A3(new_n403_), .A4(new_n404_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n398_), .A2(new_n400_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n413_), .A2(new_n403_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n407_), .A2(new_n411_), .A3(new_n412_), .A4(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT33), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n414_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT33), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n418_), .A2(new_n419_), .A3(new_n411_), .A4(new_n412_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n417_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G226gat), .A2(G233gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT19), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT91), .B(G204gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(G197gat), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n425_), .B1(G197gat), .B2(G204gat), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT21), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G211gat), .B(G218gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(G204gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(G197gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT90), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT92), .ZN(new_n434_));
  INV_X1    g233(.A(G197gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n424_), .A2(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n433_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n437_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n430_), .B1(new_n438_), .B2(KEYINPUT21), .ZN(new_n439_));
  NOR3_X1   g238(.A1(new_n426_), .A2(new_n427_), .A3(new_n429_), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(G183gat), .ZN(new_n442_));
  INV_X1    g241(.A(G190gat), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT23), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT81), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT23), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(G183gat), .A3(G190gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G169gat), .A2(G176gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT24), .ZN(new_n451_));
  INV_X1    g250(.A(G169gat), .ZN(new_n452_));
  INV_X1    g251(.A(G176gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  MUX2_X1   g253(.A(KEYINPUT24), .B(new_n451_), .S(new_n454_), .Z(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT26), .B(G190gat), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT25), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT80), .B1(new_n457_), .B2(G183gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT25), .B(G183gat), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n456_), .B(new_n458_), .C1(new_n459_), .C2(KEYINPUT80), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n449_), .A2(new_n455_), .A3(new_n460_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n444_), .A2(new_n448_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(G183gat), .A2(G190gat), .ZN(new_n463_));
  XOR2_X1   g262(.A(KEYINPUT83), .B(G176gat), .Z(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT82), .B1(new_n452_), .B2(KEYINPUT22), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT22), .B(G169gat), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n467_), .A2(KEYINPUT82), .ZN(new_n468_));
  OAI221_X1 g267(.A(new_n450_), .B1(new_n462_), .B2(new_n463_), .C1(new_n466_), .C2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n461_), .A2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT20), .B1(new_n441_), .B2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n462_), .B1(new_n459_), .B2(new_n456_), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n472_), .A2(new_n455_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT95), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n467_), .B(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(new_n464_), .ZN(new_n476_));
  XOR2_X1   g275(.A(new_n450_), .B(KEYINPUT94), .Z(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT96), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n476_), .A2(KEYINPUT96), .A3(new_n477_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n449_), .B1(G183gat), .B2(G190gat), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n473_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n439_), .A2(new_n440_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n423_), .B1(new_n471_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n470_), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT20), .B1(new_n485_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n423_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n484_), .A2(new_n485_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G8gat), .B(G36gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT18), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G64gat), .B(G92gat), .ZN(new_n496_));
  XOR2_X1   g295(.A(new_n495_), .B(new_n496_), .Z(new_n497_));
  NAND3_X1  g296(.A1(new_n487_), .A2(new_n493_), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n487_), .A2(new_n493_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n497_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n403_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n401_), .A2(new_n502_), .A3(new_n404_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n411_), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n503_), .B(new_n504_), .C1(new_n413_), .C2(new_n502_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n421_), .A2(new_n498_), .A3(new_n501_), .A4(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n497_), .A2(KEYINPUT32), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n484_), .A2(new_n485_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n423_), .B1(new_n508_), .B2(new_n489_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT20), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n510_), .B1(new_n485_), .B2(new_n488_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n511_), .B(new_n491_), .C1(new_n484_), .C2(new_n485_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n507_), .B1(new_n509_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT99), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  AOI211_X1 g314(.A(KEYINPUT99), .B(new_n507_), .C1(new_n509_), .C2(new_n512_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n507_), .ZN(new_n517_));
  OAI22_X1  g316(.A1(new_n515_), .A2(new_n516_), .B1(new_n499_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT100), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n416_), .A2(new_n519_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n418_), .A2(KEYINPUT100), .A3(new_n411_), .A4(new_n412_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n407_), .A2(new_n412_), .A3(new_n415_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(new_n504_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n520_), .A2(new_n521_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n506_), .B1(new_n518_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT29), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n393_), .A2(new_n527_), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n528_), .A2(KEYINPUT89), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(KEYINPUT89), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G22gat), .B(G50gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT28), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n531_), .B(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G78gat), .B(G106gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G228gat), .A2(G233gat), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n393_), .A2(new_n527_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n536_), .B1(new_n441_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n536_), .ZN(new_n540_));
  NOR3_X1   g339(.A1(new_n485_), .A2(new_n540_), .A3(new_n537_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n535_), .B1(new_n539_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n541_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n540_), .B1(new_n485_), .B2(new_n537_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n535_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n534_), .A2(new_n542_), .A3(KEYINPUT93), .A4(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT93), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n542_), .A2(new_n549_), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n550_), .A2(new_n534_), .B1(new_n542_), .B2(new_n546_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n548_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G227gat), .A2(G233gat), .ZN(new_n553_));
  INV_X1    g352(.A(G15gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(G71gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT84), .B(G43gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(G99gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n556_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT85), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT30), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n470_), .B(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT86), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n470_), .B(KEYINPUT30), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT85), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n565_), .A2(new_n566_), .A3(new_n559_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n563_), .A2(new_n564_), .A3(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT31), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT31), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n563_), .A2(new_n567_), .A3(new_n564_), .A4(new_n570_), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n569_), .A2(new_n397_), .A3(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n397_), .B1(new_n569_), .B2(new_n571_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n552_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n526_), .A2(new_n575_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n568_), .A2(KEYINPUT31), .ZN(new_n577_));
  INV_X1    g376(.A(new_n571_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n399_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n569_), .A2(new_n397_), .A3(new_n571_), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n579_), .B(new_n580_), .C1(new_n548_), .C2(new_n551_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n550_), .A2(new_n534_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n546_), .A2(new_n542_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n584_), .B(new_n547_), .C1(new_n572_), .C2(new_n573_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n581_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n498_), .A2(KEYINPUT27), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n497_), .B1(new_n509_), .B2(new_n512_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(KEYINPUT27), .B1(new_n501_), .B2(new_n498_), .ZN(new_n590_));
  NOR3_X1   g389(.A1(new_n589_), .A2(new_n590_), .A3(new_n524_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n586_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n576_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G113gat), .B(G141gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G169gat), .B(G197gat), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n594_), .B(new_n595_), .Z(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n225_), .A2(new_n353_), .A3(new_n348_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n344_), .A2(new_n347_), .A3(new_n334_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n333_), .B1(new_n352_), .B2(new_n343_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n262_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G229gat), .A2(G233gat), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n598_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT78), .ZN(new_n605_));
  INV_X1    g404(.A(new_n262_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n348_), .A2(new_n353_), .A3(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n606_), .B1(new_n348_), .B2(new_n353_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n605_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n348_), .A2(new_n353_), .A3(new_n606_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n601_), .A2(KEYINPUT78), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n602_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n604_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n597_), .B1(new_n614_), .B2(KEYINPUT79), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT79), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n602_), .B1(new_n609_), .B2(new_n611_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n616_), .B(new_n596_), .C1(new_n617_), .C2(new_n604_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n615_), .A2(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n371_), .B1(new_n593_), .B2(new_n619_), .ZN(new_n620_));
  AOI22_X1  g419(.A1(new_n526_), .A2(new_n575_), .B1(new_n586_), .B2(new_n591_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n619_), .ZN(new_n622_));
  NOR3_X1   g421(.A1(new_n621_), .A2(KEYINPUT101), .A3(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n370_), .B1(new_n620_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT102), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  OAI211_X1 g425(.A(KEYINPUT102), .B(new_n370_), .C1(new_n620_), .C2(new_n623_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n626_), .A2(new_n524_), .A3(new_n345_), .A4(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT38), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n629_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT103), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n279_), .A2(new_n282_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n632_), .B1(new_n621_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n633_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n593_), .A2(KEYINPUT103), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n330_), .A2(new_n619_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n638_), .A2(new_n367_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n640_), .A2(new_n524_), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n630_), .B(new_n631_), .C1(new_n337_), .C2(new_n641_), .ZN(G1324gat));
  INV_X1    g441(.A(new_n589_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n590_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n626_), .A2(new_n336_), .A3(new_n645_), .A4(new_n627_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n637_), .A2(new_n645_), .A3(new_n639_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n647_), .A2(G8gat), .A3(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n647_), .B2(G8gat), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n646_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT40), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OAI211_X1 g452(.A(new_n646_), .B(KEYINPUT40), .C1(new_n649_), .C2(new_n650_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1325gat));
  NAND4_X1  g454(.A1(new_n626_), .A2(new_n554_), .A3(new_n574_), .A4(new_n627_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n640_), .A2(new_n574_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n657_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT41), .B1(new_n657_), .B2(G15gat), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n656_), .B1(new_n658_), .B2(new_n659_), .ZN(G1326gat));
  INV_X1    g459(.A(G22gat), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n626_), .A2(new_n661_), .A3(new_n552_), .A4(new_n627_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT42), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n640_), .A2(new_n552_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n664_), .B2(G22gat), .ZN(new_n665_));
  AOI211_X1 g464(.A(KEYINPUT42), .B(new_n661_), .C1(new_n640_), .C2(new_n552_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n662_), .B1(new_n665_), .B2(new_n666_), .ZN(G1327gat));
  NAND3_X1  g466(.A1(new_n330_), .A2(new_n367_), .A3(new_n633_), .ZN(new_n668_));
  OAI21_X1  g467(.A(KEYINPUT101), .B1(new_n621_), .B2(new_n622_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n593_), .A2(new_n371_), .A3(new_n619_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n668_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(G29gat), .B1(new_n671_), .B2(new_n524_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n638_), .A2(new_n368_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT105), .Z(new_n674_));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n633_), .A2(KEYINPUT37), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n279_), .A2(new_n202_), .A3(new_n282_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n675_), .B1(new_n593_), .B2(new_n678_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n621_), .A2(KEYINPUT43), .A3(new_n285_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n674_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682_));
  AOI211_X1 g481(.A(new_n213_), .B(new_n525_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n673_), .B(KEYINPUT105), .ZN(new_n684_));
  OAI21_X1  g483(.A(KEYINPUT43), .B1(new_n621_), .B2(new_n285_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n593_), .A2(new_n675_), .A3(new_n678_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n684_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT44), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n672_), .B1(new_n683_), .B2(new_n688_), .ZN(G1328gat));
  INV_X1    g488(.A(KEYINPUT46), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT107), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n690_), .A2(KEYINPUT107), .ZN(new_n692_));
  INV_X1    g491(.A(new_n645_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n693_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n211_), .B1(new_n694_), .B2(new_n688_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n645_), .B(KEYINPUT106), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n696_), .A2(G36gat), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n671_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT45), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n671_), .A2(KEYINPUT45), .A3(new_n697_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n691_), .B(new_n692_), .C1(new_n695_), .C2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n688_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n645_), .B1(new_n687_), .B2(KEYINPUT44), .ZN(new_n705_));
  OAI21_X1  g504(.A(G36gat), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n701_), .ZN(new_n707_));
  AOI21_X1  g506(.A(KEYINPUT45), .B1(new_n671_), .B2(new_n697_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n706_), .A2(new_n709_), .A3(KEYINPUT107), .A4(new_n690_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n703_), .A2(new_n710_), .ZN(G1329gat));
  OAI211_X1 g510(.A(G43gat), .B(new_n574_), .C1(new_n687_), .C2(KEYINPUT44), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n671_), .A2(new_n574_), .ZN(new_n713_));
  OAI22_X1  g512(.A1(new_n704_), .A2(new_n712_), .B1(new_n713_), .B2(G43gat), .ZN(new_n714_));
  XOR2_X1   g513(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n715_));
  XNOR2_X1  g514(.A(new_n714_), .B(new_n715_), .ZN(G1330gat));
  OAI21_X1  g515(.A(new_n552_), .B1(new_n687_), .B2(KEYINPUT44), .ZN(new_n717_));
  OAI21_X1  g516(.A(G50gat), .B1(new_n704_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n671_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n548_), .A2(new_n551_), .A3(G50gat), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT109), .Z(new_n721_));
  OAI21_X1  g520(.A(new_n718_), .B1(new_n719_), .B2(new_n721_), .ZN(G1331gat));
  NOR2_X1   g521(.A1(new_n621_), .A2(new_n619_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n330_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n678_), .A2(new_n367_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n723_), .A2(new_n724_), .A3(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(G57gat), .B1(new_n726_), .B2(new_n524_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n330_), .A2(new_n619_), .A3(new_n367_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n637_), .A2(new_n728_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n525_), .A2(KEYINPUT110), .ZN(new_n730_));
  MUX2_X1   g529(.A(KEYINPUT110), .B(new_n730_), .S(G57gat), .Z(new_n731_));
  AOI21_X1  g530(.A(new_n727_), .B1(new_n729_), .B2(new_n731_), .ZN(G1332gat));
  INV_X1    g531(.A(G64gat), .ZN(new_n733_));
  INV_X1    g532(.A(new_n696_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n726_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n729_), .A2(new_n734_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(G64gat), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n737_), .A2(KEYINPUT48), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n737_), .A2(KEYINPUT48), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n738_), .B2(new_n739_), .ZN(G1333gat));
  NAND3_X1  g539(.A1(new_n726_), .A2(new_n299_), .A3(new_n574_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT112), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n637_), .A2(new_n574_), .A3(new_n728_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n743_), .B2(G71gat), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n743_), .A2(new_n742_), .A3(G71gat), .ZN(new_n746_));
  XOR2_X1   g545(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n747_));
  AND3_X1   g546(.A1(new_n745_), .A2(new_n746_), .A3(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n741_), .B1(new_n748_), .B2(new_n749_), .ZN(G1334gat));
  NAND2_X1  g549(.A1(new_n552_), .A2(new_n297_), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT113), .Z(new_n752_));
  NAND2_X1  g551(.A1(new_n726_), .A2(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT103), .B1(new_n593_), .B2(new_n635_), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n621_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n552_), .B(new_n728_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT50), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n756_), .A2(new_n757_), .A3(G78gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n756_), .B2(G78gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n753_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT114), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n760_), .B(new_n761_), .ZN(G1335gat));
  NOR3_X1   g561(.A1(new_n330_), .A2(new_n368_), .A3(new_n635_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n723_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n765_), .A2(new_n236_), .A3(new_n524_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT115), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n767_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n330_), .A2(new_n368_), .A3(new_n619_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT116), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n685_), .A2(new_n686_), .A3(KEYINPUT115), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n768_), .A2(new_n770_), .A3(new_n771_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n772_), .A2(new_n524_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n766_), .B1(new_n773_), .B2(new_n236_), .ZN(G1336gat));
  AOI21_X1  g573(.A(G92gat), .B1(new_n765_), .B2(new_n645_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n696_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n772_), .B2(new_n776_), .ZN(G1337gat));
  NAND4_X1  g576(.A1(new_n768_), .A2(new_n574_), .A3(new_n770_), .A4(new_n771_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(G99gat), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n765_), .A2(new_n574_), .A3(new_n232_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g581(.A1(new_n765_), .A2(new_n233_), .A3(new_n552_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n552_), .B(new_n770_), .C1(new_n679_), .C2(new_n680_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n784_), .A2(new_n785_), .A3(G106gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n784_), .B2(G106gat), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n783_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g588(.A(KEYINPUT54), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n725_), .A2(new_n790_), .A3(new_n622_), .A4(new_n330_), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT54), .B1(new_n369_), .B2(new_n619_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  OAI22_X1  g593(.A1(new_n314_), .A2(new_n315_), .B1(new_n312_), .B2(new_n260_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n286_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n316_), .A2(new_n797_), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n311_), .B(KEYINPUT55), .C1(new_n314_), .C2(new_n315_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n796_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n326_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT56), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n803_), .B2(KEYINPUT118), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n801_), .A2(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n320_), .A2(new_n326_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n805_), .A2(new_n618_), .A3(new_n615_), .A4(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n800_), .A2(new_n802_), .A3(new_n326_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT118), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT56), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(KEYINPUT119), .B1(new_n808_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n809_), .A2(new_n810_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n803_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n615_), .A2(new_n618_), .A3(new_n807_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT119), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n814_), .A2(new_n815_), .A3(new_n816_), .A4(new_n805_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n612_), .A2(new_n602_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n598_), .A2(new_n601_), .A3(new_n613_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n596_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n607_), .A2(new_n608_), .A3(new_n605_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT78), .B1(new_n601_), .B2(new_n610_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n613_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n597_), .B1(new_n823_), .B2(new_n603_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n820_), .A2(new_n824_), .ZN(new_n825_));
  OR2_X1    g624(.A1(new_n825_), .A2(new_n329_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n812_), .A2(new_n817_), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n635_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT121), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n807_), .B1(new_n820_), .B2(new_n824_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n803_), .B1(new_n800_), .B2(new_n326_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n800_), .A2(new_n803_), .A3(new_n326_), .ZN(new_n835_));
  AOI21_X1  g634(.A(KEYINPUT58), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n831_), .B1(new_n836_), .B2(new_n285_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n801_), .A2(KEYINPUT56), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n613_), .B1(new_n609_), .B2(new_n611_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n819_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n597_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n596_), .B1(new_n617_), .B2(new_n604_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n806_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n838_), .A2(new_n835_), .A3(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n678_), .A2(KEYINPUT121), .A3(new_n846_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n838_), .A2(KEYINPUT58), .A3(new_n843_), .A4(new_n835_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT122), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n848_), .B(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n837_), .A2(new_n847_), .A3(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n829_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n827_), .A2(new_n635_), .A3(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n830_), .A2(new_n851_), .A3(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n794_), .B1(new_n854_), .B2(new_n367_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n645_), .A2(new_n581_), .A3(new_n525_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(G113gat), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n858_), .A2(new_n859_), .A3(new_n619_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n861_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n851_), .A2(new_n853_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n368_), .B1(new_n863_), .B2(new_n830_), .ZN(new_n864_));
  OAI211_X1 g663(.A(KEYINPUT59), .B(new_n856_), .C1(new_n864_), .C2(new_n794_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n622_), .B1(new_n862_), .B2(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n860_), .B1(new_n866_), .B2(new_n859_), .ZN(G1340gat));
  INV_X1    g666(.A(KEYINPUT123), .ZN(new_n868_));
  INV_X1    g667(.A(G120gat), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n862_), .A2(new_n865_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n870_), .B2(new_n724_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n858_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n869_), .B1(new_n330_), .B2(KEYINPUT60), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(KEYINPUT60), .B2(new_n869_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n872_), .A2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n868_), .B1(new_n871_), .B2(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n330_), .B1(new_n862_), .B2(new_n865_), .ZN(new_n877_));
  OAI221_X1 g676(.A(KEYINPUT123), .B1(new_n872_), .B2(new_n874_), .C1(new_n877_), .C2(new_n869_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(G1341gat));
  INV_X1    g678(.A(G127gat), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n880_), .B1(new_n870_), .B2(new_n368_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n368_), .A2(new_n880_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n872_), .A2(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(KEYINPUT124), .B1(new_n881_), .B2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT124), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n367_), .B1(new_n862_), .B2(new_n865_), .ZN(new_n886_));
  OAI221_X1 g685(.A(new_n885_), .B1(new_n872_), .B2(new_n882_), .C1(new_n886_), .C2(new_n880_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n884_), .A2(new_n887_), .ZN(G1342gat));
  AOI21_X1  g687(.A(G134gat), .B1(new_n858_), .B2(new_n633_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT125), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n890_), .ZN(new_n892_));
  AND2_X1   g691(.A1(new_n678_), .A2(G134gat), .ZN(new_n893_));
  AOI22_X1  g692(.A1(new_n891_), .A2(new_n892_), .B1(new_n870_), .B2(new_n893_), .ZN(G1343gat));
  NOR4_X1   g693(.A1(new_n855_), .A2(new_n585_), .A3(new_n525_), .A4(new_n734_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n619_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n724_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g698(.A1(new_n895_), .A2(new_n368_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(KEYINPUT61), .B(G155gat), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(G1346gat));
  INV_X1    g701(.A(G162gat), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n895_), .A2(new_n903_), .A3(new_n633_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n895_), .A2(new_n678_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n905_), .B2(new_n903_), .ZN(G1347gat));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n696_), .A2(new_n581_), .A3(new_n524_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n855_), .A2(new_n622_), .A3(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(KEYINPUT126), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(G169gat), .B1(new_n910_), .B2(KEYINPUT126), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n907_), .B1(new_n912_), .B2(new_n913_), .ZN(new_n914_));
  OR2_X1    g713(.A1(new_n910_), .A2(KEYINPUT126), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n915_), .A2(KEYINPUT62), .A3(new_n911_), .A4(G169gat), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n910_), .A2(new_n475_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n914_), .A2(new_n916_), .A3(new_n917_), .ZN(G1348gat));
  NOR2_X1   g717(.A1(new_n855_), .A2(new_n909_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(new_n724_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n453_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n921_), .B1(new_n464_), .B2(new_n920_), .ZN(G1349gat));
  NAND2_X1  g721(.A1(new_n919_), .A2(new_n368_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n459_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n924_), .B1(new_n442_), .B2(new_n923_), .ZN(G1350gat));
  INV_X1    g724(.A(new_n919_), .ZN(new_n926_));
  OAI21_X1  g725(.A(G190gat), .B1(new_n926_), .B2(new_n285_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n919_), .A2(new_n456_), .A3(new_n633_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(G1351gat));
  NOR4_X1   g728(.A1(new_n855_), .A2(new_n585_), .A3(new_n524_), .A4(new_n696_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(new_n619_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g731(.A1(new_n930_), .A2(new_n424_), .A3(new_n724_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n855_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n585_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n696_), .A2(new_n524_), .ZN(new_n936_));
  NAND4_X1  g735(.A1(new_n934_), .A2(new_n935_), .A3(new_n724_), .A4(new_n936_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(new_n431_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n933_), .A2(new_n938_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(KEYINPUT127), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT127), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n933_), .A2(new_n938_), .A3(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n940_), .A2(new_n942_), .ZN(G1353gat));
  NAND2_X1  g742(.A1(new_n930_), .A2(new_n368_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n944_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n945_));
  XOR2_X1   g744(.A(KEYINPUT63), .B(G211gat), .Z(new_n946_));
  OAI21_X1  g745(.A(new_n945_), .B1(new_n944_), .B2(new_n946_), .ZN(G1354gat));
  INV_X1    g746(.A(G218gat), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n930_), .A2(new_n948_), .A3(new_n633_), .ZN(new_n949_));
  AND2_X1   g748(.A1(new_n930_), .A2(new_n678_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n949_), .B1(new_n950_), .B2(new_n948_), .ZN(G1355gat));
endmodule


