//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 1 1 1 0 1 0 0 1 0 0 0 0 0 1 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_;
  XNOR2_X1  g000(.A(G120gat), .B(G148gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT5), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT73), .ZN(new_n204_));
  XOR2_X1   g003(.A(G176gat), .B(G204gat), .Z(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT74), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT6), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n208_), .B(KEYINPUT6), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT65), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT7), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n212_), .A2(new_n214_), .A3(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(KEYINPUT66), .B(KEYINPUT8), .Z(new_n218_));
  XNOR2_X1  g017(.A(G85gat), .B(G92gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n219_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT7), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n215_), .B(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n221_), .B1(new_n223_), .B2(new_n210_), .ZN(new_n224_));
  AOI22_X1  g023(.A1(new_n217_), .A2(new_n220_), .B1(KEYINPUT8), .B2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n212_), .A2(new_n214_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT9), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(G85gat), .A3(G92gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT10), .B(G99gat), .ZN(new_n229_));
  OAI221_X1 g028(.A(new_n228_), .B1(new_n219_), .B2(new_n227_), .C1(G106gat), .C2(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n226_), .A2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n225_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G57gat), .B(G64gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT11), .ZN(new_n234_));
  XOR2_X1   g033(.A(G71gat), .B(G78gat), .Z(new_n235_));
  OR2_X1    g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n235_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n233_), .A2(KEYINPUT11), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n236_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n232_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT67), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n232_), .A2(new_n242_), .A3(new_n239_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n232_), .A2(new_n239_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT69), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n241_), .A2(KEYINPUT68), .A3(new_n243_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n246_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G230gat), .A2(G233gat), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n251_), .B(KEYINPUT64), .Z(new_n252_));
  NAND3_X1  g051(.A1(new_n250_), .A2(KEYINPUT70), .A3(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n252_), .B1(new_n232_), .B2(new_n239_), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n254_), .A2(KEYINPUT72), .ZN(new_n255_));
  INV_X1    g054(.A(new_n252_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n240_), .A2(KEYINPUT72), .A3(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT12), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n258_), .B1(new_n232_), .B2(new_n239_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT71), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n231_), .A2(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT71), .B1(new_n226_), .B2(new_n230_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n225_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  OR2_X1    g062(.A1(new_n239_), .A2(new_n258_), .ZN(new_n264_));
  OR2_X1    g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n255_), .A2(new_n257_), .A3(new_n259_), .A4(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n253_), .A2(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(KEYINPUT70), .B1(new_n250_), .B2(new_n252_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n207_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n250_), .A2(new_n252_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n272_), .A2(new_n253_), .A3(new_n266_), .A4(new_n206_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n269_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT75), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT13), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(KEYINPUT75), .A2(KEYINPUT13), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n275_), .A2(new_n276_), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n269_), .A2(new_n273_), .A3(new_n278_), .A4(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n277_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G29gat), .B(G36gat), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n282_), .A2(KEYINPUT78), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(KEYINPUT78), .ZN(new_n284_));
  XOR2_X1   g083(.A(G43gat), .B(G50gat), .Z(new_n285_));
  OR3_X1    g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n285_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G15gat), .B(G22gat), .ZN(new_n289_));
  INV_X1    g088(.A(G1gat), .ZN(new_n290_));
  INV_X1    g089(.A(G8gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT14), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G1gat), .B(G8gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n288_), .B(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G229gat), .A2(G233gat), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT83), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n288_), .A2(KEYINPUT15), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT15), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n286_), .A2(new_n287_), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  MUX2_X1   g104(.A(new_n288_), .B(new_n305_), .S(new_n295_), .Z(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(new_n297_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n301_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G113gat), .B(G141gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G169gat), .B(G197gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n311_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n301_), .A2(new_n307_), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n281_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT27), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT98), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT21), .ZN(new_n320_));
  INV_X1    g119(.A(G211gat), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n321_), .A2(G218gat), .ZN(new_n322_));
  INV_X1    g121(.A(G218gat), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n323_), .A2(G211gat), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n320_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G197gat), .B(G204gat), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n323_), .A2(G211gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n321_), .A2(G218gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n328_), .A2(new_n329_), .A3(KEYINPUT21), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n325_), .A2(new_n327_), .A3(new_n330_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n326_), .A2(KEYINPUT21), .A3(new_n328_), .A4(new_n329_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G183gat), .A2(G190gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT23), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT23), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n336_), .A2(G183gat), .A3(G190gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(G183gat), .ZN(new_n339_));
  INV_X1    g138(.A(G190gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT22), .ZN(new_n343_));
  OAI211_X1 g142(.A(KEYINPUT85), .B(G169gat), .C1(new_n343_), .C2(KEYINPUT84), .ZN(new_n344_));
  NAND2_X1  g143(.A1(KEYINPUT85), .A2(G169gat), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT84), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(new_n346_), .A3(KEYINPUT22), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT85), .ZN(new_n348_));
  INV_X1    g147(.A(G169gat), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n348_), .B1(new_n349_), .B2(KEYINPUT22), .ZN(new_n350_));
  INV_X1    g149(.A(G176gat), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n344_), .A2(new_n347_), .A3(new_n350_), .A4(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G169gat), .A2(G176gat), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n342_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n339_), .A2(KEYINPUT25), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT25), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(G183gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n340_), .A2(KEYINPUT26), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT26), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(G190gat), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n355_), .A2(new_n357_), .A3(new_n358_), .A4(new_n360_), .ZN(new_n361_));
  OR3_X1    g160(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n349_), .A2(new_n351_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(KEYINPUT24), .A3(new_n353_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n361_), .A2(new_n338_), .A3(new_n362_), .A4(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n354_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT86), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT86), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n354_), .A2(new_n368_), .A3(new_n365_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n333_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n343_), .A2(G169gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n349_), .A2(KEYINPUT22), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(new_n372_), .A3(new_n351_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n353_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT97), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT97), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n373_), .A2(new_n376_), .A3(new_n353_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(new_n342_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n358_), .A2(new_n360_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT96), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n355_), .A2(new_n357_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n358_), .A2(new_n360_), .A3(KEYINPUT96), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n338_), .A2(new_n364_), .A3(new_n362_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n333_), .A2(new_n378_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388_));
  XOR2_X1   g187(.A(new_n388_), .B(KEYINPUT19), .Z(new_n389_));
  AND2_X1   g188(.A1(new_n389_), .A2(KEYINPUT20), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n387_), .A2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n319_), .B1(new_n370_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n331_), .A2(new_n332_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n354_), .A2(new_n368_), .A3(new_n365_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n368_), .B1(new_n354_), .B2(new_n365_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n393_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n396_), .A2(KEYINPUT98), .A3(new_n387_), .A4(new_n390_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n392_), .A2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n393_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n378_), .A2(new_n393_), .A3(new_n386_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT20), .B1(new_n399_), .B2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n389_), .B(KEYINPUT95), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G64gat), .B(G92gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT100), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G8gat), .B(G36gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n398_), .A2(new_n404_), .A3(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n411_), .B1(new_n398_), .B2(new_n404_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n318_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT104), .B(KEYINPUT20), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n367_), .A2(new_n369_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n415_), .B1(new_n416_), .B2(new_n393_), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n378_), .A2(KEYINPUT105), .A3(new_n386_), .ZN(new_n418_));
  AOI21_X1  g217(.A(KEYINPUT105), .B1(new_n378_), .B2(new_n386_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n333_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n389_), .B1(new_n417_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT20), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n333_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n423_));
  AOI211_X1 g222(.A(new_n422_), .B(new_n403_), .C1(new_n423_), .C2(new_n400_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n410_), .B1(new_n421_), .B2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n398_), .A2(new_n404_), .A3(new_n411_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n426_), .A3(KEYINPUT27), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n414_), .A2(KEYINPUT107), .A3(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(KEYINPUT107), .B1(new_n414_), .B2(new_n427_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT106), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT94), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT93), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n432_), .B1(new_n433_), .B2(KEYINPUT3), .ZN(new_n434_));
  NOR2_X1   g233(.A1(G141gat), .A2(G148gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  OAI221_X1 g235(.A(new_n432_), .B1(G141gat), .B2(G148gat), .C1(new_n433_), .C2(KEYINPUT3), .ZN(new_n437_));
  NAND3_X1  g236(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G141gat), .A2(G148gat), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT2), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT3), .ZN(new_n441_));
  AOI22_X1  g240(.A1(new_n439_), .A2(new_n440_), .B1(new_n441_), .B2(KEYINPUT94), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .A4(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(G155gat), .A2(G162gat), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G155gat), .A2(G162gat), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n443_), .A2(new_n447_), .ZN(new_n448_));
  XOR2_X1   g247(.A(G141gat), .B(G148gat), .Z(new_n449_));
  INV_X1    g248(.A(KEYINPUT92), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n446_), .A2(new_n450_), .A3(KEYINPUT1), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n451_), .B(new_n445_), .C1(KEYINPUT1), .C2(new_n446_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n450_), .B1(new_n446_), .B2(KEYINPUT1), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n449_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n448_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(G134gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(G127gat), .ZN(new_n457_));
  INV_X1    g256(.A(G127gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(G134gat), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT90), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n457_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n460_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT91), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n458_), .A2(G134gat), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n456_), .A2(G127gat), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT90), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT91), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n457_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G113gat), .B(G120gat), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n463_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n471_), .B1(new_n463_), .B2(new_n469_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n455_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G225gat), .A2(G233gat), .ZN(new_n475_));
  NOR3_X1   g274(.A1(new_n461_), .A2(new_n462_), .A3(KEYINPUT91), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n467_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n470_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n448_), .A2(new_n454_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n463_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n474_), .A2(new_n475_), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT4), .B1(new_n448_), .B2(new_n454_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n484_), .A2(new_n480_), .A3(new_n478_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT101), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT101), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n484_), .A2(new_n478_), .A3(new_n487_), .A4(new_n480_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n475_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n474_), .A2(KEYINPUT4), .A3(new_n481_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n483_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G1gat), .B(G29gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT0), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(G57gat), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n492_), .A2(KEYINPUT0), .ZN(new_n495_));
  INV_X1    g294(.A(G57gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n492_), .A2(KEYINPUT0), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n494_), .A2(new_n498_), .A3(G85gat), .ZN(new_n499_));
  AOI21_X1  g298(.A(G85gat), .B1(new_n494_), .B2(new_n498_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n431_), .B1(new_n491_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n475_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n472_), .A2(new_n473_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n487_), .B1(new_n505_), .B2(new_n484_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n488_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n490_), .B(new_n504_), .C1(new_n506_), .C2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(new_n482_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n509_), .A2(KEYINPUT106), .A3(new_n501_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n508_), .A2(new_n482_), .A3(new_n502_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n503_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT29), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n455_), .A2(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n515_), .B(KEYINPUT28), .Z(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G228gat), .A2(G233gat), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n393_), .B(new_n518_), .C1(new_n455_), .C2(new_n514_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n514_), .B1(new_n448_), .B2(new_n454_), .ZN(new_n520_));
  OAI211_X1 g319(.A(G228gat), .B(G233gat), .C1(new_n520_), .C2(new_n333_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G78gat), .B(G106gat), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n519_), .A2(new_n521_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n523_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n526_));
  XOR2_X1   g325(.A(G22gat), .B(G50gat), .Z(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NOR3_X1   g327(.A1(new_n525_), .A2(new_n526_), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n519_), .A2(new_n521_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(new_n522_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n527_), .B1(new_n531_), .B2(new_n524_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n517_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n528_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n531_), .A2(new_n524_), .A3(new_n527_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(new_n516_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n533_), .A2(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(KEYINPUT87), .B(KEYINPUT30), .Z(new_n538_));
  OAI21_X1  g337(.A(new_n538_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n538_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n367_), .A2(new_n369_), .A3(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G15gat), .B(G43gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT88), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G71gat), .B(G99gat), .ZN(new_n544_));
  AND2_X1   g343(.A1(G227gat), .A2(G233gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n543_), .B(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n539_), .A2(new_n541_), .A3(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n539_), .A2(new_n541_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n547_), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT89), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT89), .ZN(new_n552_));
  AOI211_X1 g351(.A(new_n552_), .B(new_n547_), .C1(new_n539_), .C2(new_n541_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n548_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT31), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT31), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n556_), .B(new_n548_), .C1(new_n551_), .C2(new_n553_), .ZN(new_n557_));
  AND3_X1   g356(.A1(new_n555_), .A2(new_n505_), .A3(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n505_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n513_), .B(new_n537_), .C1(new_n558_), .C2(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(KEYINPUT108), .B1(new_n430_), .B2(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n558_), .A2(new_n559_), .ZN(new_n562_));
  AND3_X1   g361(.A1(new_n534_), .A2(new_n535_), .A3(new_n516_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n516_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n398_), .A2(new_n404_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n421_), .A2(new_n424_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT32), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n410_), .A2(new_n568_), .ZN(new_n569_));
  MUX2_X1   g368(.A(new_n566_), .B(new_n567_), .S(new_n569_), .Z(new_n570_));
  NAND2_X1  g369(.A1(new_n512_), .A2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n412_), .A2(new_n413_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n474_), .A2(new_n504_), .A3(new_n481_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(new_n501_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n504_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n574_), .B1(new_n575_), .B2(new_n490_), .ZN(new_n576_));
  XOR2_X1   g375(.A(KEYINPUT103), .B(KEYINPUT33), .Z(new_n577_));
  AOI21_X1  g376(.A(new_n576_), .B1(new_n511_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT33), .ZN(new_n579_));
  OAI21_X1  g378(.A(KEYINPUT102), .B1(new_n511_), .B2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT102), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n491_), .A2(new_n581_), .A3(KEYINPUT33), .A4(new_n502_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n572_), .A2(new_n578_), .A3(new_n580_), .A4(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n565_), .B1(new_n571_), .B2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n414_), .A2(new_n427_), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n585_), .A2(new_n512_), .A3(new_n537_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n562_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT107), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n566_), .A2(new_n410_), .ZN(new_n589_));
  AOI21_X1  g388(.A(KEYINPUT27), .B1(new_n589_), .B2(new_n426_), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n425_), .A2(new_n426_), .A3(KEYINPUT27), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n588_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n414_), .A2(KEYINPUT107), .A3(new_n427_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n555_), .A2(new_n557_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n505_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n555_), .A2(new_n505_), .A3(new_n557_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n565_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT108), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n594_), .A2(new_n599_), .A3(new_n600_), .A4(new_n513_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n561_), .A2(new_n587_), .A3(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n317_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT81), .ZN(new_n604_));
  XOR2_X1   g403(.A(G190gat), .B(G218gat), .Z(new_n605_));
  XNOR2_X1  g404(.A(G134gat), .B(G162gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT36), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n232_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n609_));
  XOR2_X1   g408(.A(KEYINPUT76), .B(KEYINPUT34), .Z(new_n610_));
  NAND2_X1  g409(.A1(G232gat), .A2(G233gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n612_), .A2(KEYINPUT35), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n609_), .B(new_n613_), .C1(new_n263_), .C2(new_n305_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(KEYINPUT35), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT77), .ZN(new_n616_));
  OAI21_X1  g415(.A(KEYINPUT79), .B1(new_n263_), .B2(new_n305_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n614_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n614_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n608_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n614_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n617_), .A2(new_n616_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT36), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n624_), .A2(new_n625_), .A3(new_n607_), .A4(new_n618_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n621_), .A2(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n604_), .B1(new_n627_), .B2(KEYINPUT37), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT37), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n621_), .A2(new_n626_), .A3(KEYINPUT81), .A4(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(KEYINPUT80), .B1(new_n627_), .B2(KEYINPUT37), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT80), .ZN(new_n632_));
  AOI211_X1 g431(.A(new_n632_), .B(new_n629_), .C1(new_n621_), .C2(new_n626_), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n628_), .B(new_n630_), .C1(new_n631_), .C2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(G231gat), .A2(G233gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n295_), .B(new_n636_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n637_), .B(new_n239_), .Z(new_n638_));
  XOR2_X1   g437(.A(G127gat), .B(G155gat), .Z(new_n639_));
  XNOR2_X1  g438(.A(G183gat), .B(G211gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  XOR2_X1   g440(.A(KEYINPUT82), .B(KEYINPUT16), .Z(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT17), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n638_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(KEYINPUT17), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n645_), .B1(new_n647_), .B2(new_n638_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n635_), .A2(new_n649_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n603_), .A2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n651_), .A2(new_n290_), .A3(new_n512_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT38), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n602_), .A2(new_n627_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n317_), .A2(new_n654_), .A3(new_n648_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G1gat), .B1(new_n655_), .B2(new_n513_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n653_), .A2(new_n656_), .ZN(G1324gat));
  INV_X1    g456(.A(KEYINPUT39), .ZN(new_n658_));
  OAI21_X1  g457(.A(G8gat), .B1(new_n655_), .B2(new_n594_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(KEYINPUT109), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n659_), .A2(KEYINPUT109), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n658_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n662_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n664_), .A2(KEYINPUT39), .A3(new_n660_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n651_), .A2(new_n291_), .A3(new_n430_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n663_), .A2(new_n665_), .A3(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT40), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n663_), .A2(new_n665_), .A3(KEYINPUT40), .A4(new_n666_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1325gat));
  INV_X1    g470(.A(G15gat), .ZN(new_n672_));
  INV_X1    g471(.A(new_n562_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n651_), .A2(new_n672_), .A3(new_n673_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT110), .Z(new_n675_));
  OAI21_X1  g474(.A(G15gat), .B1(new_n655_), .B2(new_n562_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT41), .Z(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(G1326gat));
  OAI21_X1  g477(.A(G22gat), .B1(new_n655_), .B2(new_n537_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT42), .ZN(new_n680_));
  INV_X1    g479(.A(G22gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n651_), .A2(new_n681_), .A3(new_n565_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(G1327gat));
  NOR2_X1   g482(.A1(new_n627_), .A2(new_n648_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n603_), .A2(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(G29gat), .B1(new_n685_), .B2(new_n512_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n602_), .A2(new_n635_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT112), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT111), .B1(new_n602_), .B2(new_n635_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n689_), .B(new_n690_), .C1(new_n688_), .C2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT111), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n687_), .A2(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n694_), .A2(KEYINPUT112), .A3(KEYINPUT43), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n281_), .A2(new_n316_), .A3(new_n648_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n692_), .A2(new_n695_), .A3(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n699_), .A2(G29gat), .A3(new_n512_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n692_), .A2(KEYINPUT44), .A3(new_n695_), .A4(new_n696_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n686_), .B1(new_n700_), .B2(new_n701_), .ZN(G1328gat));
  NAND3_X1  g501(.A1(new_n699_), .A2(new_n430_), .A3(new_n701_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(G36gat), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n594_), .A2(G36gat), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n603_), .A2(new_n684_), .A3(new_n705_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT45), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n704_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT46), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n704_), .A2(KEYINPUT46), .A3(new_n707_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1329gat));
  NAND2_X1  g511(.A1(new_n699_), .A2(new_n701_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n673_), .A2(G43gat), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n685_), .A2(new_n673_), .ZN(new_n715_));
  OAI22_X1  g514(.A1(new_n713_), .A2(new_n714_), .B1(new_n715_), .B2(G43gat), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g516(.A(G50gat), .B1(new_n685_), .B2(new_n565_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n699_), .A2(G50gat), .A3(new_n565_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n719_), .B2(new_n701_), .ZN(G1331gat));
  NAND4_X1  g519(.A1(new_n654_), .A2(new_n316_), .A3(new_n281_), .A4(new_n648_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT113), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n722_), .A2(G57gat), .A3(new_n512_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT114), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n281_), .A2(new_n602_), .A3(new_n316_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n650_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(G57gat), .B1(new_n727_), .B2(new_n512_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n724_), .A2(new_n728_), .ZN(G1332gat));
  OR3_X1    g528(.A1(new_n726_), .A2(G64gat), .A3(new_n594_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n722_), .A2(new_n430_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(KEYINPUT115), .B(KEYINPUT48), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n731_), .A2(G64gat), .A3(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n731_), .B2(G64gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n730_), .B1(new_n733_), .B2(new_n734_), .ZN(G1333gat));
  OR3_X1    g534(.A1(new_n726_), .A2(G71gat), .A3(new_n562_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n722_), .A2(new_n673_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(G71gat), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(KEYINPUT49), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(KEYINPUT49), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n736_), .B1(new_n739_), .B2(new_n740_), .ZN(G1334gat));
  NAND2_X1  g540(.A1(new_n722_), .A2(new_n565_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(G78gat), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n743_), .A2(KEYINPUT50), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(KEYINPUT50), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n537_), .A2(G78gat), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT116), .ZN(new_n747_));
  OAI22_X1  g546(.A1(new_n744_), .A2(new_n745_), .B1(new_n726_), .B2(new_n747_), .ZN(G1335gat));
  INV_X1    g547(.A(new_n281_), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n749_), .A2(new_n315_), .A3(new_n648_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n692_), .A2(new_n695_), .A3(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT117), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT117), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n692_), .A2(new_n753_), .A3(new_n695_), .A4(new_n750_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n513_), .B1(new_n752_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(G85gat), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n725_), .A2(new_n684_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n512_), .A2(new_n756_), .ZN(new_n758_));
  OAI22_X1  g557(.A1(new_n755_), .A2(new_n756_), .B1(new_n757_), .B2(new_n758_), .ZN(G1336gat));
  AOI21_X1  g558(.A(new_n594_), .B1(new_n752_), .B2(new_n754_), .ZN(new_n760_));
  INV_X1    g559(.A(G92gat), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n430_), .A2(new_n761_), .ZN(new_n762_));
  OAI22_X1  g561(.A1(new_n760_), .A2(new_n761_), .B1(new_n757_), .B2(new_n762_), .ZN(G1337gat));
  AOI21_X1  g562(.A(new_n562_), .B1(new_n752_), .B2(new_n754_), .ZN(new_n764_));
  INV_X1    g563(.A(G99gat), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n562_), .A2(new_n229_), .ZN(new_n766_));
  OAI22_X1  g565(.A1(new_n764_), .A2(new_n765_), .B1(new_n757_), .B2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT51), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n769_));
  OAI221_X1 g568(.A(new_n769_), .B1(new_n757_), .B2(new_n766_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(G1338gat));
  NAND4_X1  g570(.A1(new_n692_), .A2(new_n565_), .A3(new_n695_), .A4(new_n750_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n772_), .A2(new_n773_), .A3(G106gat), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n773_), .B1(new_n772_), .B2(G106gat), .ZN(new_n775_));
  OR2_X1    g574(.A1(new_n537_), .A2(G106gat), .ZN(new_n776_));
  OAI22_X1  g575(.A1(new_n774_), .A2(new_n775_), .B1(new_n757_), .B2(new_n776_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n266_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n265_), .A2(new_n259_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n782_), .A2(KEYINPUT55), .A3(new_n257_), .A4(new_n255_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n252_), .B1(new_n781_), .B2(new_n244_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n780_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n785_), .A2(KEYINPUT56), .A3(new_n207_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT56), .B1(new_n785_), .B2(new_n207_), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n273_), .A2(new_n315_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n306_), .A2(new_n298_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n313_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n793_), .A2(KEYINPUT120), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(KEYINPUT120), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n794_), .A2(new_n314_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n274_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n790_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(KEYINPUT57), .A3(new_n627_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT121), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n786_), .A2(new_n787_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n273_), .A2(new_n796_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n800_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT58), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT58), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n800_), .B(new_n805_), .C1(new_n801_), .C2(new_n802_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n804_), .A2(new_n635_), .A3(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n788_), .A2(new_n789_), .B1(new_n274_), .B2(new_n796_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n627_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n808_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n799_), .A2(new_n807_), .A3(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n649_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n316_), .A2(KEYINPUT118), .A3(new_n648_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT118), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n315_), .B2(new_n649_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n816_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n277_), .A2(new_n280_), .A3(new_n634_), .A4(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT54), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT119), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n818_), .A2(new_n821_), .A3(KEYINPUT54), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n818_), .A2(KEYINPUT54), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n820_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n813_), .A2(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n430_), .A2(new_n513_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n599_), .A3(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(G113gat), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n829_), .A3(new_n315_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT122), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT59), .B1(new_n825_), .B2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n827_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n599_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n834_), .B1(new_n813_), .B2(new_n824_), .ZN(new_n835_));
  AOI21_X1  g634(.A(KEYINPUT122), .B1(new_n813_), .B2(new_n824_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n826_), .B(new_n835_), .C1(new_n836_), .C2(KEYINPUT59), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n316_), .B1(new_n833_), .B2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n830_), .B1(new_n838_), .B2(new_n829_), .ZN(G1340gat));
  INV_X1    g638(.A(KEYINPUT60), .ZN(new_n840_));
  INV_X1    g639(.A(G120gat), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n281_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n828_), .A2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n749_), .B1(new_n833_), .B2(new_n837_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n845_), .B2(new_n841_), .ZN(G1341gat));
  AOI21_X1  g645(.A(G127gat), .B1(new_n828_), .B2(new_n648_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n833_), .A2(new_n837_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n648_), .A2(KEYINPUT123), .A3(G127gat), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(KEYINPUT123), .B2(G127gat), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n847_), .B1(new_n848_), .B2(new_n850_), .ZN(G1342gat));
  NAND2_X1  g650(.A1(new_n635_), .A2(G134gat), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n833_), .B2(new_n837_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n835_), .A2(new_n810_), .A3(new_n826_), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n854_), .A2(KEYINPUT124), .A3(new_n456_), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT124), .B1(new_n854_), .B2(new_n456_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n853_), .A2(new_n855_), .A3(new_n856_), .ZN(G1343gat));
  NOR2_X1   g656(.A1(new_n673_), .A2(new_n537_), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n825_), .A2(new_n826_), .A3(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n315_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n281_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g662(.A1(new_n859_), .A2(new_n648_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT61), .B(G155gat), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1346gat));
  INV_X1    g665(.A(G162gat), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n859_), .A2(new_n867_), .A3(new_n810_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n859_), .A2(new_n635_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(new_n867_), .ZN(G1347gat));
  NOR2_X1   g669(.A1(new_n594_), .A2(new_n512_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n835_), .A2(new_n315_), .A3(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(G169gat), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT62), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n872_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n371_), .A2(new_n372_), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n875_), .B(new_n876_), .C1(new_n877_), .C2(new_n872_), .ZN(G1348gat));
  AND2_X1   g677(.A1(new_n835_), .A2(new_n871_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n281_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g680(.A1(new_n835_), .A2(new_n648_), .A3(new_n871_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT126), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n835_), .A2(KEYINPUT126), .A3(new_n648_), .A4(new_n871_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n382_), .ZN(new_n887_));
  NAND4_X1  g686(.A1(new_n879_), .A2(KEYINPUT125), .A3(new_n887_), .A4(new_n648_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT125), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n889_), .B1(new_n882_), .B2(new_n382_), .ZN(new_n890_));
  AOI22_X1  g689(.A1(new_n886_), .A2(new_n339_), .B1(new_n888_), .B2(new_n890_), .ZN(G1350gat));
  NAND4_X1  g690(.A1(new_n879_), .A2(new_n810_), .A3(new_n381_), .A4(new_n383_), .ZN(new_n892_));
  AND2_X1   g691(.A1(new_n879_), .A2(new_n635_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n340_), .ZN(G1351gat));
  AND2_X1   g693(.A1(new_n858_), .A2(new_n871_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n825_), .A2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n315_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g698(.A1(new_n896_), .A2(new_n749_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(G1353gat));
  NOR2_X1   g701(.A1(new_n896_), .A2(new_n649_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n904_));
  AND2_X1   g703(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n903_), .B1(new_n904_), .B2(new_n905_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n906_), .B1(new_n903_), .B2(new_n904_), .ZN(G1354gat));
  OAI21_X1  g706(.A(G218gat), .B1(new_n896_), .B2(new_n634_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n810_), .A2(new_n323_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n896_), .B2(new_n909_), .ZN(G1355gat));
endmodule


