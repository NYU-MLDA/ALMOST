//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 0 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 0 0 1 0 1 1 0 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n869_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_;
  INV_X1    g000(.A(KEYINPUT20), .ZN(new_n202_));
  OR2_X1    g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n203_), .A2(KEYINPUT24), .A3(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT76), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(G183gat), .A3(G190gat), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n208_), .A2(KEYINPUT77), .ZN(new_n209_));
  INV_X1    g008(.A(G183gat), .ZN(new_n210_));
  INV_X1    g009(.A(G190gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT23), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n208_), .A2(KEYINPUT77), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n209_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n203_), .A2(KEYINPUT24), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT75), .ZN(new_n216_));
  OR3_X1    g015(.A1(new_n216_), .A2(new_n211_), .A3(KEYINPUT26), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT26), .B1(new_n216_), .B2(new_n211_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT25), .B(G183gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n206_), .A2(new_n214_), .A3(new_n215_), .A4(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n212_), .A2(new_n208_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n222_), .B1(G183gat), .B2(G190gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n204_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT22), .B(G169gat), .ZN(new_n225_));
  INV_X1    g024(.A(G176gat), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n224_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n223_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n221_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT78), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G211gat), .B(G218gat), .ZN(new_n231_));
  INV_X1    g030(.A(G204gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(G197gat), .ZN(new_n233_));
  INV_X1    g032(.A(G197gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(G204gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT21), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n233_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT88), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n238_), .B1(new_n234_), .B2(G204gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n232_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(new_n235_), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n241_), .A2(KEYINPUT89), .A3(KEYINPUT21), .ZN(new_n242_));
  AOI21_X1  g041(.A(KEYINPUT89), .B1(new_n241_), .B2(KEYINPUT21), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n231_), .B(new_n237_), .C1(new_n242_), .C2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT90), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n245_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n231_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n236_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n248_), .A2(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n202_), .B1(new_n230_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G226gat), .A2(G233gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT19), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n251_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n214_), .B1(G183gat), .B2(G190gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(new_n227_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT96), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT26), .B(G190gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n219_), .A2(new_n262_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n263_), .A2(new_n215_), .A3(new_n222_), .A4(new_n205_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT96), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n259_), .A2(new_n265_), .A3(new_n227_), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n261_), .A2(new_n264_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n258_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n254_), .A2(new_n257_), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT97), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n258_), .A2(new_n267_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT78), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n229_), .B(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n258_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n271_), .A2(KEYINPUT20), .A3(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n256_), .B(KEYINPUT95), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT97), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n254_), .A2(new_n279_), .A3(new_n257_), .A4(new_n268_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n270_), .A2(new_n278_), .A3(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G8gat), .B(G36gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(G92gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT18), .B(G64gat), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n283_), .B(new_n284_), .Z(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n281_), .A2(new_n286_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n270_), .A2(new_n278_), .A3(new_n285_), .A4(new_n280_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT98), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT98), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n287_), .A2(new_n291_), .A3(new_n288_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G113gat), .B(G120gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT80), .B(KEYINPUT81), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G127gat), .B(G134gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298_));
  NOR2_X1   g097(.A1(G141gat), .A2(G148gat), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT84), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n303_), .B1(KEYINPUT1), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(KEYINPUT1), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT85), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n298_), .B(new_n300_), .C1(new_n305_), .C2(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n299_), .B(KEYINPUT3), .Z(new_n309_));
  NOR2_X1   g108(.A1(KEYINPUT86), .A2(KEYINPUT2), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(new_n298_), .ZN(new_n311_));
  AOI22_X1  g110(.A1(KEYINPUT86), .A2(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n311_), .B1(new_n312_), .B2(new_n310_), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n303_), .B(new_n304_), .C1(new_n309_), .C2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n308_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n297_), .B(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT4), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G225gat), .A2(G233gat), .ZN(new_n318_));
  INV_X1    g117(.A(new_n297_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT4), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(new_n320_), .A3(new_n315_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n317_), .A2(new_n318_), .A3(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G1gat), .B(G29gat), .ZN(new_n323_));
  INV_X1    g122(.A(G85gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT0), .B(G57gat), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n325_), .B(new_n326_), .Z(new_n327_));
  INV_X1    g126(.A(new_n318_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n316_), .A2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n322_), .A2(new_n327_), .A3(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n317_), .A2(new_n328_), .A3(new_n321_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n316_), .A2(new_n318_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n327_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n331_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT33), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n290_), .A2(new_n292_), .A3(new_n330_), .A4(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n331_), .A2(new_n332_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n327_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(new_n334_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT20), .B1(new_n273_), .B2(new_n258_), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n258_), .A2(new_n264_), .A3(new_n260_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n256_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n271_), .A2(new_n274_), .A3(KEYINPUT20), .A4(new_n276_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n285_), .A2(KEYINPUT32), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n339_), .B(new_n346_), .C1(new_n281_), .C2(new_n345_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT99), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n336_), .A2(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G15gat), .B(G43gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G71gat), .B(G99gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G227gat), .A2(G233gat), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n353_), .B(new_n354_), .Z(new_n355_));
  INV_X1    g154(.A(KEYINPUT79), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n230_), .A2(KEYINPUT30), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT30), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n273_), .A2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n357_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n355_), .B(new_n356_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n358_), .A2(new_n360_), .A3(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n362_), .A2(KEYINPUT83), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT83), .ZN(new_n366_));
  INV_X1    g165(.A(new_n364_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n366_), .B1(new_n367_), .B2(new_n361_), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n297_), .B(KEYINPUT82), .Z(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT31), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n365_), .A2(new_n368_), .A3(new_n371_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n362_), .A2(KEYINPUT83), .A3(new_n370_), .A4(new_n364_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n315_), .A2(KEYINPUT29), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G228gat), .A2(G233gat), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n377_), .B(KEYINPUT87), .Z(new_n378_));
  NAND3_X1  g177(.A1(new_n253_), .A2(new_n376_), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n378_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n376_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n380_), .B1(new_n258_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G78gat), .B(G106gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT91), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  OR2_X1    g185(.A1(new_n315_), .A2(KEYINPUT29), .ZN(new_n387_));
  INV_X1    g186(.A(G50gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT28), .B(G22gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n387_), .B(G50gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n390_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n391_), .A2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n386_), .B1(new_n395_), .B2(KEYINPUT92), .ZN(new_n396_));
  AOI21_X1  g195(.A(KEYINPUT92), .B1(new_n391_), .B2(new_n394_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n386_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n383_), .A2(new_n385_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n383_), .A2(KEYINPUT93), .A3(new_n385_), .ZN(new_n401_));
  AOI21_X1  g200(.A(KEYINPUT93), .B1(new_n383_), .B2(new_n385_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n395_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n396_), .A2(new_n400_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT94), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n396_), .A2(new_n400_), .A3(new_n403_), .A4(KEYINPUT94), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n350_), .A2(new_n375_), .A3(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n339_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT27), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n289_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n344_), .A2(new_n286_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n288_), .A2(new_n413_), .A3(KEYINPUT27), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n406_), .A2(new_n374_), .A3(new_n407_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n374_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n417_));
  OAI211_X1 g216(.A(new_n410_), .B(new_n415_), .C1(new_n416_), .C2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n409_), .A2(new_n418_), .ZN(new_n419_));
  AND2_X1   g218(.A1(G230gat), .A2(G233gat), .ZN(new_n420_));
  XOR2_X1   g219(.A(G85gat), .B(G92gat), .Z(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT9), .ZN(new_n422_));
  AND3_X1   g221(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(G106gat), .ZN(new_n426_));
  INV_X1    g225(.A(G99gat), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n427_), .A2(KEYINPUT10), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(KEYINPUT10), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n426_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(G92gat), .ZN(new_n431_));
  OR3_X1    g230(.A1(new_n324_), .A2(new_n431_), .A3(KEYINPUT9), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n422_), .A2(new_n425_), .A3(new_n430_), .A4(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(G57gat), .ZN(new_n434_));
  INV_X1    g233(.A(G64gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G57gat), .A2(G64gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT11), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G71gat), .B(G78gat), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT11), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n436_), .A2(new_n442_), .A3(new_n437_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n439_), .A2(new_n441_), .A3(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n438_), .A2(new_n440_), .A3(KEYINPUT11), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT8), .ZN(new_n447_));
  NAND2_X1  g246(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n448_));
  OAI22_X1  g247(.A1(KEYINPUT64), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT64), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT7), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n450_), .A2(new_n451_), .A3(new_n427_), .A4(new_n426_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n425_), .A2(new_n448_), .A3(new_n449_), .A4(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n447_), .B1(new_n453_), .B2(new_n421_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n449_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G99gat), .A2(G106gat), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(new_n459_), .A3(new_n448_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n447_), .B(new_n421_), .C1(new_n455_), .C2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n433_), .B(new_n446_), .C1(new_n454_), .C2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n421_), .B1(new_n455_), .B2(new_n460_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT8), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n461_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n446_), .B1(new_n467_), .B2(new_n433_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n420_), .B1(new_n464_), .B2(new_n468_), .ZN(new_n469_));
  AOI211_X1 g268(.A(KEYINPUT12), .B(new_n446_), .C1(new_n467_), .C2(new_n433_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n464_), .A2(new_n468_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n470_), .B1(new_n471_), .B2(KEYINPUT12), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n469_), .B1(new_n472_), .B2(new_n420_), .ZN(new_n473_));
  XOR2_X1   g272(.A(KEYINPUT65), .B(G204gat), .Z(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT5), .B(G176gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G120gat), .B(G148gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n473_), .B(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT13), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G29gat), .B(G36gat), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G43gat), .B(G50gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(G43gat), .B(G50gat), .Z(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n482_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G1gat), .B(G8gat), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT68), .ZN(new_n491_));
  AND2_X1   g290(.A1(KEYINPUT67), .A2(G1gat), .ZN(new_n492_));
  NOR2_X1   g291(.A1(KEYINPUT67), .A2(G1gat), .ZN(new_n493_));
  INV_X1    g292(.A(G8gat), .ZN(new_n494_));
  NOR3_X1   g293(.A1(new_n492_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT14), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n491_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  OR2_X1    g296(.A1(KEYINPUT67), .A2(G1gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(KEYINPUT67), .A2(G1gat), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n498_), .A2(G8gat), .A3(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(KEYINPUT68), .A3(KEYINPUT14), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n497_), .A2(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(G15gat), .B(G22gat), .Z(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n490_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n490_), .ZN(new_n506_));
  AOI211_X1 g305(.A(new_n503_), .B(new_n506_), .C1(new_n497_), .C2(new_n501_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n489_), .B1(new_n505_), .B2(new_n507_), .ZN(new_n508_));
  NOR3_X1   g307(.A1(new_n495_), .A2(new_n491_), .A3(new_n496_), .ZN(new_n509_));
  AOI21_X1  g308(.A(KEYINPUT68), .B1(new_n500_), .B2(KEYINPUT14), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n504_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n506_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT15), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n488_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n485_), .A2(new_n487_), .A3(KEYINPUT15), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n502_), .A2(new_n504_), .A3(new_n490_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n512_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G229gat), .A2(G233gat), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n508_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n512_), .A2(new_n488_), .A3(new_n517_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n519_), .B1(new_n508_), .B2(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G113gat), .B(G141gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G169gat), .B(G197gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n523_), .A2(KEYINPUT73), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT73), .ZN(new_n529_));
  INV_X1    g328(.A(new_n519_), .ZN(new_n530_));
  NOR3_X1   g329(.A1(new_n505_), .A2(new_n507_), .A3(new_n489_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n488_), .B1(new_n512_), .B2(new_n517_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n530_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n508_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n529_), .B1(new_n535_), .B2(new_n526_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n528_), .A2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n526_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT72), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT72), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n535_), .A2(new_n540_), .A3(new_n526_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT74), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n537_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n543_), .B1(new_n537_), .B2(new_n542_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n481_), .A2(new_n546_), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n419_), .A2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n433_), .B1(new_n454_), .B2(new_n462_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n549_), .A2(new_n516_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n488_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G232gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT34), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT35), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n555_), .A2(new_n556_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n552_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT36), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G190gat), .B(G218gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G134gat), .B(G162gat), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n562_), .B(new_n563_), .Z(new_n564_));
  OAI211_X1 g363(.A(KEYINPUT35), .B(new_n554_), .C1(new_n550_), .C2(new_n551_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n560_), .A2(new_n561_), .A3(new_n564_), .A4(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT66), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n560_), .A2(new_n565_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n564_), .B(KEYINPUT36), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n567_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT37), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n567_), .A2(new_n570_), .A3(KEYINPUT37), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G127gat), .B(G155gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(G211gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(KEYINPUT16), .B(G183gat), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n577_), .B(new_n578_), .Z(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT71), .B(KEYINPUT17), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G231gat), .A2(G233gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n446_), .B(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n512_), .A2(new_n517_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n586_), .A2(KEYINPUT69), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT70), .B(KEYINPUT17), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n588_), .B1(new_n586_), .B2(KEYINPUT69), .ZN(new_n589_));
  OAI221_X1 g388(.A(new_n580_), .B1(new_n581_), .B2(new_n585_), .C1(new_n587_), .C2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n581_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n579_), .B1(new_n585_), .B2(new_n591_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n575_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n548_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n596_), .B(new_n339_), .C1(new_n493_), .C2(new_n492_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT38), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n419_), .A2(new_n571_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT100), .ZN(new_n600_));
  INV_X1    g399(.A(new_n593_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT100), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n419_), .A2(new_n602_), .A3(new_n571_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n600_), .A2(new_n547_), .A3(new_n601_), .A4(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(G1gat), .B1(new_n604_), .B2(new_n410_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n598_), .A2(new_n605_), .ZN(G1324gat));
  NOR3_X1   g405(.A1(new_n595_), .A2(G8gat), .A3(new_n415_), .ZN(new_n607_));
  OAI21_X1  g406(.A(G8gat), .B1(new_n604_), .B2(new_n415_), .ZN(new_n608_));
  XOR2_X1   g407(.A(KEYINPUT101), .B(KEYINPUT39), .Z(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n609_), .ZN(new_n611_));
  OAI211_X1 g410(.A(G8gat), .B(new_n611_), .C1(new_n604_), .C2(new_n415_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n607_), .B1(new_n610_), .B2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT102), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n613_), .B(new_n615_), .Z(G1325gat));
  INV_X1    g415(.A(G15gat), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n596_), .A2(new_n617_), .A3(new_n374_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n604_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n617_), .B1(new_n619_), .B2(new_n374_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(KEYINPUT41), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n620_), .A2(KEYINPUT41), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n618_), .B1(new_n622_), .B2(new_n623_), .ZN(G1326gat));
  INV_X1    g423(.A(G22gat), .ZN(new_n625_));
  INV_X1    g424(.A(new_n408_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n596_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n625_), .B1(new_n619_), .B2(new_n626_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT42), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n628_), .A2(new_n629_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n627_), .B1(new_n631_), .B2(new_n632_), .ZN(G1327gat));
  NAND2_X1  g432(.A1(new_n547_), .A2(new_n593_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT43), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n636_), .B1(new_n575_), .B2(KEYINPUT104), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n638_), .B1(new_n419_), .B2(new_n575_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n575_), .ZN(new_n640_));
  AOI211_X1 g439(.A(new_n640_), .B(new_n637_), .C1(new_n409_), .C2(new_n418_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n635_), .B1(new_n639_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT44), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  OAI211_X1 g443(.A(KEYINPUT44), .B(new_n635_), .C1(new_n639_), .C2(new_n641_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n644_), .A2(new_n339_), .A3(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT105), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n644_), .A2(KEYINPUT105), .A3(new_n339_), .A4(new_n645_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n648_), .A2(G29gat), .A3(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n571_), .B1(new_n409_), .B2(new_n418_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n651_), .A2(new_n635_), .ZN(new_n652_));
  INV_X1    g451(.A(G29gat), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(new_n653_), .A3(new_n339_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n650_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT106), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n650_), .A2(new_n657_), .A3(new_n654_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(G1328gat));
  INV_X1    g458(.A(new_n415_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n644_), .A2(new_n660_), .A3(new_n645_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(G36gat), .ZN(new_n662_));
  INV_X1    g461(.A(G36gat), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n651_), .A2(new_n663_), .A3(new_n660_), .A4(new_n635_), .ZN(new_n664_));
  XOR2_X1   g463(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n665_));
  XOR2_X1   g464(.A(new_n664_), .B(new_n665_), .Z(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n662_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT46), .ZN(new_n669_));
  AOI21_X1  g468(.A(KEYINPUT108), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n666_), .B1(new_n661_), .B2(G36gat), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT108), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n671_), .A2(new_n672_), .A3(KEYINPUT46), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n671_), .A2(KEYINPUT109), .A3(KEYINPUT46), .ZN(new_n674_));
  AOI21_X1  g473(.A(KEYINPUT109), .B1(new_n671_), .B2(KEYINPUT46), .ZN(new_n675_));
  OAI22_X1  g474(.A1(new_n670_), .A2(new_n673_), .B1(new_n674_), .B2(new_n675_), .ZN(G1329gat));
  NAND2_X1  g475(.A1(new_n644_), .A2(new_n645_), .ZN(new_n677_));
  OAI21_X1  g476(.A(G43gat), .B1(new_n677_), .B2(new_n375_), .ZN(new_n678_));
  INV_X1    g477(.A(G43gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n652_), .A2(new_n679_), .A3(new_n374_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT47), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n681_), .B(new_n682_), .ZN(G1330gat));
  OAI21_X1  g482(.A(G50gat), .B1(new_n677_), .B2(new_n408_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n652_), .A2(new_n388_), .A3(new_n626_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1331gat));
  AND2_X1   g485(.A1(new_n600_), .A2(new_n603_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n687_), .A2(new_n601_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n546_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n689_), .A2(new_n480_), .ZN(new_n690_));
  AND4_X1   g489(.A1(G57gat), .A2(new_n688_), .A3(new_n339_), .A4(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n594_), .A2(new_n481_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT110), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n693_), .A2(new_n419_), .A3(new_n546_), .ZN(new_n694_));
  AOI21_X1  g493(.A(G57gat), .B1(new_n694_), .B2(new_n339_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n691_), .A2(new_n695_), .ZN(G1332gat));
  NAND3_X1  g495(.A1(new_n694_), .A2(new_n435_), .A3(new_n660_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n688_), .A2(new_n660_), .A3(new_n690_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(KEYINPUT111), .B(KEYINPUT48), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n698_), .A2(G64gat), .A3(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n699_), .B1(new_n698_), .B2(G64gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n697_), .B1(new_n701_), .B2(new_n702_), .ZN(G1333gat));
  INV_X1    g502(.A(G71gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n694_), .A2(new_n704_), .A3(new_n374_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n688_), .A2(new_n374_), .A3(new_n690_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT49), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n706_), .A2(new_n707_), .A3(G71gat), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n707_), .B1(new_n706_), .B2(G71gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n705_), .B1(new_n709_), .B2(new_n710_), .ZN(G1334gat));
  INV_X1    g510(.A(G78gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n694_), .A2(new_n712_), .A3(new_n626_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n688_), .A2(new_n626_), .A3(new_n690_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT50), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n714_), .A2(new_n715_), .A3(G78gat), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n715_), .B1(new_n714_), .B2(G78gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n713_), .B1(new_n717_), .B2(new_n718_), .ZN(G1335gat));
  NOR3_X1   g518(.A1(new_n601_), .A2(new_n689_), .A3(new_n480_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n651_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(G85gat), .B1(new_n722_), .B2(new_n339_), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n639_), .A2(new_n641_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n724_), .A2(new_n720_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n410_), .A2(new_n324_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n723_), .B1(new_n725_), .B2(new_n726_), .ZN(G1336gat));
  NOR3_X1   g526(.A1(new_n721_), .A2(G92gat), .A3(new_n415_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n725_), .A2(new_n660_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(G92gat), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT112), .Z(G1337gat));
  NAND2_X1  g530(.A1(new_n725_), .A2(new_n374_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(G99gat), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n722_), .B(new_n374_), .C1(new_n428_), .C2(new_n429_), .ZN(new_n734_));
  AOI211_X1 g533(.A(KEYINPUT113), .B(KEYINPUT51), .C1(new_n733_), .C2(new_n734_), .ZN(new_n735_));
  OR2_X1    g534(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n736_));
  NAND2_X1  g535(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n737_));
  AND4_X1   g536(.A1(new_n736_), .A2(new_n733_), .A3(new_n737_), .A4(new_n734_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n735_), .A2(new_n738_), .ZN(G1338gat));
  NAND3_X1  g538(.A1(new_n722_), .A2(new_n426_), .A3(new_n626_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n724_), .A2(new_n626_), .A3(new_n720_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT52), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n741_), .A2(new_n742_), .A3(G106gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n741_), .B2(G106gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g545(.A1(new_n415_), .A2(new_n339_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(new_n416_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n473_), .A2(new_n478_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n508_), .A2(new_n518_), .A3(new_n530_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n530_), .B1(new_n508_), .B2(new_n521_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n752_), .A2(new_n753_), .A3(new_n527_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n754_), .B1(new_n528_), .B2(new_n536_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT115), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT55), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n756_), .B(new_n757_), .C1(new_n472_), .C2(new_n420_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n446_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n549_), .A2(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n760_), .A2(KEYINPUT12), .A3(new_n463_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT12), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n468_), .A2(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n420_), .B1(new_n761_), .B2(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(KEYINPUT115), .B1(new_n764_), .B2(KEYINPUT55), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n472_), .A2(new_n420_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(KEYINPUT55), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n758_), .A2(new_n765_), .A3(new_n766_), .A4(new_n767_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n768_), .A2(KEYINPUT56), .A3(new_n478_), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT56), .B1(new_n768_), .B2(new_n478_), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n751_), .B(new_n755_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT58), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n768_), .A2(new_n478_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT56), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n768_), .A2(KEYINPUT56), .A3(new_n478_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n778_), .A2(KEYINPUT58), .A3(new_n751_), .A4(new_n755_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n773_), .A2(new_n779_), .A3(new_n575_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n571_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n776_), .A2(new_n782_), .A3(new_n777_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n768_), .A2(KEYINPUT116), .A3(KEYINPUT56), .A4(new_n478_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT73), .B1(new_n523_), .B2(new_n527_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n535_), .A2(new_n529_), .A3(new_n526_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n540_), .B1(new_n535_), .B2(new_n526_), .ZN(new_n787_));
  AOI211_X1 g586(.A(KEYINPUT72), .B(new_n527_), .C1(new_n533_), .C2(new_n534_), .ZN(new_n788_));
  OAI22_X1  g587(.A1(new_n785_), .A2(new_n786_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT74), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n537_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n750_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n783_), .A2(new_n784_), .A3(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n479_), .A2(new_n755_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n781_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n780_), .B1(new_n795_), .B2(KEYINPUT57), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n769_), .A2(new_n770_), .A3(KEYINPUT116), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n784_), .B(new_n751_), .C1(new_n544_), .C2(new_n545_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n794_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n571_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT57), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(KEYINPUT117), .B1(new_n796_), .B2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT57), .B1(new_n799_), .B2(new_n571_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n795_), .A2(KEYINPUT57), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT117), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n805_), .A2(new_n806_), .A3(new_n807_), .A4(new_n780_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n803_), .A2(new_n593_), .A3(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n594_), .A2(new_n810_), .A3(new_n546_), .A4(new_n480_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n594_), .A2(new_n546_), .A3(new_n480_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT54), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n811_), .A2(new_n812_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n813_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n749_), .B1(new_n809_), .B2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(G113gat), .B1(new_n818_), .B2(new_n689_), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n773_), .A2(new_n779_), .A3(new_n575_), .ZN(new_n820_));
  OAI21_X1  g619(.A(KEYINPUT119), .B1(new_n804_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n822_), .B(new_n780_), .C1(new_n795_), .C2(KEYINPUT57), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n821_), .A2(new_n806_), .A3(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT120), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n824_), .A2(new_n825_), .A3(new_n593_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n825_), .B1(new_n824_), .B2(new_n593_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT59), .B1(new_n828_), .B2(new_n817_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n749_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n809_), .A2(new_n817_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n830_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(KEYINPUT118), .A3(KEYINPUT59), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT59), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n818_), .B2(new_n835_), .ZN(new_n836_));
  AOI22_X1  g635(.A1(new_n829_), .A2(new_n830_), .B1(new_n833_), .B2(new_n836_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n689_), .A2(G113gat), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n819_), .B1(new_n837_), .B2(new_n838_), .ZN(G1340gat));
  INV_X1    g638(.A(KEYINPUT121), .ZN(new_n840_));
  INV_X1    g639(.A(G120gat), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n841_), .B1(new_n837_), .B2(new_n481_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n841_), .A2(KEYINPUT60), .ZN(new_n843_));
  AOI21_X1  g642(.A(KEYINPUT60), .B1(new_n481_), .B2(new_n841_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n832_), .A2(new_n843_), .A3(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n840_), .B1(new_n842_), .B2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n833_), .A2(new_n836_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n827_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n824_), .A2(new_n825_), .A3(new_n593_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n817_), .A3(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n850_), .A2(new_n835_), .A3(new_n830_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n847_), .A2(new_n481_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(G120gat), .ZN(new_n853_));
  INV_X1    g652(.A(new_n845_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(KEYINPUT121), .A3(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n846_), .A2(new_n855_), .ZN(G1341gat));
  AOI21_X1  g655(.A(G127gat), .B1(new_n818_), .B2(new_n601_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n601_), .A2(G127gat), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n857_), .B1(new_n837_), .B2(new_n858_), .ZN(G1342gat));
  INV_X1    g658(.A(G134gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n832_), .B2(new_n571_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(KEYINPUT122), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n640_), .A2(new_n860_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n862_), .B1(new_n837_), .B2(new_n863_), .ZN(G1343gat));
  AND2_X1   g663(.A1(new_n831_), .A2(new_n417_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n865_), .A2(new_n748_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n689_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n481_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g669(.A1(new_n866_), .A2(new_n601_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(KEYINPUT61), .B(G155gat), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(G1346gat));
  AOI21_X1  g672(.A(G162gat), .B1(new_n866_), .B2(new_n781_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n575_), .A2(G162gat), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n866_), .B2(new_n875_), .ZN(G1347gat));
  NOR2_X1   g675(.A1(new_n415_), .A2(new_n339_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n374_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(KEYINPUT123), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(new_n626_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n850_), .A2(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(G169gat), .B1(new_n881_), .B2(new_n546_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n881_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n885_), .A2(new_n689_), .A3(new_n225_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n882_), .A2(new_n883_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n884_), .A2(new_n886_), .A3(new_n887_), .ZN(G1348gat));
  AOI21_X1  g687(.A(G176gat), .B1(new_n885_), .B2(new_n481_), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n880_), .A2(new_n831_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n480_), .A2(new_n226_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n889_), .B1(new_n890_), .B2(new_n891_), .ZN(G1349gat));
  NOR3_X1   g691(.A1(new_n881_), .A2(new_n593_), .A3(new_n219_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n890_), .A2(new_n601_), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n894_), .B(KEYINPUT125), .Z(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n895_), .B2(new_n210_), .ZN(G1350gat));
  OAI21_X1  g695(.A(G190gat), .B1(new_n881_), .B2(new_n640_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n781_), .A2(new_n262_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n881_), .B2(new_n898_), .ZN(G1351gat));
  NAND2_X1  g698(.A1(new_n865_), .A2(new_n877_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n900_), .A2(new_n546_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(new_n234_), .ZN(G1352gat));
  NOR2_X1   g701(.A1(new_n900_), .A2(new_n480_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT126), .B(G204gat), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1353gat));
  INV_X1    g704(.A(new_n900_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n601_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n908_));
  AND2_X1   g707(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n907_), .A2(new_n908_), .A3(new_n909_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n910_), .B1(new_n907_), .B2(new_n908_), .ZN(G1354gat));
  NAND3_X1  g710(.A1(new_n906_), .A2(KEYINPUT127), .A3(new_n781_), .ZN(new_n912_));
  INV_X1    g711(.A(G218gat), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT127), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n914_), .B1(new_n900_), .B2(new_n571_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n912_), .A2(new_n913_), .A3(new_n915_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n906_), .A2(G218gat), .A3(new_n575_), .ZN(new_n917_));
  AND2_X1   g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1355gat));
endmodule


