//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 1 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n644_, new_n645_, new_n646_, new_n647_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n827_, new_n828_, new_n829_, new_n831_, new_n832_, new_n834_,
    new_n835_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n874_, new_n875_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT22), .B(G169gat), .ZN(new_n203_));
  INV_X1    g002(.A(G176gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n207_), .A2(KEYINPUT95), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT23), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n210_), .B1(G183gat), .B2(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n207_), .A2(KEYINPUT95), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n208_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G169gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(new_n204_), .A3(KEYINPUT79), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT79), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n216_), .B1(G169gat), .B2(G176gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT24), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n210_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n219_), .B1(G169gat), .B2(G176gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(new_n215_), .A3(new_n217_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT26), .B(G190gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT94), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT25), .B(G183gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n222_), .B(new_n224_), .C1(new_n226_), .C2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n213_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G211gat), .B(G218gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT90), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G197gat), .B(G204gat), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT21), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n232_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n233_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n232_), .A2(KEYINPUT21), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n230_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT20), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G226gat), .A2(G233gat), .ZN(new_n243_));
  XOR2_X1   g042(.A(new_n243_), .B(KEYINPUT92), .Z(new_n244_));
  XOR2_X1   g043(.A(new_n244_), .B(KEYINPUT19), .Z(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n211_), .A2(new_n206_), .A3(new_n205_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n224_), .A2(KEYINPUT80), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT80), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n223_), .A2(new_n250_), .A3(new_n215_), .A4(new_n217_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n227_), .A2(new_n225_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n249_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT81), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n221_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n249_), .A2(KEYINPUT81), .A3(new_n251_), .A4(new_n252_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n248_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n239_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n242_), .B(new_n246_), .C1(new_n257_), .C2(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n241_), .B1(new_n230_), .B2(new_n239_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n257_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n245_), .B(KEYINPUT93), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G8gat), .B(G36gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT18), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(G64gat), .ZN(new_n267_));
  INV_X1    g066(.A(G92gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n259_), .A2(new_n264_), .A3(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n269_), .B1(new_n259_), .B2(new_n264_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n202_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n270_), .A2(new_n202_), .ZN(new_n273_));
  OR2_X1    g072(.A1(new_n262_), .A2(new_n263_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n242_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n275_));
  AOI22_X1  g074(.A1(new_n274_), .A2(KEYINPUT98), .B1(new_n275_), .B2(new_n245_), .ZN(new_n276_));
  OR3_X1    g075(.A1(new_n262_), .A2(KEYINPUT98), .A3(new_n263_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n269_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n272_), .B1(new_n273_), .B2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G57gat), .B(G85gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G1gat), .B(G29gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n282_), .B(new_n283_), .Z(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT4), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G127gat), .B(G134gat), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n287_), .B(KEYINPUT83), .Z(new_n288_));
  XNOR2_X1  g087(.A(G113gat), .B(G120gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n287_), .B(KEYINPUT83), .ZN(new_n291_));
  INV_X1    g090(.A(new_n289_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n290_), .A2(new_n293_), .A3(KEYINPUT84), .ZN(new_n294_));
  OR3_X1    g093(.A1(new_n291_), .A2(KEYINPUT84), .A3(new_n292_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(G155gat), .B(G162gat), .Z(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n298_), .A2(KEYINPUT1), .ZN(new_n299_));
  NOR2_X1   g098(.A1(G141gat), .A2(G148gat), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G141gat), .A2(G148gat), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n301_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n299_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n300_), .B(KEYINPUT3), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n303_), .B(KEYINPUT2), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT87), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n307_), .A2(KEYINPUT87), .A3(new_n308_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n311_), .A2(new_n297_), .A3(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n306_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n296_), .A2(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n298_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n305_), .B1(new_n316_), .B2(new_n312_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n290_), .A2(new_n293_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n286_), .B1(new_n315_), .B2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G225gat), .A2(G233gat), .ZN(new_n321_));
  AOI21_X1  g120(.A(KEYINPUT4), .B1(new_n296_), .B2(new_n314_), .ZN(new_n322_));
  NOR3_X1   g121(.A1(new_n320_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n315_), .A2(new_n319_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(new_n321_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n285_), .B1(new_n323_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n324_), .A2(KEYINPUT4), .ZN(new_n328_));
  INV_X1    g127(.A(new_n321_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n322_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n328_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n331_), .A2(new_n284_), .A3(new_n325_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n327_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT99), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT99), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n327_), .A2(new_n332_), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n279_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT30), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n255_), .A2(new_n256_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n339_), .B1(new_n340_), .B2(new_n248_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n257_), .A2(KEYINPUT30), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n341_), .A2(KEYINPUT82), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT82), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n257_), .A2(KEYINPUT30), .ZN(new_n345_));
  AOI211_X1 g144(.A(new_n339_), .B(new_n248_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n344_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  XOR2_X1   g146(.A(G15gat), .B(G43gat), .Z(new_n348_));
  NAND2_X1  g147(.A1(G227gat), .A2(G233gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G71gat), .B(G99gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n343_), .A2(new_n347_), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n352_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n341_), .A2(KEYINPUT82), .A3(new_n342_), .A4(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT85), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT86), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT86), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n353_), .A2(new_n359_), .A3(new_n355_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n296_), .B(KEYINPUT31), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n358_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n361_), .ZN(new_n363_));
  OAI211_X1 g162(.A(KEYINPUT86), .B(new_n363_), .C1(new_n356_), .C2(new_n357_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n258_), .B1(KEYINPUT29), .B2(new_n314_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT89), .ZN(new_n367_));
  AOI22_X1  g166(.A1(new_n239_), .A2(new_n367_), .B1(G228gat), .B2(G233gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n366_), .B(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(G22gat), .B(G50gat), .Z(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT28), .B1(new_n314_), .B2(KEYINPUT29), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT28), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT29), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n317_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT88), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n371_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n375_), .B1(new_n371_), .B2(new_n374_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n370_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n371_), .A2(new_n374_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT88), .ZN(new_n380_));
  INV_X1    g179(.A(new_n370_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n371_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G78gat), .B(G106gat), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n385_), .A2(KEYINPUT91), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n378_), .A2(new_n383_), .A3(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n385_), .B1(new_n378_), .B2(new_n383_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n369_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n369_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n378_), .A2(new_n383_), .A3(new_n386_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n378_), .A2(new_n383_), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n390_), .B(new_n391_), .C1(new_n392_), .C2(new_n385_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n389_), .A2(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n365_), .A2(new_n394_), .ZN(new_n395_));
  AOI22_X1  g194(.A1(new_n362_), .A2(new_n364_), .B1(new_n389_), .B2(new_n393_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n338_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n284_), .B1(new_n324_), .B2(new_n321_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n328_), .A2(new_n330_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n398_), .B1(new_n399_), .B2(new_n321_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT33), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n400_), .B1(new_n327_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT97), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n403_), .B1(new_n327_), .B2(new_n401_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n284_), .B1(new_n331_), .B2(new_n325_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n405_), .A2(KEYINPUT97), .A3(KEYINPUT33), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n270_), .A2(new_n271_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n402_), .A2(new_n404_), .A3(new_n406_), .A4(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n269_), .A2(KEYINPUT32), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n259_), .A2(new_n264_), .A3(new_n409_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n276_), .A2(new_n277_), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n333_), .B(new_n410_), .C1(new_n411_), .C2(new_n409_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n408_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n394_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(new_n365_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n397_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G57gat), .B(G64gat), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n417_), .A2(KEYINPUT11), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(KEYINPUT11), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G71gat), .B(G78gat), .ZN(new_n420_));
  OR3_X1    g219(.A1(new_n418_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n417_), .A2(new_n420_), .A3(KEYINPUT11), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT12), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT69), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT65), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n427_), .A2(G92gat), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n268_), .A2(KEYINPUT65), .ZN(new_n429_));
  OAI21_X1  g228(.A(G85gat), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n431_));
  INV_X1    g230(.A(G85gat), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n432_), .A2(new_n268_), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n430_), .A2(new_n431_), .B1(KEYINPUT9), .B2(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(KEYINPUT64), .A2(G106gat), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  OR2_X1    g235(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(KEYINPUT64), .A2(G106gat), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .A4(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT6), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT66), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT66), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT6), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G99gat), .A2(G106gat), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n442_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n445_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n440_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT67), .B1(new_n434_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n445_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n443_), .A2(KEYINPUT6), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n441_), .A2(KEYINPUT66), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n450_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n442_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n454_));
  XOR2_X1   g253(.A(KEYINPUT10), .B(G99gat), .Z(new_n455_));
  INV_X1    g254(.A(new_n439_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n456_), .A2(new_n435_), .ZN(new_n457_));
  AOI22_X1  g256(.A1(new_n453_), .A2(new_n454_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT67), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n433_), .A2(KEYINPUT9), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n268_), .A2(KEYINPUT65), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n427_), .A2(G92gat), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n432_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n431_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n460_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n458_), .A2(new_n459_), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n449_), .A2(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(G99gat), .A2(G106gat), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT7), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n470_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G85gat), .B(G92gat), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT8), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT8), .ZN(new_n474_));
  INV_X1    g273(.A(new_n472_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n453_), .A2(new_n454_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n474_), .B(new_n475_), .C1(new_n477_), .C2(new_n470_), .ZN(new_n478_));
  AOI22_X1  g277(.A1(new_n467_), .A2(KEYINPUT68), .B1(new_n473_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT68), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n449_), .A2(new_n480_), .A3(new_n466_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n426_), .B1(new_n479_), .B2(new_n481_), .ZN(new_n482_));
  AND4_X1   g281(.A1(new_n459_), .A2(new_n465_), .A3(new_n476_), .A4(new_n440_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n459_), .B1(new_n458_), .B2(new_n465_), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT68), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n473_), .A2(new_n478_), .ZN(new_n486_));
  AND4_X1   g285(.A1(new_n426_), .A2(new_n485_), .A3(new_n481_), .A4(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n425_), .B1(new_n482_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n467_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(new_n486_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n490_), .A2(new_n422_), .A3(new_n421_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(new_n424_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n489_), .A2(new_n486_), .A3(new_n423_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G230gat), .A2(G233gat), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n488_), .A2(new_n492_), .A3(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n491_), .A2(new_n493_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n494_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n496_), .A2(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(G120gat), .B(G148gat), .Z(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(G204gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(KEYINPUT5), .B(G176gat), .ZN(new_n503_));
  XOR2_X1   g302(.A(new_n502_), .B(new_n503_), .Z(new_n504_));
  OR2_X1    g303(.A1(new_n500_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n500_), .A2(new_n504_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT13), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n505_), .A2(KEYINPUT13), .A3(new_n506_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(G29gat), .B(G36gat), .Z(new_n512_));
  XOR2_X1   g311(.A(G43gat), .B(G50gat), .Z(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G29gat), .B(G36gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G43gat), .B(G50gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT15), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G15gat), .B(G22gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G1gat), .A2(G8gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT14), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G1gat), .B(G8gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n519_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT76), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n525_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n518_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G229gat), .A2(G233gat), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n528_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n518_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n525_), .B(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n531_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n532_), .A2(new_n536_), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n537_), .A2(KEYINPUT77), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G113gat), .B(G141gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(G169gat), .ZN(new_n540_));
  INV_X1    g339(.A(G197gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n542_), .B1(new_n537_), .B2(KEYINPUT77), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n532_), .A2(new_n536_), .A3(new_n542_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n544_), .A2(KEYINPUT78), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(KEYINPUT78), .ZN(new_n546_));
  AOI22_X1  g345(.A1(new_n538_), .A2(new_n543_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n511_), .A2(new_n547_), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n416_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT72), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n550_), .A2(KEYINPUT37), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(KEYINPUT37), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G232gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT34), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT35), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  OAI22_X1  g356(.A1(new_n490_), .A2(new_n533_), .B1(KEYINPUT35), .B2(new_n554_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n519_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n485_), .A2(new_n481_), .A3(new_n486_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT69), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n479_), .A2(new_n426_), .A3(new_n481_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n560_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n559_), .B1(new_n564_), .B2(KEYINPUT70), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n519_), .B1(new_n482_), .B2(new_n487_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT70), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n557_), .B1(new_n565_), .B2(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(G190gat), .B(G218gat), .Z(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT71), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(G134gat), .ZN(new_n572_));
  INV_X1    g371(.A(G162gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT36), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n558_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n557_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n564_), .A2(KEYINPUT70), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n577_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n569_), .A2(new_n576_), .A3(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n574_), .B(KEYINPUT36), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n583_), .B1(new_n569_), .B2(new_n580_), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n551_), .B(new_n552_), .C1(new_n581_), .C2(new_n584_), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n565_), .A2(new_n568_), .A3(new_n557_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n578_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n582_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n569_), .A2(new_n580_), .A3(new_n576_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n588_), .A2(new_n550_), .A3(KEYINPUT37), .A4(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n585_), .A2(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(G183gat), .B(G211gat), .Z(new_n592_));
  XNOR2_X1  g391(.A(G127gat), .B(G155gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(KEYINPUT73), .B(KEYINPUT16), .Z(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n596_), .A2(KEYINPUT17), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(KEYINPUT17), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n423_), .B(new_n529_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  AOI211_X1 g400(.A(new_n597_), .B(new_n598_), .C1(new_n601_), .C2(KEYINPUT75), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n602_), .B1(KEYINPUT75), .B2(new_n601_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n597_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT74), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n603_), .A2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n591_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n549_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n337_), .ZN(new_n610_));
  OR3_X1    g409(.A1(new_n609_), .A2(G1gat), .A3(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT101), .ZN(new_n614_));
  INV_X1    g413(.A(new_n607_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n548_), .A2(KEYINPUT102), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n588_), .A2(new_n589_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n618_), .B1(new_n397_), .B2(new_n415_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT102), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n620_), .B1(new_n511_), .B2(new_n547_), .ZN(new_n621_));
  AND4_X1   g420(.A1(new_n615_), .A2(new_n616_), .A3(new_n619_), .A4(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(new_n337_), .ZN(new_n623_));
  AOI22_X1  g422(.A1(new_n611_), .A2(new_n612_), .B1(G1gat), .B2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n614_), .A2(new_n624_), .ZN(G1324gat));
  INV_X1    g424(.A(new_n279_), .ZN(new_n626_));
  OR3_X1    g425(.A1(new_n609_), .A2(G8gat), .A3(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n622_), .A2(new_n279_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(G8gat), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n629_), .A2(KEYINPUT39), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(KEYINPUT39), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n627_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT40), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n633_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(G1325gat));
  INV_X1    g435(.A(G15gat), .ZN(new_n637_));
  INV_X1    g436(.A(new_n365_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n622_), .B2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT41), .ZN(new_n640_));
  INV_X1    g439(.A(new_n609_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n641_), .A2(new_n637_), .A3(new_n638_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(G1326gat));
  INV_X1    g442(.A(G22gat), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n622_), .B2(new_n394_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT42), .Z(new_n646_));
  NAND3_X1  g445(.A1(new_n641_), .A2(new_n644_), .A3(new_n394_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(G1327gat));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n585_), .A2(KEYINPUT103), .A3(new_n590_), .ZN(new_n650_));
  AOI21_X1  g449(.A(KEYINPUT103), .B1(new_n585_), .B2(new_n590_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n416_), .A2(new_n650_), .A3(new_n652_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n585_), .A2(new_n590_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n654_), .A2(KEYINPUT43), .ZN(new_n655_));
  AOI22_X1  g454(.A1(new_n653_), .A2(KEYINPUT43), .B1(new_n416_), .B2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n616_), .A2(new_n607_), .A3(new_n621_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n649_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n616_), .A2(new_n607_), .A3(new_n621_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT43), .ZN(new_n660_));
  INV_X1    g459(.A(new_n650_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n661_), .A2(new_n651_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n660_), .B1(new_n662_), .B2(new_n416_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n655_), .A2(new_n416_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n659_), .B(KEYINPUT44), .C1(new_n663_), .C2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n658_), .A2(new_n666_), .A3(new_n337_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT104), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT104), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n658_), .A2(new_n666_), .A3(new_n669_), .A4(new_n337_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n668_), .A2(G29gat), .A3(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n617_), .A2(new_n615_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT105), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n549_), .A2(new_n673_), .ZN(new_n674_));
  OR3_X1    g473(.A1(new_n674_), .A2(G29gat), .A3(new_n610_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n671_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT106), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n671_), .A2(new_n678_), .A3(new_n675_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(G1328gat));
  NOR3_X1   g479(.A1(new_n674_), .A2(G36gat), .A3(new_n626_), .ZN(new_n681_));
  XOR2_X1   g480(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n682_));
  XOR2_X1   g481(.A(new_n681_), .B(new_n682_), .Z(new_n683_));
  NAND3_X1  g482(.A1(new_n658_), .A2(new_n666_), .A3(new_n279_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(G36gat), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT46), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(G1329gat));
  AND2_X1   g487(.A1(new_n658_), .A2(new_n666_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(G43gat), .A3(new_n638_), .ZN(new_n690_));
  INV_X1    g489(.A(G43gat), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n691_), .B1(new_n674_), .B2(new_n365_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g493(.A(G50gat), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n414_), .A2(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n549_), .A2(new_n394_), .A3(new_n673_), .ZN(new_n697_));
  AOI22_X1  g496(.A1(new_n689_), .A2(new_n696_), .B1(new_n695_), .B2(new_n697_), .ZN(G1331gat));
  AND2_X1   g497(.A1(new_n509_), .A2(new_n510_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n538_), .A2(new_n543_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n545_), .A2(new_n546_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n699_), .A2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n619_), .A2(new_n703_), .A3(new_n615_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G57gat), .B1(new_n704_), .B2(new_n610_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n703_), .A2(new_n416_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(new_n608_), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n610_), .A2(G57gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n705_), .B1(new_n707_), .B2(new_n708_), .ZN(G1332gat));
  OAI21_X1  g508(.A(G64gat), .B1(new_n704_), .B2(new_n626_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT48), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n626_), .A2(G64gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n711_), .B1(new_n707_), .B2(new_n712_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT108), .Z(G1333gat));
  OAI21_X1  g513(.A(G71gat), .B1(new_n704_), .B2(new_n365_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT49), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n365_), .A2(G71gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n707_), .B2(new_n717_), .ZN(G1334gat));
  OAI21_X1  g517(.A(G78gat), .B1(new_n704_), .B2(new_n414_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT50), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n414_), .A2(G78gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n720_), .B1(new_n707_), .B2(new_n721_), .ZN(G1335gat));
  INV_X1    g521(.A(KEYINPUT109), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n703_), .A2(new_n607_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n723_), .B1(new_n656_), .B2(new_n724_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n699_), .A2(new_n615_), .A3(new_n702_), .ZN(new_n726_));
  OAI211_X1 g525(.A(KEYINPUT109), .B(new_n726_), .C1(new_n663_), .C2(new_n665_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G85gat), .B1(new_n729_), .B2(new_n610_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n706_), .A2(new_n673_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n731_), .A2(new_n432_), .A3(new_n337_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(G1336gat));
  AOI21_X1  g532(.A(G92gat), .B1(new_n731_), .B2(new_n279_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n626_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n728_), .B2(new_n735_), .ZN(G1337gat));
  INV_X1    g535(.A(G99gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n728_), .B2(new_n638_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n731_), .A2(new_n455_), .A3(new_n638_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT110), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n739_), .A2(KEYINPUT111), .A3(new_n741_), .A4(KEYINPUT51), .ZN(new_n742_));
  NAND2_X1  g541(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n743_));
  OR2_X1    g542(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n740_), .B(new_n745_), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n743_), .B(new_n744_), .C1(new_n746_), .C2(new_n738_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n742_), .A2(new_n747_), .ZN(G1338gat));
  XOR2_X1   g547(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n749_));
  OAI211_X1 g548(.A(new_n394_), .B(new_n726_), .C1(new_n663_), .C2(new_n665_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n750_), .B2(G106gat), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT113), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n750_), .A2(G106gat), .A3(new_n749_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n394_), .A2(new_n457_), .ZN(new_n756_));
  AOI22_X1  g555(.A1(new_n751_), .A2(new_n752_), .B1(new_n731_), .B2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT53), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT53), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n755_), .A2(new_n760_), .A3(new_n757_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1339gat));
  AOI21_X1  g561(.A(new_n547_), .B1(new_n500_), .B2(new_n504_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n488_), .A2(new_n493_), .A3(new_n492_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n498_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n496_), .A2(new_n766_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n488_), .A2(KEYINPUT55), .A3(new_n492_), .A4(new_n495_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n765_), .A2(new_n767_), .A3(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT114), .ZN(new_n770_));
  INV_X1    g569(.A(new_n504_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n765_), .A2(new_n767_), .A3(new_n772_), .A4(new_n768_), .ZN(new_n773_));
  AND4_X1   g572(.A1(KEYINPUT56), .A2(new_n770_), .A3(new_n771_), .A4(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n504_), .B1(new_n769_), .B2(KEYINPUT114), .ZN(new_n775_));
  AOI21_X1  g574(.A(KEYINPUT56), .B1(new_n775_), .B2(new_n773_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n763_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n528_), .A2(new_n530_), .A3(new_n535_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n542_), .B1(new_n534_), .B2(new_n531_), .ZN(new_n779_));
  AOI22_X1  g578(.A1(new_n545_), .A2(new_n546_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n507_), .A2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n618_), .B1(new_n777_), .B2(new_n781_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n780_), .A2(new_n506_), .ZN(new_n783_));
  OAI211_X1 g582(.A(KEYINPUT58), .B(new_n783_), .C1(new_n774_), .C2(new_n776_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n591_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n770_), .A2(new_n771_), .A3(new_n773_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT56), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n775_), .A2(KEYINPUT56), .A3(new_n773_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT58), .B1(new_n790_), .B2(new_n783_), .ZN(new_n791_));
  OAI22_X1  g590(.A1(new_n782_), .A2(KEYINPUT57), .B1(new_n785_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT57), .ZN(new_n793_));
  AOI211_X1 g592(.A(new_n793_), .B(new_n618_), .C1(new_n777_), .C2(new_n781_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n607_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n608_), .A2(new_n699_), .A3(new_n547_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT54), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n395_), .A2(new_n337_), .A3(new_n626_), .ZN(new_n799_));
  XOR2_X1   g598(.A(new_n799_), .B(KEYINPUT115), .Z(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(G113gat), .B1(new_n802_), .B2(new_n702_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(KEYINPUT59), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT59), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n798_), .A2(new_n805_), .A3(new_n800_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n804_), .A2(new_n806_), .ZN(new_n807_));
  XOR2_X1   g606(.A(KEYINPUT116), .B(G113gat), .Z(new_n808_));
  NAND2_X1  g607(.A1(new_n702_), .A2(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT117), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n803_), .B1(new_n807_), .B2(new_n810_), .ZN(G1340gat));
  INV_X1    g610(.A(KEYINPUT60), .ZN(new_n812_));
  XOR2_X1   g611(.A(KEYINPUT118), .B(G120gat), .Z(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n812_), .B1(new_n699_), .B2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n699_), .B1(new_n802_), .B2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n802_), .A2(new_n812_), .A3(new_n815_), .ZN(new_n817_));
  AOI22_X1  g616(.A1(new_n807_), .A2(new_n816_), .B1(new_n817_), .B2(new_n813_), .ZN(G1341gat));
  INV_X1    g617(.A(KEYINPUT119), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n615_), .A2(G127gat), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n804_), .A2(new_n819_), .A3(new_n806_), .A4(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(G127gat), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n821_), .A2(KEYINPUT119), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n802_), .B(new_n615_), .C1(new_n805_), .C2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(G1342gat));
  NAND3_X1  g625(.A1(new_n804_), .A2(new_n591_), .A3(new_n806_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(G134gat), .ZN(new_n828_));
  OR2_X1    g627(.A1(new_n617_), .A2(G134gat), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n801_), .B2(new_n829_), .ZN(G1343gat));
  AND4_X1   g629(.A1(new_n396_), .A2(new_n798_), .A3(new_n337_), .A4(new_n626_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n702_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n511_), .ZN(new_n834_));
  XOR2_X1   g633(.A(KEYINPUT120), .B(G148gat), .Z(new_n835_));
  XNOR2_X1  g634(.A(new_n834_), .B(new_n835_), .ZN(G1345gat));
  NAND2_X1  g635(.A1(new_n831_), .A2(new_n615_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(KEYINPUT61), .B(G155gat), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(KEYINPUT121), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n837_), .B(new_n839_), .ZN(G1346gat));
  AOI21_X1  g639(.A(G162gat), .B1(new_n831_), .B2(new_n618_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n661_), .A2(new_n573_), .A3(new_n651_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n841_), .B1(new_n831_), .B2(new_n842_), .ZN(G1347gat));
  NOR2_X1   g642(.A1(new_n626_), .A2(new_n337_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n638_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n845_), .A2(new_n394_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n847_), .B1(new_n795_), .B2(new_n797_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n848_), .A2(new_n702_), .A3(new_n203_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n214_), .B1(new_n848_), .B2(new_n702_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(KEYINPUT62), .ZN(new_n851_));
  AOI211_X1 g650(.A(new_n547_), .B(new_n847_), .C1(new_n795_), .C2(new_n797_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT62), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n852_), .A2(new_n853_), .A3(new_n214_), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT122), .B1(new_n851_), .B2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n850_), .A2(KEYINPUT62), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n853_), .B1(new_n852_), .B2(new_n214_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n856_), .A2(new_n857_), .A3(new_n858_), .A4(new_n849_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n855_), .A2(new_n859_), .ZN(G1348gat));
  AOI21_X1  g659(.A(G176gat), .B1(new_n848_), .B2(new_n511_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n394_), .B1(new_n795_), .B2(new_n797_), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n862_), .A2(KEYINPUT123), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(KEYINPUT123), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n845_), .A2(new_n699_), .A3(new_n204_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n861_), .B1(new_n865_), .B2(new_n866_), .ZN(G1349gat));
  INV_X1    g666(.A(new_n848_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n868_), .A2(new_n607_), .A3(new_n227_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n845_), .A2(new_n607_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n863_), .A2(new_n864_), .A3(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(G183gat), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n869_), .B1(new_n871_), .B2(new_n872_), .ZN(G1350gat));
  OAI21_X1  g672(.A(G190gat), .B1(new_n868_), .B2(new_n654_), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n617_), .A2(new_n226_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n868_), .B2(new_n875_), .ZN(G1351gat));
  NAND4_X1  g675(.A1(new_n798_), .A2(new_n702_), .A3(new_n396_), .A4(new_n844_), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n877_), .A2(KEYINPUT124), .A3(new_n541_), .ZN(new_n878_));
  AOI21_X1  g677(.A(KEYINPUT124), .B1(new_n877_), .B2(new_n541_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n877_), .A2(new_n541_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n878_), .A2(new_n879_), .A3(new_n880_), .ZN(G1352gat));
  NAND2_X1  g680(.A1(new_n798_), .A2(new_n396_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n844_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n511_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g685(.A(KEYINPUT125), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n882_), .A2(new_n607_), .A3(new_n883_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n887_), .B1(new_n888_), .B2(new_n890_), .ZN(new_n891_));
  AOI211_X1 g690(.A(new_n638_), .B(new_n414_), .C1(new_n795_), .C2(new_n797_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n844_), .ZN(new_n893_));
  OAI211_X1 g692(.A(KEYINPUT125), .B(new_n889_), .C1(new_n893_), .C2(new_n607_), .ZN(new_n894_));
  XOR2_X1   g693(.A(KEYINPUT63), .B(G211gat), .Z(new_n895_));
  AOI22_X1  g694(.A1(new_n891_), .A2(new_n894_), .B1(new_n888_), .B2(new_n895_), .ZN(G1354gat));
  NAND3_X1  g695(.A1(new_n892_), .A2(new_n618_), .A3(new_n844_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT126), .ZN(new_n898_));
  AOI21_X1  g697(.A(G218gat), .B1(new_n897_), .B2(new_n898_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n884_), .A2(KEYINPUT126), .A3(new_n618_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n591_), .A2(G218gat), .ZN(new_n901_));
  XOR2_X1   g700(.A(new_n901_), .B(KEYINPUT127), .Z(new_n902_));
  AOI22_X1  g701(.A1(new_n899_), .A2(new_n900_), .B1(new_n884_), .B2(new_n902_), .ZN(G1355gat));
endmodule


