//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 0 0 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n844_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n871_, new_n872_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_;
  XOR2_X1   g000(.A(G113gat), .B(G120gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G127gat), .B(G134gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  AND3_X1   g003(.A1(KEYINPUT85), .A2(G141gat), .A3(G148gat), .ZN(new_n205_));
  AOI21_X1  g004(.A(KEYINPUT85), .B1(G141gat), .B2(G148gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT87), .B1(new_n207_), .B2(KEYINPUT2), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT87), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n209_), .B(new_n210_), .C1(new_n205_), .C2(new_n206_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT88), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND4_X1  g013(.A1(KEYINPUT88), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n215_));
  INV_X1    g014(.A(G141gat), .ZN(new_n216_));
  INV_X1    g015(.A(G148gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(new_n217_), .A3(KEYINPUT3), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n219_), .B1(G141gat), .B2(G148gat), .ZN(new_n220_));
  AOI22_X1  g019(.A1(new_n214_), .A2(new_n215_), .B1(new_n218_), .B2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n208_), .A2(new_n211_), .A3(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G155gat), .A2(G162gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n222_), .A2(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n207_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n225_), .B1(KEYINPUT1), .B2(new_n223_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT86), .ZN(new_n230_));
  OAI22_X1  g029(.A1(new_n229_), .A2(new_n230_), .B1(KEYINPUT1), .B2(new_n223_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n229_), .A2(new_n230_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n228_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n227_), .A2(KEYINPUT89), .A3(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT89), .B1(new_n227_), .B2(new_n233_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n204_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT98), .B1(new_n236_), .B2(KEYINPUT4), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n227_), .A2(new_n233_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n238_), .A2(new_n204_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n236_), .A2(KEYINPUT4), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT89), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n227_), .A2(KEYINPUT89), .A3(new_n233_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT98), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n244_), .A2(new_n245_), .A3(new_n246_), .A4(new_n204_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G225gat), .A2(G233gat), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n237_), .A2(new_n240_), .A3(new_n247_), .A4(new_n249_), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n236_), .A2(new_n239_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n248_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G1gat), .B(G29gat), .ZN(new_n253_));
  INV_X1    g052(.A(G85gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT0), .B(G57gat), .ZN(new_n256_));
  XOR2_X1   g055(.A(new_n255_), .B(new_n256_), .Z(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n250_), .A2(new_n252_), .A3(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n259_), .A2(KEYINPUT99), .A3(KEYINPUT33), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT99), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n250_), .A2(new_n252_), .A3(new_n258_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT33), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n261_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G8gat), .B(G36gat), .ZN(new_n265_));
  INV_X1    g064(.A(G92gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT18), .B(G64gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G226gat), .A2(G233gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT20), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G183gat), .A2(G190gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT23), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(G183gat), .B2(G190gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT22), .B(G169gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT97), .ZN(new_n283_));
  XOR2_X1   g082(.A(KEYINPUT83), .B(G176gat), .Z(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n281_), .A2(new_n285_), .ZN(new_n286_));
  OR3_X1    g085(.A1(KEYINPUT82), .A2(G169gat), .A3(G176gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(KEYINPUT82), .B1(G169gat), .B2(G176gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT26), .B(G190gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT25), .B(G183gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  AND3_X1   g094(.A1(new_n292_), .A2(new_n277_), .A3(new_n295_), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n287_), .A2(new_n288_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n297_), .A2(new_n279_), .A3(new_n290_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n286_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G211gat), .B(G218gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT92), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT21), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G197gat), .B(G204gat), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT93), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n303_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n302_), .B(new_n307_), .C1(new_n306_), .C2(new_n305_), .ZN(new_n308_));
  INV_X1    g107(.A(G197gat), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n309_), .A2(G204gat), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT21), .B1(new_n310_), .B2(KEYINPUT91), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n311_), .A2(new_n304_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n304_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n312_), .A2(new_n301_), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n308_), .A2(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n275_), .B1(new_n300_), .B2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n297_), .A2(KEYINPUT24), .A3(new_n279_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT24), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n289_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(G183gat), .ZN(new_n320_));
  OR3_X1    g119(.A1(new_n320_), .A2(KEYINPUT81), .A3(KEYINPUT25), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT25), .B1(new_n320_), .B2(KEYINPUT81), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n321_), .A2(new_n293_), .A3(new_n322_), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n317_), .A2(new_n319_), .A3(new_n277_), .A4(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n284_), .A2(new_n282_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n278_), .A2(new_n279_), .A3(new_n325_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n308_), .A2(new_n324_), .A3(new_n314_), .A4(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n274_), .B1(new_n316_), .B2(new_n327_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n286_), .A2(new_n299_), .A3(new_n314_), .A4(new_n308_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n324_), .A2(new_n326_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n315_), .A2(new_n330_), .ZN(new_n331_));
  AND4_X1   g130(.A1(KEYINPUT20), .A2(new_n329_), .A3(new_n331_), .A4(new_n274_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n270_), .B1(new_n328_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n315_), .ZN(new_n334_));
  AOI22_X1  g133(.A1(new_n281_), .A2(new_n285_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n275_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n336_), .A2(new_n274_), .A3(new_n331_), .ZN(new_n337_));
  OAI211_X1 g136(.A(KEYINPUT20), .B(new_n327_), .C1(new_n334_), .C2(new_n335_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(new_n273_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n339_), .A3(new_n269_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n333_), .A2(new_n340_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n237_), .A2(new_n240_), .A3(new_n247_), .A4(new_n248_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n258_), .B1(new_n251_), .B2(new_n249_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n341_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n262_), .A2(new_n263_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n260_), .A2(new_n264_), .A3(new_n344_), .A4(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n269_), .A2(KEYINPUT32), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NOR3_X1   g147(.A1(new_n328_), .A2(new_n332_), .A3(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n336_), .A2(new_n331_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n273_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n351_), .B1(new_n273_), .B2(new_n338_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n349_), .B1(new_n352_), .B2(new_n348_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n258_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n353_), .B1(new_n259_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT100), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n353_), .B(KEYINPUT100), .C1(new_n259_), .C2(new_n354_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n346_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  XOR2_X1   g158(.A(G78gat), .B(G106gat), .Z(new_n360_));
  INV_X1    g159(.A(G228gat), .ZN(new_n361_));
  INV_X1    g160(.A(G233gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n238_), .A2(KEYINPUT29), .ZN(new_n363_));
  AOI211_X1 g162(.A(new_n361_), .B(new_n362_), .C1(new_n363_), .C2(new_n315_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n334_), .B1(G228gat), .B2(G233gat), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n234_), .A2(new_n235_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n366_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n360_), .B1(new_n365_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n365_), .A2(new_n369_), .A3(new_n360_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT94), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n370_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n376_), .B1(new_n244_), .B2(KEYINPUT29), .ZN(new_n377_));
  INV_X1    g176(.A(new_n376_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n367_), .A2(new_n368_), .A3(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G22gat), .B(G50gat), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n377_), .A2(new_n379_), .A3(new_n381_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n373_), .B1(new_n375_), .B2(new_n385_), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n383_), .A2(new_n384_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n387_), .A2(new_n374_), .A3(new_n372_), .A4(new_n371_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT101), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n391_), .B1(new_n259_), .B2(new_n354_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n354_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n393_), .A2(KEYINPUT101), .A3(new_n262_), .ZN(new_n394_));
  AOI22_X1  g193(.A1(new_n392_), .A2(new_n394_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n352_), .A2(new_n270_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n396_), .A2(KEYINPUT27), .A3(new_n340_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT27), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n341_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  AOI22_X1  g200(.A1(new_n359_), .A2(new_n390_), .B1(new_n395_), .B2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n330_), .B(KEYINPUT30), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT84), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n403_), .B(new_n404_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G71gat), .B(G99gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G227gat), .A2(G233gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(G15gat), .B(G43gat), .Z(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  MUX2_X1   g210(.A(new_n405_), .B(new_n406_), .S(new_n411_), .Z(new_n412_));
  XOR2_X1   g211(.A(new_n204_), .B(KEYINPUT31), .Z(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n390_), .A2(new_n401_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n394_), .A2(new_n392_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  OAI22_X1  g216(.A1(new_n402_), .A2(new_n414_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G229gat), .A2(G233gat), .ZN(new_n419_));
  XOR2_X1   g218(.A(G1gat), .B(G8gat), .Z(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G15gat), .B(G22gat), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT75), .ZN(new_n423_));
  INV_X1    g222(.A(G1gat), .ZN(new_n424_));
  INV_X1    g223(.A(G8gat), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT14), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n422_), .A2(new_n423_), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n423_), .B1(new_n422_), .B2(new_n426_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n421_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n429_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n431_), .A2(new_n427_), .A3(new_n420_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G29gat), .B(G36gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G43gat), .B(G50gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n433_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n430_), .A2(new_n432_), .A3(new_n436_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT79), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n438_), .A2(KEYINPUT79), .A3(new_n439_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n419_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n436_), .B(KEYINPUT15), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n433_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(new_n419_), .A3(new_n439_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT80), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT80), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n447_), .A2(new_n450_), .A3(new_n419_), .A4(new_n439_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G113gat), .B(G141gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G169gat), .B(G197gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n445_), .A2(new_n449_), .A3(new_n451_), .A4(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n449_), .A2(new_n451_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n454_), .B1(new_n457_), .B2(new_n444_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n418_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT102), .ZN(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G127gat), .B(G155gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  XOR2_X1   g263(.A(G183gat), .B(G211gat), .Z(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G231gat), .A2(G233gat), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n430_), .A2(new_n432_), .A3(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n467_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G57gat), .B(G64gat), .ZN(new_n470_));
  OR2_X1    g269(.A1(new_n470_), .A2(KEYINPUT11), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(KEYINPUT11), .ZN(new_n472_));
  XOR2_X1   g271(.A(G71gat), .B(G78gat), .Z(new_n473_));
  NAND3_X1  g272(.A1(new_n471_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  OR2_X1    g273(.A1(new_n472_), .A2(new_n473_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  OR3_X1    g275(.A1(new_n468_), .A2(new_n469_), .A3(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n476_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n466_), .B1(new_n479_), .B2(KEYINPUT17), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n466_), .A2(KEYINPUT17), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n477_), .A2(KEYINPUT77), .A3(new_n478_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT13), .ZN(new_n485_));
  XOR2_X1   g284(.A(G176gat), .B(G204gat), .Z(new_n486_));
  XNOR2_X1  g285(.A(G120gat), .B(G148gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n488_), .B(new_n489_), .Z(new_n490_));
  NAND2_X1  g289(.A1(new_n254_), .A2(new_n266_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT9), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G85gat), .A2(G92gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n491_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n493_), .A2(KEYINPUT64), .A3(new_n492_), .ZN(new_n495_));
  AOI21_X1  g294(.A(KEYINPUT64), .B1(new_n493_), .B2(new_n492_), .ZN(new_n496_));
  NOR3_X1   g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  AND3_X1   g296(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n498_));
  AOI21_X1  g297(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT10), .B(G99gat), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n500_), .B1(G106gat), .B2(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n497_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(G99gat), .ZN(new_n505_));
  INV_X1    g304(.A(G106gat), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(new_n506_), .A3(KEYINPUT66), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n507_), .A2(KEYINPUT65), .A3(KEYINPUT7), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT65), .ZN(new_n509_));
  NOR2_X1   g308(.A1(G99gat), .A2(G106gat), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n509_), .B1(new_n510_), .B2(KEYINPUT66), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT7), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n512_), .B1(new_n510_), .B2(new_n509_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n508_), .B(new_n500_), .C1(new_n511_), .C2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT8), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n491_), .A2(new_n493_), .ZN(new_n516_));
  AND3_X1   g315(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n515_), .B1(new_n514_), .B2(new_n516_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n504_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n476_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n504_), .B(new_n476_), .C1(new_n517_), .C2(new_n518_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(G230gat), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n523_), .A2(new_n524_), .A3(new_n362_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n362_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n521_), .A2(KEYINPUT12), .A3(new_n522_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT12), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n519_), .A2(new_n528_), .A3(new_n520_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n526_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n490_), .B1(new_n525_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NOR3_X1   g331(.A1(new_n525_), .A2(new_n530_), .A3(new_n490_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n485_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n533_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n535_), .A2(KEYINPUT13), .A3(new_n531_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n484_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT74), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n436_), .B(new_n504_), .C1(new_n517_), .C2(new_n518_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n514_), .A2(new_n516_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT8), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n503_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT15), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n436_), .B(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n539_), .B1(new_n543_), .B2(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(KEYINPUT68), .B(KEYINPUT34), .Z(new_n547_));
  NAND2_X1  g346(.A1(G232gat), .A2(G233gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT35), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n546_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT69), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT69), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n546_), .A2(new_n554_), .A3(new_n551_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n549_), .B(KEYINPUT35), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n539_), .B(new_n556_), .C1(new_n543_), .C2(new_n545_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT70), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n519_), .A2(new_n446_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n560_), .A2(KEYINPUT70), .A3(new_n539_), .A4(new_n556_), .ZN(new_n561_));
  AOI22_X1  g360(.A1(new_n553_), .A2(new_n555_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(G190gat), .B(G218gat), .Z(new_n563_));
  XOR2_X1   g362(.A(G134gat), .B(G162gat), .Z(new_n564_));
  XOR2_X1   g363(.A(new_n563_), .B(new_n564_), .Z(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT36), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT72), .B1(new_n562_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT72), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n546_), .A2(new_n554_), .A3(new_n551_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n554_), .B1(new_n546_), .B2(new_n551_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n559_), .A2(new_n561_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n569_), .B(new_n566_), .C1(new_n572_), .C2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n565_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n575_), .A2(KEYINPUT36), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n562_), .A2(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(KEYINPUT73), .B(KEYINPUT37), .Z(new_n578_));
  NAND4_X1  g377(.A1(new_n568_), .A2(new_n574_), .A3(new_n577_), .A4(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n553_), .A2(new_n555_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n559_), .A2(new_n561_), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n580_), .A2(new_n581_), .A3(new_n576_), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n566_), .B(KEYINPUT71), .Z(new_n583_));
  AOI21_X1  g382(.A(new_n583_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n584_));
  OAI21_X1  g383(.A(KEYINPUT37), .B1(new_n582_), .B2(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n538_), .B1(new_n579_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n579_), .A2(new_n538_), .A3(new_n585_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n537_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n589_), .B(KEYINPUT78), .Z(new_n590_));
  AND2_X1   g389(.A1(new_n461_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n416_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n591_), .A2(new_n424_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT38), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n568_), .A2(new_n577_), .A3(new_n574_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n534_), .A2(new_n536_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n598_), .A2(new_n459_), .A3(new_n484_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n596_), .B1(new_n599_), .B2(KEYINPUT103), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n600_), .B1(KEYINPUT103), .B2(new_n599_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(new_n418_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n602_), .A2(KEYINPUT104), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(KEYINPUT104), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(G1gat), .B1(new_n605_), .B2(new_n416_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n593_), .A2(new_n594_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n595_), .A2(new_n606_), .A3(new_n607_), .ZN(G1324gat));
  NAND3_X1  g407(.A1(new_n591_), .A2(new_n425_), .A3(new_n400_), .ZN(new_n609_));
  OAI21_X1  g408(.A(G8gat), .B1(new_n602_), .B2(new_n401_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT39), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(G1325gat));
  INV_X1    g413(.A(new_n414_), .ZN(new_n615_));
  OAI21_X1  g414(.A(G15gat), .B1(new_n605_), .B2(new_n615_), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n616_), .A2(KEYINPUT41), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(KEYINPUT41), .ZN(new_n618_));
  INV_X1    g417(.A(G15gat), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n591_), .A2(new_n619_), .A3(new_n414_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n617_), .A2(new_n618_), .A3(new_n620_), .ZN(G1326gat));
  INV_X1    g420(.A(G22gat), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n591_), .A2(new_n622_), .A3(new_n389_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT42), .ZN(new_n624_));
  INV_X1    g423(.A(new_n605_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(new_n389_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n624_), .B1(new_n626_), .B2(G22gat), .ZN(new_n627_));
  AOI211_X1 g426(.A(KEYINPUT42), .B(new_n622_), .C1(new_n625_), .C2(new_n389_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n623_), .B1(new_n627_), .B2(new_n628_), .ZN(G1327gat));
  NOR3_X1   g428(.A1(new_n597_), .A2(new_n596_), .A3(new_n484_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n461_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(G29gat), .B1(new_n632_), .B2(new_n592_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n415_), .A2(new_n417_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n359_), .A2(new_n390_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n395_), .A2(new_n401_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n634_), .B1(new_n637_), .B2(new_n615_), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n579_), .A2(new_n538_), .A3(new_n585_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n639_), .A2(new_n586_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(KEYINPUT43), .B1(new_n638_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT43), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n418_), .A2(new_n643_), .A3(new_n640_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n459_), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n597_), .A2(new_n646_), .A3(new_n484_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n648_), .A2(new_n649_), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n652_), .A2(G29gat), .A3(new_n592_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n633_), .B1(new_n651_), .B2(new_n653_), .ZN(G1328gat));
  NOR2_X1   g453(.A1(new_n401_), .A2(G36gat), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n461_), .A2(new_n630_), .A3(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT45), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n652_), .A2(new_n400_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G36gat), .B1(new_n658_), .B2(new_n650_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT107), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n657_), .A2(new_n659_), .A3(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n661_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1329gat));
  NAND3_X1  g463(.A1(new_n652_), .A2(G43gat), .A3(new_n414_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n631_), .A2(new_n615_), .ZN(new_n666_));
  OAI22_X1  g465(.A1(new_n665_), .A2(new_n650_), .B1(new_n666_), .B2(G43gat), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g467(.A(G50gat), .B1(new_n632_), .B2(new_n389_), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n652_), .A2(G50gat), .A3(new_n389_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n669_), .B1(new_n651_), .B2(new_n670_), .ZN(G1331gat));
  INV_X1    g470(.A(new_n484_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n598_), .A2(new_n459_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n638_), .A2(new_n672_), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(new_n596_), .ZN(new_n676_));
  INV_X1    g475(.A(G57gat), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n676_), .A2(new_n677_), .A3(new_n416_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n679_), .A2(KEYINPUT108), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n675_), .A2(new_n641_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n677_), .B1(new_n681_), .B2(new_n416_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n679_), .A2(KEYINPUT108), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n680_), .A2(new_n682_), .A3(new_n683_), .ZN(G1332gat));
  OR3_X1    g483(.A1(new_n681_), .A2(G64gat), .A3(new_n401_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n675_), .A2(new_n400_), .A3(new_n596_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n686_), .A2(G64gat), .A3(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n687_), .B1(new_n686_), .B2(G64gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n685_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT110), .Z(G1333gat));
  OAI21_X1  g491(.A(G71gat), .B1(new_n676_), .B2(new_n615_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT49), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n615_), .A2(G71gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n694_), .B1(new_n681_), .B2(new_n695_), .ZN(G1334gat));
  OAI21_X1  g495(.A(G78gat), .B1(new_n676_), .B2(new_n390_), .ZN(new_n697_));
  XOR2_X1   g496(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n390_), .A2(G78gat), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n699_), .B1(new_n681_), .B2(new_n700_), .ZN(G1335gat));
  NOR2_X1   g500(.A1(new_n638_), .A2(new_n674_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n484_), .A2(new_n596_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT112), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n702_), .A2(KEYINPUT112), .A3(new_n703_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(G85gat), .B1(new_n708_), .B2(new_n592_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n674_), .A2(new_n484_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n645_), .A2(new_n710_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n416_), .A2(new_n254_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n709_), .B1(new_n711_), .B2(new_n712_), .ZN(G1336gat));
  AOI21_X1  g512(.A(G92gat), .B1(new_n708_), .B2(new_n400_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n400_), .A2(G92gat), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT113), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n714_), .B1(new_n711_), .B2(new_n716_), .ZN(G1337gat));
  INV_X1    g516(.A(KEYINPUT51), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT115), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n645_), .A2(new_n414_), .A3(new_n710_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(G99gat), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT114), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n718_), .A2(KEYINPUT115), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n615_), .A2(new_n501_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n708_), .B2(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n719_), .B1(new_n722_), .B2(new_n725_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n721_), .A2(KEYINPUT114), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT114), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n720_), .B2(G99gat), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n725_), .B(new_n719_), .C1(new_n727_), .C2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n726_), .A2(new_n731_), .ZN(G1338gat));
  XNOR2_X1  g531(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT118), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n418_), .A2(new_n643_), .A3(new_n640_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n643_), .B1(new_n418_), .B2(new_n640_), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n389_), .B(new_n710_), .C1(new_n735_), .C2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT116), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT116), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n645_), .A2(new_n739_), .A3(new_n389_), .A4(new_n710_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n738_), .A2(G106gat), .A3(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT52), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT52), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n738_), .A2(new_n740_), .A3(new_n743_), .A4(G106gat), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(new_n745_));
  AOI211_X1 g544(.A(G106gat), .B(new_n390_), .C1(new_n706_), .C2(new_n707_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n734_), .B1(new_n745_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n734_), .ZN(new_n749_));
  AOI211_X1 g548(.A(new_n746_), .B(new_n749_), .C1(new_n742_), .C2(new_n744_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n748_), .A2(new_n750_), .ZN(G1339gat));
  INV_X1    g550(.A(KEYINPUT125), .ZN(new_n752_));
  INV_X1    g551(.A(new_n537_), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n753_), .B(new_n646_), .C1(new_n639_), .C2(new_n586_), .ZN(new_n754_));
  XOR2_X1   g553(.A(KEYINPUT119), .B(KEYINPUT54), .Z(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT121), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT120), .ZN(new_n759_));
  INV_X1    g558(.A(new_n755_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n589_), .A2(new_n759_), .A3(new_n646_), .A4(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT120), .B1(new_n754_), .B2(new_n755_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n754_), .A2(KEYINPUT121), .A3(new_n755_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n758_), .A2(new_n761_), .A3(new_n762_), .A4(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n419_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n447_), .A2(new_n765_), .A3(new_n439_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(new_n454_), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n766_), .A2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n535_), .A2(new_n456_), .A3(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT55), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n771_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n526_), .A2(KEYINPUT122), .ZN(new_n773_));
  OAI22_X1  g572(.A1(KEYINPUT55), .A2(new_n530_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n772_), .A2(new_n773_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n490_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT56), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  OAI211_X1 g577(.A(KEYINPUT56), .B(new_n490_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n770_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n780_), .A2(KEYINPUT58), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(KEYINPUT58), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(new_n640_), .A3(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n459_), .A2(new_n535_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n784_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n456_), .A2(new_n769_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n786_), .B1(new_n531_), .B2(new_n535_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n596_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT57), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  OAI211_X1 g589(.A(KEYINPUT57), .B(new_n596_), .C1(new_n785_), .C2(new_n787_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n783_), .A2(new_n790_), .A3(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(new_n672_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n764_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT59), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n390_), .A2(new_n401_), .A3(new_n414_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n796_), .A2(new_n416_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n794_), .A2(new_n795_), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n764_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n791_), .A2(KEYINPUT123), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT58), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n780_), .B(new_n801_), .ZN(new_n802_));
  AOI22_X1  g601(.A1(new_n800_), .A2(new_n790_), .B1(new_n802_), .B2(new_n640_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n788_), .A2(KEYINPUT123), .A3(new_n789_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n484_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n797_), .B1(new_n799_), .B2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT124), .B1(new_n806_), .B2(KEYINPUT59), .ZN(new_n807_));
  INV_X1    g606(.A(new_n797_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n800_), .A2(new_n790_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n809_), .A2(new_n804_), .A3(new_n783_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n672_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n808_), .B1(new_n811_), .B2(new_n764_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT124), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n812_), .A2(new_n813_), .A3(new_n795_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n459_), .B(new_n798_), .C1(new_n807_), .C2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(G113gat), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n806_), .A2(G113gat), .A3(new_n646_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n752_), .B1(new_n816_), .B2(new_n818_), .ZN(new_n819_));
  AOI211_X1 g618(.A(KEYINPUT125), .B(new_n817_), .C1(new_n815_), .C2(G113gat), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(G1340gat));
  INV_X1    g620(.A(G120gat), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n822_), .B1(new_n598_), .B2(KEYINPUT60), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n812_), .B(new_n823_), .C1(KEYINPUT60), .C2(new_n822_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n807_), .A2(new_n814_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n798_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n825_), .A2(new_n598_), .A3(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n824_), .B1(new_n827_), .B2(new_n822_), .ZN(G1341gat));
  NOR2_X1   g627(.A1(new_n764_), .A2(new_n672_), .ZN(new_n829_));
  INV_X1    g628(.A(G127gat), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n797_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n825_), .A2(new_n672_), .A3(new_n826_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(new_n830_), .ZN(G1342gat));
  INV_X1    g632(.A(new_n596_), .ZN(new_n834_));
  AOI21_X1  g633(.A(G134gat), .B1(new_n812_), .B2(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n825_), .A2(new_n826_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n640_), .A2(G134gat), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n835_), .B1(new_n836_), .B2(new_n837_), .ZN(G1343gat));
  AOI21_X1  g637(.A(new_n414_), .B1(new_n811_), .B2(new_n764_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n390_), .A2(new_n416_), .A3(new_n400_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(new_n646_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(new_n216_), .ZN(G1344gat));
  NOR2_X1   g642(.A1(new_n841_), .A2(new_n598_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(new_n217_), .ZN(G1345gat));
  NOR2_X1   g644(.A1(new_n841_), .A2(new_n672_), .ZN(new_n846_));
  XOR2_X1   g645(.A(KEYINPUT61), .B(G155gat), .Z(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(G1346gat));
  INV_X1    g647(.A(new_n841_), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n849_), .A2(G162gat), .A3(new_n640_), .ZN(new_n850_));
  AOI21_X1  g649(.A(G162gat), .B1(new_n849_), .B2(new_n834_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1347gat));
  INV_X1    g651(.A(KEYINPUT62), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n417_), .A2(new_n389_), .A3(new_n401_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n794_), .A2(new_n854_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n855_), .A2(new_n646_), .ZN(new_n856_));
  INV_X1    g655(.A(G169gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n853_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  OAI211_X1 g657(.A(KEYINPUT62), .B(G169gat), .C1(new_n855_), .C2(new_n646_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n856_), .A2(new_n283_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n858_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  XOR2_X1   g660(.A(new_n861_), .B(KEYINPUT126), .Z(G1348gat));
  NAND3_X1  g661(.A1(new_n854_), .A2(G176gat), .A3(new_n597_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n863_), .B1(new_n811_), .B2(new_n764_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n855_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n597_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n864_), .B1(new_n866_), .B2(new_n284_), .ZN(G1349gat));
  AOI21_X1  g666(.A(G183gat), .B1(new_n829_), .B2(new_n854_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n672_), .A2(new_n294_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n865_), .B2(new_n869_), .ZN(G1350gat));
  OAI21_X1  g669(.A(G190gat), .B1(new_n855_), .B2(new_n641_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n834_), .A2(new_n293_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n855_), .B2(new_n872_), .ZN(G1351gat));
  AND2_X1   g672(.A1(new_n395_), .A2(new_n400_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n839_), .A2(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n646_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(new_n309_), .ZN(G1352gat));
  INV_X1    g676(.A(new_n875_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n597_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g679(.A(KEYINPUT63), .ZN(new_n881_));
  INV_X1    g680(.A(G211gat), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n484_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  XOR2_X1   g682(.A(new_n883_), .B(KEYINPUT127), .Z(new_n884_));
  NAND2_X1  g683(.A1(new_n878_), .A2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n881_), .A2(new_n882_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n885_), .B(new_n886_), .ZN(G1354gat));
  AND3_X1   g686(.A1(new_n878_), .A2(G218gat), .A3(new_n640_), .ZN(new_n888_));
  AOI21_X1  g687(.A(G218gat), .B1(new_n878_), .B2(new_n834_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n888_), .A2(new_n889_), .ZN(G1355gat));
endmodule


