//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 0 0 0 1 1 0 1 0 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n632_, new_n633_, new_n634_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n848_, new_n849_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n891_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT25), .B(G183gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT26), .B(G190gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  OR2_X1    g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n206_), .A2(KEYINPUT24), .A3(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n205_), .A2(new_n208_), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n209_), .A2(KEYINPUT81), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT82), .B(KEYINPUT23), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT83), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT83), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n211_), .A2(new_n215_), .A3(new_n212_), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n214_), .B(new_n216_), .C1(KEYINPUT23), .C2(new_n212_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n209_), .A2(KEYINPUT81), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n206_), .A2(KEYINPUT24), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n210_), .A2(new_n217_), .A3(new_n218_), .A4(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT22), .B(G169gat), .ZN(new_n222_));
  INV_X1    g021(.A(G176gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(new_n207_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n211_), .A2(new_n212_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n227_), .B1(KEYINPUT23), .B2(new_n212_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n226_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n221_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT84), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G71gat), .B(G99gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G227gat), .A2(G233gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n232_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT84), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n231_), .B(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n235_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G15gat), .B(G43gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT30), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n236_), .A2(new_n240_), .A3(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n242_), .B1(new_n236_), .B2(new_n240_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n202_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n236_), .A2(new_n240_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n242_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n236_), .A2(new_n240_), .A3(new_n242_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(KEYINPUT85), .A3(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G127gat), .B(G134gat), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n251_), .A2(G113gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(G113gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(G120gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n252_), .A2(G120gat), .A3(new_n253_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n258_), .B(KEYINPUT31), .Z(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n245_), .A2(new_n250_), .A3(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT0), .B(G57gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(G85gat), .ZN(new_n263_));
  XOR2_X1   g062(.A(G1gat), .B(G29gat), .Z(new_n264_));
  XOR2_X1   g063(.A(new_n263_), .B(new_n264_), .Z(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G225gat), .A2(G233gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G141gat), .A2(G148gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT2), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n270_));
  OR3_X1    g069(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT87), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G155gat), .B(G162gat), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT87), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n269_), .A2(new_n276_), .A3(new_n270_), .A4(new_n271_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n273_), .A2(new_n275_), .A3(new_n277_), .ZN(new_n278_));
  AND2_X1   g077(.A1(G155gat), .A2(G162gat), .ZN(new_n279_));
  AOI22_X1  g078(.A1(new_n279_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n280_));
  OAI221_X1 g079(.A(new_n280_), .B1(G141gat), .B2(G148gat), .C1(KEYINPUT1), .C2(new_n274_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(new_n258_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n283_), .A2(KEYINPUT4), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n278_), .A2(new_n281_), .A3(new_n257_), .A4(new_n256_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n283_), .A2(new_n286_), .A3(KEYINPUT4), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n267_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n267_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n289_), .B1(new_n283_), .B2(new_n286_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n266_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n287_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n289_), .B1(new_n292_), .B2(new_n284_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n290_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(new_n265_), .A3(new_n294_), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n291_), .A2(new_n295_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n248_), .A2(KEYINPUT85), .A3(new_n249_), .A4(new_n259_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n261_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G226gat), .A2(G233gat), .ZN(new_n299_));
  XOR2_X1   g098(.A(new_n299_), .B(KEYINPUT94), .Z(new_n300_));
  XOR2_X1   g099(.A(new_n300_), .B(KEYINPUT19), .Z(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n229_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n217_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n226_), .ZN(new_n305_));
  NOR3_X1   g104(.A1(new_n228_), .A2(new_n209_), .A3(new_n219_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT89), .B(G197gat), .ZN(new_n309_));
  INV_X1    g108(.A(G204gat), .ZN(new_n310_));
  OR3_X1    g109(.A1(new_n309_), .A2(KEYINPUT91), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT21), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(G197gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT91), .B1(new_n309_), .B2(new_n310_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n311_), .A2(new_n312_), .A3(new_n313_), .A4(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n310_), .A2(G197gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT90), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n309_), .A2(new_n310_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT21), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  XOR2_X1   g118(.A(G211gat), .B(G218gat), .Z(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n315_), .A2(new_n319_), .A3(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n311_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(KEYINPUT21), .A3(new_n320_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n308_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n221_), .A2(new_n230_), .A3(new_n322_), .A4(new_n324_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT20), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n302_), .B1(new_n327_), .B2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT18), .B(G64gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(G92gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G8gat), .B(G36gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n332_), .B(new_n333_), .Z(new_n334_));
  AOI21_X1  g133(.A(new_n306_), .B1(new_n226_), .B2(new_n304_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(new_n322_), .A3(new_n324_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n231_), .A2(new_n325_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n336_), .A2(new_n337_), .A3(KEYINPUT20), .A4(new_n301_), .ZN(new_n338_));
  AND3_X1   g137(.A1(new_n330_), .A2(new_n334_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n326_), .A2(new_n328_), .A3(KEYINPUT20), .A4(new_n301_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT97), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n328_), .A2(KEYINPUT20), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT97), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n343_), .A2(new_n344_), .A3(new_n301_), .A4(new_n326_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n342_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT96), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n308_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n335_), .A2(KEYINPUT96), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT92), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n322_), .A2(new_n350_), .A3(new_n324_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n350_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n348_), .B(new_n349_), .C1(new_n352_), .C2(new_n353_), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n337_), .A2(KEYINPUT20), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n301_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n346_), .A2(new_n356_), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n340_), .B(KEYINPUT27), .C1(new_n357_), .C2(new_n334_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n353_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n282_), .A2(KEYINPUT29), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n359_), .A2(new_n351_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(G228gat), .ZN(new_n362_));
  INV_X1    g161(.A(G233gat), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n361_), .A2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G78gat), .B(G106gat), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n366_), .B(KEYINPUT93), .Z(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n360_), .B(new_n325_), .C1(new_n362_), .C2(new_n363_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n365_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n368_), .B1(new_n365_), .B2(new_n369_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G22gat), .B(G50gat), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  XOR2_X1   g173(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n375_));
  OR3_X1    g174(.A1(new_n282_), .A2(KEYINPUT29), .A3(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n375_), .B1(new_n282_), .B2(KEYINPUT29), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n374_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n376_), .A2(new_n374_), .A3(new_n377_), .ZN(new_n379_));
  OAI22_X1  g178(.A1(new_n371_), .A2(new_n372_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n365_), .A2(new_n369_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n367_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n379_), .A2(new_n378_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(new_n383_), .A3(new_n370_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n380_), .A2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT98), .B(KEYINPUT27), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n334_), .B1(new_n330_), .B2(new_n338_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n386_), .B1(new_n339_), .B2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n358_), .A2(new_n385_), .A3(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n298_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n358_), .A2(new_n388_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n380_), .A2(new_n296_), .A3(new_n384_), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT99), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n380_), .A2(new_n296_), .A3(new_n384_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT99), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n394_), .A2(new_n395_), .A3(new_n388_), .A4(new_n358_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n285_), .A2(new_n267_), .A3(new_n287_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n283_), .A2(new_n286_), .A3(new_n289_), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n397_), .A2(new_n265_), .A3(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n265_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT33), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n339_), .A2(new_n387_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT33), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n291_), .A2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n401_), .A2(new_n402_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n334_), .A2(KEYINPUT32), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n407_), .B1(new_n346_), .B2(new_n356_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n291_), .A2(new_n295_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n330_), .A2(new_n338_), .A3(new_n406_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT95), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n330_), .A2(KEYINPUT95), .A3(new_n338_), .A4(new_n406_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n408_), .A2(new_n409_), .A3(new_n412_), .A4(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n405_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n385_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n393_), .A2(new_n396_), .A3(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT86), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n261_), .A2(new_n418_), .A3(new_n297_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n418_), .B1(new_n261_), .B2(new_n297_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n390_), .B1(new_n417_), .B2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G169gat), .B(G197gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT79), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(G113gat), .ZN(new_n425_));
  INV_X1    g224(.A(G141gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G29gat), .B(G36gat), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n429_), .A2(G43gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(G43gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(G50gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n430_), .A2(G50gat), .A3(new_n431_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(G1gat), .B(G8gat), .Z(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G15gat), .B(G22gat), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT74), .ZN(new_n440_));
  INV_X1    g239(.A(G1gat), .ZN(new_n441_));
  INV_X1    g240(.A(G8gat), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT14), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n439_), .A2(new_n440_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n440_), .B1(new_n439_), .B2(new_n443_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n438_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n446_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n448_), .A2(new_n437_), .A3(new_n444_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n436_), .A2(new_n450_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n430_), .A2(G50gat), .A3(new_n431_), .ZN(new_n452_));
  AOI21_X1  g251(.A(G50gat), .B1(new_n430_), .B2(new_n431_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT15), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT15), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n436_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n451_), .B1(new_n458_), .B2(new_n450_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G229gat), .A2(G233gat), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n460_), .B(KEYINPUT78), .Z(new_n461_));
  NAND3_X1  g260(.A1(new_n454_), .A2(new_n449_), .A3(new_n447_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n436_), .A2(new_n450_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n460_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n459_), .A2(new_n461_), .B1(new_n464_), .B2(KEYINPUT77), .ZN(new_n465_));
  OR2_X1    g264(.A1(new_n464_), .A2(KEYINPUT77), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n428_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n458_), .A2(new_n450_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(new_n462_), .A3(new_n461_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n464_), .A2(KEYINPUT77), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n466_), .A2(new_n469_), .A3(new_n470_), .A4(new_n428_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT80), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT80), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n465_), .A2(new_n466_), .A3(new_n473_), .A4(new_n428_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n467_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G57gat), .B(G64gat), .ZN(new_n476_));
  OR2_X1    g275(.A1(new_n476_), .A2(KEYINPUT11), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(KEYINPUT11), .ZN(new_n478_));
  XOR2_X1   g277(.A(G71gat), .B(G78gat), .Z(new_n479_));
  NAND3_X1  g278(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n478_), .A2(new_n479_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT6), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT64), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT64), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT6), .ZN(new_n487_));
  AND2_X1   g286(.A1(G99gat), .A2(G106gat), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n485_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n488_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT65), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n488_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n486_), .A2(KEYINPUT6), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n484_), .A2(KEYINPUT64), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n492_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT65), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n485_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(G99gat), .A2(G106gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT7), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n491_), .A2(new_n498_), .A3(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(G85gat), .B(G92gat), .Z(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT8), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n489_), .A2(new_n490_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n500_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT8), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(new_n507_), .A3(new_n502_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n504_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n502_), .A2(KEYINPUT9), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT9), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n511_), .A2(G85gat), .A3(G92gat), .ZN(new_n512_));
  XOR2_X1   g311(.A(KEYINPUT10), .B(G99gat), .Z(new_n513_));
  INV_X1    g312(.A(G106gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n505_), .A2(new_n510_), .A3(new_n512_), .A4(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT66), .B1(new_n509_), .B2(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n507_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n506_), .A2(new_n507_), .A3(new_n502_), .ZN(new_n519_));
  OAI211_X1 g318(.A(KEYINPUT66), .B(new_n516_), .C1(new_n518_), .C2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(KEYINPUT12), .B(new_n483_), .C1(new_n517_), .C2(new_n521_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n482_), .B(new_n516_), .C1(new_n518_), .C2(new_n519_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  AND2_X1   g323(.A1(G230gat), .A2(G233gat), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n516_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n527_));
  AOI21_X1  g326(.A(KEYINPUT12), .B1(new_n527_), .B2(new_n483_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n528_), .A2(KEYINPUT67), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT67), .ZN(new_n530_));
  AOI211_X1 g329(.A(new_n530_), .B(KEYINPUT12), .C1(new_n527_), .C2(new_n483_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n522_), .B(new_n526_), .C1(new_n529_), .C2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n482_), .B1(new_n509_), .B2(new_n516_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n525_), .B1(new_n533_), .B2(new_n524_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G120gat), .B(G148gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(new_n310_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT5), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(new_n223_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n532_), .A2(new_n534_), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n538_), .B1(new_n532_), .B2(new_n534_), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT13), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n541_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT13), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(new_n544_), .A3(new_n539_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NOR3_X1   g346(.A1(new_n422_), .A2(new_n475_), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT37), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n454_), .B(new_n516_), .C1(new_n518_), .C2(new_n519_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT66), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n527_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(new_n520_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n551_), .B1(new_n554_), .B2(new_n458_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT68), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G232gat), .A2(G233gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n557_), .A2(new_n561_), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n555_), .A2(KEYINPUT35), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n555_), .A2(new_n556_), .A3(new_n560_), .ZN(new_n564_));
  AND3_X1   g363(.A1(new_n562_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT69), .B(G190gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(G218gat), .ZN(new_n567_));
  XOR2_X1   g366(.A(G134gat), .B(G162gat), .Z(new_n568_));
  XOR2_X1   g367(.A(new_n567_), .B(new_n568_), .Z(new_n569_));
  XOR2_X1   g368(.A(new_n569_), .B(KEYINPUT36), .Z(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n549_), .B1(new_n565_), .B2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n562_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n573_));
  XOR2_X1   g372(.A(KEYINPUT70), .B(KEYINPUT36), .Z(new_n574_));
  NAND2_X1  g373(.A1(new_n569_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT71), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT72), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n573_), .A2(KEYINPUT72), .A3(new_n576_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n572_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n570_), .B1(new_n573_), .B2(KEYINPUT73), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT73), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n562_), .A2(new_n563_), .A3(new_n583_), .A4(new_n564_), .ZN(new_n584_));
  AOI22_X1  g383(.A1(new_n582_), .A2(new_n584_), .B1(new_n573_), .B2(new_n576_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n581_), .B1(new_n585_), .B2(KEYINPUT37), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G231gat), .A2(G233gat), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n588_), .B(KEYINPUT75), .Z(new_n589_));
  XNOR2_X1  g388(.A(new_n482_), .B(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n450_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT17), .ZN(new_n593_));
  XNOR2_X1  g392(.A(KEYINPUT16), .B(G183gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(G211gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G127gat), .B(G155gat), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n595_), .B(new_n596_), .Z(new_n597_));
  NOR3_X1   g396(.A1(new_n592_), .A2(new_n593_), .A3(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n593_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n598_), .B1(new_n592_), .B2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT76), .Z(new_n602_));
  NAND3_X1  g401(.A1(new_n548_), .A2(new_n587_), .A3(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT100), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n604_), .A2(G1gat), .A3(new_n296_), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n605_), .A2(KEYINPUT38), .ZN(new_n606_));
  INV_X1    g405(.A(new_n585_), .ZN(new_n607_));
  AND3_X1   g406(.A1(new_n548_), .A2(new_n601_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(G1gat), .B1(new_n609_), .B2(new_n296_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n605_), .A2(KEYINPUT38), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n606_), .A2(new_n610_), .A3(new_n611_), .ZN(G1324gat));
  INV_X1    g411(.A(new_n391_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G8gat), .B1(new_n609_), .B2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(KEYINPUT101), .B(KEYINPUT39), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n391_), .A2(new_n442_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n604_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n617_), .A2(KEYINPUT40), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT40), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n622_), .B1(new_n616_), .B2(new_n619_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(G1325gat));
  OAI21_X1  g423(.A(G15gat), .B1(new_n609_), .B2(new_n421_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT102), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT41), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n627_), .ZN(new_n629_));
  OR3_X1    g428(.A1(new_n603_), .A2(G15gat), .A3(new_n421_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n628_), .A2(new_n629_), .A3(new_n630_), .ZN(G1326gat));
  OAI21_X1  g430(.A(G22gat), .B1(new_n609_), .B2(new_n385_), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n632_), .B(KEYINPUT42), .Z(new_n633_));
  NOR3_X1   g432(.A1(new_n603_), .A2(G22gat), .A3(new_n385_), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n633_), .A2(new_n634_), .ZN(G1327gat));
  NOR2_X1   g434(.A1(new_n547_), .A2(new_n475_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n602_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT43), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT103), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n582_), .A2(new_n584_), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT37), .B1(new_n640_), .B2(new_n577_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n572_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n639_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n581_), .B(KEYINPUT103), .C1(new_n585_), .C2(KEYINPUT37), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n417_), .A2(new_n421_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n390_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n638_), .B1(new_n645_), .B2(new_n648_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n422_), .A2(new_n587_), .A3(KEYINPUT43), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n636_), .B(new_n637_), .C1(new_n649_), .C2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT44), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n648_), .A2(new_n638_), .A3(new_n586_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n422_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n654_), .B1(new_n655_), .B2(new_n638_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n656_), .A2(KEYINPUT44), .A3(new_n636_), .A4(new_n637_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n653_), .A2(new_n657_), .A3(new_n409_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT104), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n653_), .A2(new_n657_), .A3(KEYINPUT104), .A4(new_n409_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n660_), .A2(G29gat), .A3(new_n661_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n548_), .A2(new_n585_), .A3(new_n637_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n296_), .A2(G29gat), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT105), .Z(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n662_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT106), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n662_), .A2(KEYINPUT106), .A3(new_n666_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1328gat));
  INV_X1    g470(.A(G36gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n663_), .A2(new_n672_), .A3(new_n391_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT45), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n653_), .A2(new_n657_), .A3(new_n391_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n674_), .B1(new_n675_), .B2(new_n672_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT46), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n676_), .B(new_n677_), .ZN(G1329gat));
  INV_X1    g477(.A(KEYINPUT108), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n261_), .A2(new_n297_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n681_), .A2(G43gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n653_), .A2(new_n657_), .A3(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n421_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n663_), .A2(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(KEYINPUT107), .B(G43gat), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n679_), .B1(new_n683_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n683_), .A2(new_n679_), .A3(new_n687_), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT47), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n690_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT47), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n692_), .A2(new_n693_), .A3(new_n688_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n691_), .A2(new_n694_), .ZN(G1330gat));
  INV_X1    g494(.A(new_n385_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n663_), .A2(new_n433_), .A3(new_n696_), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n653_), .A2(new_n657_), .A3(new_n696_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n697_), .B1(new_n698_), .B2(new_n433_), .ZN(G1331gat));
  NOR3_X1   g498(.A1(new_n586_), .A2(new_n546_), .A3(new_n637_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT109), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n475_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n422_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n700_), .A2(new_n701_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n702_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT110), .Z(new_n707_));
  INV_X1    g506(.A(G57gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n707_), .A2(new_n708_), .A3(new_n409_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n704_), .A2(new_n547_), .A3(new_n607_), .A4(new_n602_), .ZN(new_n710_));
  OAI21_X1  g509(.A(G57gat), .B1(new_n710_), .B2(new_n296_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT111), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n712_), .B(new_n713_), .ZN(G1332gat));
  INV_X1    g513(.A(G64gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n707_), .A2(new_n715_), .A3(new_n391_), .ZN(new_n716_));
  OAI21_X1  g515(.A(G64gat), .B1(new_n710_), .B2(new_n613_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT48), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(G1333gat));
  INV_X1    g518(.A(G71gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n707_), .A2(new_n720_), .A3(new_n684_), .ZN(new_n721_));
  OAI21_X1  g520(.A(G71gat), .B1(new_n710_), .B2(new_n421_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT49), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(G1334gat));
  INV_X1    g523(.A(G78gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n707_), .A2(new_n725_), .A3(new_n696_), .ZN(new_n726_));
  OAI21_X1  g525(.A(G78gat), .B1(new_n710_), .B2(new_n385_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT50), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1335gat));
  NAND4_X1  g528(.A1(new_n704_), .A2(new_n547_), .A3(new_n585_), .A4(new_n637_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(G85gat), .B1(new_n731_), .B2(new_n409_), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n656_), .A2(KEYINPUT112), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n656_), .A2(KEYINPUT112), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n546_), .A2(new_n703_), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n733_), .A2(new_n637_), .A3(new_n734_), .A4(new_n735_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n736_), .A2(new_n296_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n732_), .B1(new_n737_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g537(.A(G92gat), .B1(new_n731_), .B2(new_n391_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n736_), .A2(new_n613_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n740_), .B2(G92gat), .ZN(G1337gat));
  OAI21_X1  g540(.A(G99gat), .B1(new_n736_), .B2(new_n421_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n731_), .A2(new_n513_), .A3(new_n681_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT51), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT51), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n742_), .A2(new_n746_), .A3(new_n743_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(G1338gat));
  NAND4_X1  g547(.A1(new_n656_), .A2(new_n696_), .A3(new_n637_), .A4(new_n735_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(G106gat), .ZN(new_n750_));
  XOR2_X1   g549(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n751_));
  XNOR2_X1  g550(.A(new_n750_), .B(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n731_), .A2(new_n514_), .A3(new_n696_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT53), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT53), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n752_), .A2(new_n756_), .A3(new_n753_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1339gat));
  INV_X1    g557(.A(G113gat), .ZN(new_n759_));
  INV_X1    g558(.A(new_n461_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n761_));
  AOI211_X1 g560(.A(new_n761_), .B(new_n428_), .C1(new_n459_), .C2(new_n760_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n539_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT117), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT117), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n763_), .A2(new_n766_), .A3(new_n539_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n522_), .B(new_n523_), .C1(new_n529_), .C2(new_n531_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n525_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT55), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n532_), .A2(new_n771_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n528_), .B(KEYINPUT67), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n773_), .A2(KEYINPUT55), .A3(new_n526_), .A4(new_n522_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n770_), .A2(new_n772_), .A3(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n538_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n775_), .A2(KEYINPUT56), .A3(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT56), .B1(new_n775_), .B2(new_n776_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n768_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT58), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n768_), .B(KEYINPUT58), .C1(new_n777_), .C2(new_n778_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(new_n586_), .A3(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT57), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n540_), .A2(new_n475_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n786_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n785_), .B1(new_n777_), .B2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n763_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n784_), .B1(new_n790_), .B2(new_n607_), .ZN(new_n791_));
  AOI211_X1 g590(.A(KEYINPUT57), .B(new_n585_), .C1(new_n788_), .C2(new_n789_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n783_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n601_), .ZN(new_n796_));
  OAI211_X1 g595(.A(KEYINPUT118), .B(new_n783_), .C1(new_n791_), .C2(new_n792_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n795_), .A2(new_n796_), .A3(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(KEYINPUT115), .A2(KEYINPUT54), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n546_), .A2(new_n475_), .A3(new_n602_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT114), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT114), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n546_), .A2(new_n802_), .A3(new_n475_), .A4(new_n602_), .ZN(new_n803_));
  AOI211_X1 g602(.A(new_n799_), .B(new_n586_), .C1(new_n801_), .C2(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n801_), .A2(new_n803_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(new_n587_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n804_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n696_), .B1(new_n798_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n613_), .A2(new_n409_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n810_), .A2(new_n680_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n759_), .B1(new_n812_), .B2(new_n475_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT119), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(KEYINPUT59), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT120), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n793_), .A2(new_n816_), .A3(new_n637_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n808_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n816_), .B1(new_n793_), .B2(new_n637_), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT59), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n820_), .A2(new_n821_), .A3(new_n385_), .A4(new_n811_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n815_), .A2(new_n822_), .A3(G113gat), .A4(new_n703_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n824_), .B(new_n759_), .C1(new_n812_), .C2(new_n475_), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n814_), .A2(new_n823_), .A3(new_n825_), .ZN(G1340gat));
  NAND2_X1  g625(.A1(new_n815_), .A2(new_n822_), .ZN(new_n827_));
  OAI21_X1  g626(.A(G120gat), .B1(new_n827_), .B2(new_n546_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n812_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n255_), .B1(new_n546_), .B2(KEYINPUT60), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n829_), .B(new_n830_), .C1(KEYINPUT60), .C2(new_n255_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n828_), .A2(new_n831_), .ZN(G1341gat));
  NAND4_X1  g631(.A1(new_n815_), .A2(new_n822_), .A3(G127gat), .A4(new_n601_), .ZN(new_n833_));
  INV_X1    g632(.A(G127gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n812_), .B2(new_n637_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n833_), .A2(new_n835_), .ZN(G1342gat));
  AOI21_X1  g635(.A(G134gat), .B1(new_n829_), .B2(new_n585_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n827_), .ZN(new_n838_));
  XOR2_X1   g637(.A(KEYINPUT121), .B(G134gat), .Z(new_n839_));
  NAND2_X1  g638(.A1(new_n586_), .A2(new_n839_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(KEYINPUT122), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n837_), .B1(new_n838_), .B2(new_n841_), .ZN(G1343gat));
  AOI21_X1  g641(.A(new_n684_), .B1(new_n798_), .B2(new_n808_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n810_), .A2(new_n385_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n845_), .A2(new_n475_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(new_n426_), .ZN(G1344gat));
  INV_X1    g646(.A(new_n845_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n547_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g649(.A1(new_n845_), .A2(new_n637_), .ZN(new_n851_));
  XOR2_X1   g650(.A(KEYINPUT61), .B(G155gat), .Z(new_n852_));
  XNOR2_X1  g651(.A(new_n851_), .B(new_n852_), .ZN(G1346gat));
  AOI21_X1  g652(.A(G162gat), .B1(new_n848_), .B2(new_n585_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n645_), .A2(G162gat), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n848_), .B2(new_n855_), .ZN(G1347gat));
  NAND3_X1  g655(.A1(new_n684_), .A2(new_n296_), .A3(new_n391_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n475_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n385_), .B(new_n858_), .C1(new_n818_), .C2(new_n819_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(G169gat), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT62), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT124), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT123), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT62), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n859_), .A2(new_n864_), .A3(new_n865_), .A4(G169gat), .ZN(new_n866_));
  OAI21_X1  g665(.A(KEYINPUT123), .B1(new_n860_), .B2(KEYINPUT62), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n860_), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n863_), .A2(new_n866_), .A3(new_n867_), .A4(new_n868_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n820_), .A2(new_n222_), .A3(new_n385_), .A4(new_n858_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1348gat));
  INV_X1    g670(.A(new_n857_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n809_), .A2(new_n872_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n873_), .A2(new_n223_), .A3(new_n546_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n820_), .A2(new_n385_), .A3(new_n872_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n223_), .B1(new_n875_), .B2(new_n546_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT125), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  OAI211_X1 g677(.A(KEYINPUT125), .B(new_n223_), .C1(new_n875_), .C2(new_n546_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n874_), .B1(new_n878_), .B2(new_n879_), .ZN(G1349gat));
  INV_X1    g679(.A(new_n875_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n203_), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n881_), .A2(KEYINPUT126), .A3(new_n601_), .A4(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(G183gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(new_n873_), .B2(new_n637_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT126), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n820_), .A2(new_n882_), .A3(new_n385_), .A4(new_n872_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(new_n796_), .ZN(new_n888_));
  AND3_X1   g687(.A1(new_n883_), .A2(new_n885_), .A3(new_n888_), .ZN(G1350gat));
  OAI21_X1  g688(.A(G190gat), .B1(new_n875_), .B2(new_n587_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n585_), .A2(new_n204_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n875_), .B2(new_n891_), .ZN(G1351gat));
  NOR2_X1   g691(.A1(new_n613_), .A2(new_n392_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n843_), .A2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n703_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g696(.A1(new_n894_), .A2(new_n546_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(new_n310_), .ZN(G1353gat));
  NAND3_X1  g698(.A1(new_n843_), .A2(new_n601_), .A3(new_n893_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n901_));
  AND2_X1   g700(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n900_), .A2(new_n901_), .A3(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(new_n900_), .B2(new_n901_), .ZN(G1354gat));
  AOI21_X1  g703(.A(G218gat), .B1(new_n895_), .B2(new_n585_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n586_), .A2(G218gat), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(KEYINPUT127), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n905_), .B1(new_n895_), .B2(new_n907_), .ZN(G1355gat));
endmodule


