//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 0 1 0 0 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n618_,
    new_n619_, new_n620_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n803_, new_n804_, new_n805_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n838_, new_n839_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT64), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(G71gat), .B(G78gat), .Z(new_n205_));
  INV_X1    g004(.A(G57gat), .ZN(new_n206_));
  INV_X1    g005(.A(G64gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT68), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G57gat), .A2(G64gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n209_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n213_));
  NOR3_X1   g012(.A1(new_n212_), .A2(KEYINPUT11), .A3(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT11), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G57gat), .B(G64gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT68), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n215_), .B1(new_n217_), .B2(new_n211_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n205_), .B1(new_n214_), .B2(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT11), .B1(new_n212_), .B2(new_n213_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n205_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n219_), .A2(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(G85gat), .B(G92gat), .Z(new_n224_));
  INV_X1    g023(.A(KEYINPUT66), .ZN(new_n225_));
  OAI22_X1  g024(.A1(new_n225_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(KEYINPUT7), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n225_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G99gat), .A2(G106gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT6), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n229_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n224_), .B1(new_n228_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT8), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(KEYINPUT67), .A3(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(KEYINPUT10), .B(G99gat), .Z(new_n238_));
  INV_X1    g037(.A(G106gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n224_), .A2(KEYINPUT9), .ZN(new_n241_));
  NAND2_X1  g040(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n242_), .A2(KEYINPUT9), .ZN(new_n243_));
  NOR2_X1   g042(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n244_));
  OAI21_X1  g043(.A(G85gat), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  AND3_X1   g044(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n246_));
  AOI21_X1  g045(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n240_), .A2(new_n241_), .A3(new_n245_), .A4(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n226_), .A2(new_n227_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n250_), .A2(new_n248_), .A3(new_n229_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n236_), .A2(KEYINPUT67), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT8), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n251_), .A2(new_n224_), .A3(new_n252_), .A4(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n237_), .A2(new_n249_), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n223_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n223_), .A2(new_n256_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n204_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n260_), .A2(KEYINPUT69), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(KEYINPUT69), .ZN(new_n262_));
  AOI211_X1 g061(.A(new_n253_), .B(KEYINPUT8), .C1(new_n251_), .C2(new_n224_), .ZN(new_n263_));
  AND4_X1   g062(.A1(new_n224_), .A2(new_n251_), .A3(new_n252_), .A4(new_n254_), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT70), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n237_), .A2(new_n266_), .A3(new_n255_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n265_), .A2(new_n249_), .A3(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n217_), .A2(new_n215_), .A3(new_n211_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n221_), .B1(new_n220_), .B2(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n218_), .A2(new_n205_), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT71), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n219_), .A2(new_n273_), .A3(new_n222_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n268_), .A2(KEYINPUT12), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT12), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n257_), .B1(new_n259_), .B2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n276_), .A2(new_n278_), .A3(new_n203_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n261_), .A2(new_n262_), .A3(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT5), .B(G176gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(G204gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G120gat), .B(G148gat), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n282_), .B(new_n283_), .Z(new_n284_));
  NAND2_X1  g083(.A1(new_n280_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n284_), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n261_), .A2(new_n262_), .A3(new_n279_), .A4(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT13), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(G43gat), .B(G50gat), .Z(new_n291_));
  XNOR2_X1  g090(.A(G29gat), .B(G36gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT79), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G1gat), .B(G8gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT77), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT76), .B(G1gat), .ZN(new_n297_));
  INV_X1    g096(.A(G8gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT14), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G15gat), .B(G22gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n296_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n296_), .A2(new_n301_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n294_), .B(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n304_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(new_n294_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n293_), .B(KEYINPUT15), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n307_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G229gat), .A2(G233gat), .ZN(new_n310_));
  MUX2_X1   g109(.A(new_n305_), .B(new_n309_), .S(new_n310_), .Z(new_n311_));
  XOR2_X1   g110(.A(KEYINPUT81), .B(G113gat), .Z(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT82), .B(G141gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G169gat), .B(G197gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT80), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n311_), .B(new_n318_), .Z(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n290_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G127gat), .B(G134gat), .ZN(new_n323_));
  INV_X1    g122(.A(G120gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT91), .B(G113gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G15gat), .B(G43gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT31), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n327_), .B(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(G169gat), .ZN(new_n332_));
  INV_X1    g131(.A(G176gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G169gat), .A2(G176gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(KEYINPUT24), .A3(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT83), .B(G183gat), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n337_), .B1(new_n338_), .B2(KEYINPUT25), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT26), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(G190gat), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT84), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(G190gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT26), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n340_), .A2(KEYINPUT84), .A3(G190gat), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n343_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n336_), .B1(new_n339_), .B2(new_n347_), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n348_), .A2(KEYINPUT85), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT23), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n350_), .A2(G183gat), .A3(G190gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT86), .ZN(new_n352_));
  INV_X1    g151(.A(G183gat), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT23), .B1(new_n353_), .B2(new_n344_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n334_), .A2(KEYINPUT24), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n348_), .A2(KEYINPUT85), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n349_), .A2(new_n355_), .A3(new_n356_), .A4(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n354_), .A2(new_n351_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n359_), .B1(G190gat), .B2(new_n338_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n332_), .A2(KEYINPUT88), .ZN(new_n361_));
  AND2_X1   g160(.A1(KEYINPUT87), .A2(KEYINPUT22), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(KEYINPUT87), .B1(new_n332_), .B2(KEYINPUT22), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n364_), .A2(G176gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n366_), .A2(KEYINPUT89), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(KEYINPUT89), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n360_), .B(new_n335_), .C1(new_n367_), .C2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n358_), .A2(new_n369_), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n370_), .A2(G227gat), .A3(G233gat), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n370_), .B1(G227gat), .B2(G233gat), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT90), .B(KEYINPUT30), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT92), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n375_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n377_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G71gat), .B(G99gat), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n376_), .A2(new_n378_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n380_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n331_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n383_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(new_n330_), .A3(new_n381_), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n384_), .A2(new_n386_), .A3(KEYINPUT93), .ZN(new_n387_));
  AOI21_X1  g186(.A(KEYINPUT93), .B1(new_n384_), .B2(new_n386_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(G141gat), .A2(G148gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G141gat), .A2(G148gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT94), .B(KEYINPUT95), .ZN(new_n393_));
  NOR2_X1   g192(.A1(G155gat), .A2(G162gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G155gat), .A2(G162gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT1), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n391_), .B(new_n392_), .C1(new_n395_), .C2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n394_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n393_), .B(new_n399_), .ZN(new_n400_));
  XOR2_X1   g199(.A(new_n392_), .B(KEYINPUT2), .Z(new_n401_));
  XOR2_X1   g200(.A(new_n390_), .B(KEYINPUT3), .Z(new_n402_));
  OAI211_X1 g201(.A(new_n400_), .B(new_n396_), .C1(new_n401_), .C2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n398_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT96), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT96), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n398_), .A2(new_n403_), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT29), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(G22gat), .B(G50gat), .Z(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(KEYINPUT28), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n411_), .B(new_n413_), .ZN(new_n414_));
  XOR2_X1   g213(.A(G211gat), .B(G218gat), .Z(new_n415_));
  INV_X1    g214(.A(G197gat), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n416_), .A2(G204gat), .ZN(new_n417_));
  XOR2_X1   g216(.A(KEYINPUT97), .B(G197gat), .Z(new_n418_));
  AOI21_X1  g217(.A(new_n417_), .B1(new_n418_), .B2(G204gat), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT21), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n415_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G197gat), .A2(G204gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT97), .B(G197gat), .ZN(new_n423_));
  OAI211_X1 g222(.A(KEYINPUT21), .B(new_n422_), .C1(new_n423_), .C2(G204gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G211gat), .B(G218gat), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n419_), .A2(new_n425_), .ZN(new_n426_));
  AOI22_X1  g225(.A1(new_n421_), .A2(new_n424_), .B1(new_n426_), .B2(KEYINPUT21), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G228gat), .A2(G233gat), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n428_), .B(new_n429_), .C1(new_n409_), .C2(new_n410_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n410_), .B1(new_n398_), .B2(new_n403_), .ZN(new_n431_));
  OAI211_X1 g230(.A(G228gat), .B(G233gat), .C1(new_n431_), .C2(new_n427_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G78gat), .B(G106gat), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n430_), .A2(new_n432_), .A3(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n434_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n436_));
  OR3_X1    g235(.A1(new_n414_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n414_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G1gat), .B(G29gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(G85gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(KEYINPUT0), .B(G57gat), .ZN(new_n442_));
  XOR2_X1   g241(.A(new_n441_), .B(new_n442_), .Z(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n327_), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n398_), .A2(new_n403_), .A3(new_n406_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n406_), .B1(new_n398_), .B2(new_n403_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n445_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G225gat), .A2(G233gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT101), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n327_), .A2(new_n398_), .A3(new_n403_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n448_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT4), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n453_), .B1(new_n448_), .B2(new_n451_), .ZN(new_n454_));
  AOI21_X1  g253(.A(KEYINPUT4), .B1(new_n408_), .B2(new_n445_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n444_), .B(new_n452_), .C1(new_n456_), .C2(new_n450_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT25), .B(G183gat), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(new_n345_), .A3(new_n341_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n459_), .A2(new_n359_), .A3(new_n356_), .A4(new_n336_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n353_), .A2(new_n344_), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n355_), .A2(new_n461_), .B1(G169gat), .B2(G176gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT22), .B(G169gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n333_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n462_), .A2(KEYINPUT98), .A3(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT98), .B1(new_n462_), .B2(new_n464_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n460_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(new_n428_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n358_), .A2(new_n369_), .A3(new_n427_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n468_), .A2(KEYINPUT20), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G226gat), .A2(G233gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT19), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT20), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n474_), .B1(new_n370_), .B2(new_n428_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n472_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n475_), .B(new_n476_), .C1(new_n428_), .C2(new_n467_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n473_), .A2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G8gat), .B(G36gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT100), .ZN(new_n480_));
  XOR2_X1   g279(.A(G64gat), .B(G92gat), .Z(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n478_), .A2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n484_), .B1(new_n473_), .B2(new_n477_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n450_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n448_), .A2(new_n451_), .ZN(new_n490_));
  OR2_X1    g289(.A1(new_n490_), .A2(new_n450_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n489_), .A2(KEYINPUT102), .A3(new_n491_), .ZN(new_n492_));
  OR3_X1    g291(.A1(new_n490_), .A2(KEYINPUT102), .A3(new_n450_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n444_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT33), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  AOI211_X1 g295(.A(KEYINPUT33), .B(new_n444_), .C1(new_n492_), .C2(new_n493_), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n457_), .B(new_n488_), .C1(new_n496_), .C2(new_n497_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n468_), .A2(KEYINPUT20), .A3(new_n476_), .A4(new_n469_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n462_), .A2(new_n464_), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n500_), .A2(new_n427_), .A3(new_n460_), .ZN(new_n501_));
  AOI211_X1 g300(.A(new_n474_), .B(new_n501_), .C1(new_n370_), .C2(new_n428_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n499_), .B1(new_n502_), .B2(new_n476_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT103), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n484_), .A2(KEYINPUT32), .ZN(new_n505_));
  AND3_X1   g304(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n504_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n478_), .A2(new_n505_), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n492_), .A2(new_n444_), .A3(new_n493_), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n508_), .B(new_n509_), .C1(new_n510_), .C2(new_n494_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n439_), .B1(new_n498_), .B2(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n510_), .A2(new_n494_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n439_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT27), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n515_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n485_), .A2(KEYINPUT104), .ZN(new_n517_));
  OR2_X1    g316(.A1(new_n485_), .A2(KEYINPUT104), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n503_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n519_), .B(KEYINPUT27), .C1(new_n485_), .C2(new_n478_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n516_), .A2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n514_), .A2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n389_), .B1(new_n512_), .B2(new_n522_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n384_), .A2(new_n386_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n521_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n439_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n524_), .A2(new_n525_), .A3(new_n513_), .A4(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n322_), .B1(new_n523_), .B2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G232gat), .A2(G233gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT35), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n256_), .A2(new_n293_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT75), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n308_), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n268_), .A2(KEYINPUT73), .A3(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(KEYINPUT73), .B1(new_n268_), .B2(new_n537_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n533_), .B(new_n536_), .C1(new_n538_), .C2(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n531_), .A2(new_n532_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n268_), .A2(new_n537_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT73), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n268_), .A2(KEYINPUT73), .A3(new_n537_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n541_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n547_), .A2(new_n548_), .A3(new_n533_), .A4(new_n536_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n542_), .A2(new_n549_), .A3(KEYINPUT74), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G190gat), .B(G218gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G134gat), .B(G162gat), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n551_), .B(new_n552_), .Z(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n554_), .A2(KEYINPUT36), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n550_), .A2(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n535_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n548_), .B1(new_n557_), .B2(new_n533_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n540_), .A2(new_n541_), .ZN(new_n559_));
  OAI211_X1 g358(.A(KEYINPUT36), .B(new_n554_), .C1(new_n558_), .C2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n555_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n542_), .A2(new_n549_), .A3(KEYINPUT74), .A4(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n556_), .A2(new_n560_), .A3(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT37), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n275_), .B(KEYINPUT78), .Z(new_n565_));
  NAND2_X1  g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n304_), .B(new_n566_), .Z(new_n567_));
  XNOR2_X1  g366(.A(new_n565_), .B(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(G127gat), .B(G155gat), .Z(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(G211gat), .ZN(new_n570_));
  XOR2_X1   g369(.A(KEYINPUT16), .B(G183gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n568_), .A2(KEYINPUT17), .A3(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n567_), .B(new_n223_), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n572_), .B(KEYINPUT17), .Z(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT37), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n556_), .A2(new_n560_), .A3(new_n578_), .A4(new_n562_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n564_), .A2(new_n577_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n528_), .A2(new_n580_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n581_), .A2(KEYINPUT105), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(KEYINPUT105), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n513_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n297_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT107), .ZN(new_n588_));
  OR3_X1    g387(.A1(new_n587_), .A2(new_n588_), .A3(KEYINPUT38), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n563_), .B(KEYINPUT106), .Z(new_n590_));
  INV_X1    g389(.A(new_n577_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n528_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(new_n585_), .ZN(new_n595_));
  AOI22_X1  g394(.A1(new_n587_), .A2(KEYINPUT38), .B1(G1gat), .B2(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n588_), .B1(new_n587_), .B2(KEYINPUT38), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n589_), .A2(new_n596_), .A3(new_n597_), .ZN(G1324gat));
  XNOR2_X1  g397(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n594_), .A2(new_n521_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(G8gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT39), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n298_), .B(new_n521_), .C1(new_n582_), .C2(new_n583_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n599_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n601_), .A2(KEYINPUT39), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT39), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n606_), .B1(new_n600_), .B2(G8gat), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n603_), .B(new_n599_), .C1(new_n605_), .C2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n604_), .A2(new_n609_), .ZN(G1325gat));
  OAI21_X1  g409(.A(G15gat), .B1(new_n593_), .B2(new_n389_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT109), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT41), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n613_), .ZN(new_n615_));
  OR3_X1    g414(.A1(new_n581_), .A2(G15gat), .A3(new_n389_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n614_), .A2(new_n615_), .A3(new_n616_), .ZN(G1326gat));
  OAI21_X1  g416(.A(G22gat), .B1(new_n593_), .B2(new_n526_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT42), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n526_), .A2(G22gat), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n619_), .B1(new_n581_), .B2(new_n620_), .ZN(G1327gat));
  INV_X1    g420(.A(new_n563_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n622_), .A2(new_n577_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n528_), .A2(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(G29gat), .B1(new_n624_), .B2(new_n585_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n523_), .A2(new_n527_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n564_), .A2(new_n579_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT111), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n626_), .A2(new_n631_), .A3(KEYINPUT43), .A4(new_n627_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n321_), .A2(new_n591_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT110), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n630_), .A2(new_n632_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT44), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n629_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n638_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n627_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n631_), .A2(KEYINPUT43), .ZN(new_n641_));
  AOI211_X1 g440(.A(new_n640_), .B(new_n641_), .C1(new_n523_), .C2(new_n527_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n639_), .A2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n643_), .A2(KEYINPUT44), .A3(new_n634_), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n637_), .A2(new_n585_), .A3(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n625_), .B1(new_n645_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g445(.A(G36gat), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n521_), .B(KEYINPUT112), .Z(new_n648_));
  NAND4_X1  g447(.A1(new_n528_), .A2(new_n647_), .A3(new_n623_), .A4(new_n648_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT45), .Z(new_n650_));
  NAND3_X1  g449(.A1(new_n637_), .A2(new_n644_), .A3(new_n521_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n651_), .B2(G36gat), .ZN(new_n652_));
  NOR2_X1   g451(.A1(KEYINPUT113), .A2(KEYINPUT46), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n653_), .ZN(new_n655_));
  AOI211_X1 g454(.A(new_n655_), .B(new_n650_), .C1(new_n651_), .C2(G36gat), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n654_), .A2(new_n656_), .ZN(G1329gat));
  NAND4_X1  g456(.A1(new_n637_), .A2(new_n644_), .A3(G43gat), .A4(new_n524_), .ZN(new_n658_));
  INV_X1    g457(.A(G43gat), .ZN(new_n659_));
  INV_X1    g458(.A(new_n624_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n659_), .B1(new_n660_), .B2(new_n389_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n658_), .A2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(KEYINPUT114), .B(KEYINPUT47), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(G1330gat));
  AOI21_X1  g463(.A(G50gat), .B1(new_n624_), .B2(new_n439_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n637_), .A2(new_n439_), .A3(new_n644_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n666_), .B2(G50gat), .ZN(G1331gat));
  NOR2_X1   g466(.A1(new_n289_), .A2(new_n319_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n626_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(new_n592_), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n670_), .A2(new_n206_), .A3(new_n513_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n669_), .A2(new_n580_), .A3(new_n585_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n206_), .B2(new_n672_), .ZN(G1332gat));
  INV_X1    g472(.A(new_n648_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G64gat), .B1(new_n670_), .B2(new_n674_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT48), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n669_), .A2(new_n580_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n648_), .A2(new_n207_), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT115), .Z(new_n679_));
  OAI21_X1  g478(.A(new_n676_), .B1(new_n677_), .B2(new_n679_), .ZN(G1333gat));
  OAI21_X1  g479(.A(G71gat), .B1(new_n670_), .B2(new_n389_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT49), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n389_), .A2(G71gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n682_), .B1(new_n677_), .B2(new_n683_), .ZN(G1334gat));
  OAI21_X1  g483(.A(G78gat), .B1(new_n670_), .B2(new_n526_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT50), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n526_), .A2(G78gat), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n686_), .B1(new_n677_), .B2(new_n687_), .ZN(G1335gat));
  AND2_X1   g487(.A1(new_n669_), .A2(new_n623_), .ZN(new_n689_));
  AOI21_X1  g488(.A(G85gat), .B1(new_n689_), .B2(new_n585_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n630_), .A2(new_n591_), .A3(new_n632_), .A4(new_n668_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n691_), .A2(new_n513_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n690_), .B1(new_n692_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g492(.A(G92gat), .B1(new_n689_), .B2(new_n521_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n691_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n244_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n674_), .B1(new_n696_), .B2(new_n242_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n694_), .B1(new_n695_), .B2(new_n697_), .ZN(G1337gat));
  OAI21_X1  g497(.A(G99gat), .B1(new_n691_), .B2(new_n389_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n689_), .A2(new_n238_), .A3(new_n524_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g501(.A1(new_n689_), .A2(new_n239_), .A3(new_n439_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT52), .ZN(new_n704_));
  OAI211_X1 g503(.A(new_n704_), .B(G106gat), .C1(new_n691_), .C2(new_n526_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n643_), .A2(new_n591_), .A3(new_n439_), .A4(new_n668_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n704_), .B1(new_n707_), .B2(G106gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n703_), .B1(new_n706_), .B2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT53), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT53), .ZN(new_n711_));
  OAI211_X1 g510(.A(new_n711_), .B(new_n703_), .C1(new_n706_), .C2(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(G1339gat));
  INV_X1    g512(.A(KEYINPUT117), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n203_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT55), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n279_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n276_), .A2(new_n278_), .A3(KEYINPUT55), .A4(new_n203_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n284_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT56), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT56), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n719_), .A2(new_n722_), .A3(new_n284_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n721_), .A2(new_n319_), .A3(new_n287_), .A4(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n309_), .A2(G229gat), .A3(G233gat), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n305_), .A2(new_n310_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n316_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n727_), .B1(new_n316_), .B2(new_n311_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n288_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n724_), .A2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(new_n622_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT57), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n563_), .B1(new_n724_), .B2(new_n729_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT57), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n721_), .A2(new_n287_), .A3(new_n728_), .A4(new_n723_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT58), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n722_), .B1(new_n719_), .B2(new_n284_), .ZN(new_n739_));
  AOI211_X1 g538(.A(KEYINPUT56), .B(new_n286_), .C1(new_n717_), .C2(new_n718_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n741_), .A2(KEYINPUT58), .A3(new_n287_), .A4(new_n728_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n627_), .A2(new_n738_), .A3(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n733_), .A2(new_n735_), .A3(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n591_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT54), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n580_), .A2(new_n746_), .A3(new_n320_), .A4(new_n289_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n564_), .A2(new_n289_), .A3(new_n577_), .A4(new_n579_), .ZN(new_n748_));
  OAI21_X1  g547(.A(KEYINPUT54), .B1(new_n748_), .B2(new_n319_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n745_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT59), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n524_), .A2(new_n525_), .A3(new_n585_), .A4(new_n526_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n751_), .A2(new_n752_), .A3(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT116), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n745_), .A2(new_n756_), .A3(new_n750_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n745_), .B2(new_n750_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n757_), .A2(new_n758_), .A3(new_n753_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n319_), .B(new_n755_), .C1(new_n759_), .C2(new_n752_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(G113gat), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n734_), .B(new_n732_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n577_), .B1(new_n762_), .B2(new_n743_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n747_), .A2(new_n749_), .ZN(new_n764_));
  OAI21_X1  g563(.A(KEYINPUT116), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n745_), .A2(new_n756_), .A3(new_n750_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n765_), .A2(new_n319_), .A3(new_n766_), .A4(new_n754_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n767_), .A2(G113gat), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n714_), .B1(new_n761_), .B2(new_n769_), .ZN(new_n770_));
  AOI211_X1 g569(.A(KEYINPUT117), .B(new_n768_), .C1(new_n760_), .C2(G113gat), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(G1340gat));
  OAI21_X1  g571(.A(new_n324_), .B1(new_n289_), .B2(KEYINPUT60), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n759_), .B(new_n773_), .C1(KEYINPUT60), .C2(new_n324_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n755_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n759_), .ZN(new_n776_));
  AOI211_X1 g575(.A(new_n289_), .B(new_n775_), .C1(new_n776_), .C2(KEYINPUT59), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n774_), .B1(new_n777_), .B2(new_n324_), .ZN(G1341gat));
  AOI21_X1  g577(.A(G127gat), .B1(new_n759_), .B2(new_n577_), .ZN(new_n779_));
  INV_X1    g578(.A(G127gat), .ZN(new_n780_));
  AOI211_X1 g579(.A(new_n780_), .B(new_n775_), .C1(new_n776_), .C2(KEYINPUT59), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n779_), .B1(new_n781_), .B2(new_n577_), .ZN(G1342gat));
  AOI21_X1  g581(.A(G134gat), .B1(new_n759_), .B2(new_n590_), .ZN(new_n783_));
  AOI211_X1 g582(.A(new_n640_), .B(new_n775_), .C1(new_n776_), .C2(KEYINPUT59), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(G134gat), .ZN(G1343gat));
  NOR2_X1   g584(.A1(new_n757_), .A2(new_n758_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n389_), .ZN(new_n787_));
  NOR4_X1   g586(.A1(new_n648_), .A2(new_n787_), .A3(new_n513_), .A4(new_n526_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT118), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n786_), .A2(new_n789_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n790_), .A2(new_n320_), .ZN(new_n791_));
  XOR2_X1   g590(.A(KEYINPUT119), .B(G141gat), .Z(new_n792_));
  XNOR2_X1  g591(.A(new_n791_), .B(new_n792_), .ZN(G1344gat));
  NOR2_X1   g592(.A1(new_n790_), .A2(new_n289_), .ZN(new_n794_));
  XOR2_X1   g593(.A(new_n794_), .B(G148gat), .Z(G1345gat));
  OAI21_X1  g594(.A(KEYINPUT120), .B1(new_n790_), .B2(new_n591_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT120), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n786_), .A2(new_n789_), .A3(new_n797_), .A4(new_n577_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(KEYINPUT61), .B(G155gat), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n796_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n800_), .A2(new_n801_), .ZN(G1346gat));
  INV_X1    g601(.A(G162gat), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n790_), .A2(new_n803_), .A3(new_n640_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n786_), .A2(new_n789_), .A3(new_n590_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n804_), .B1(new_n803_), .B2(new_n805_), .ZN(G1347gat));
  NOR3_X1   g605(.A1(new_n674_), .A2(new_n585_), .A3(new_n389_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n751_), .A2(new_n526_), .A3(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n808_), .A2(KEYINPUT121), .A3(new_n319_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n751_), .A2(new_n319_), .A3(new_n526_), .A4(new_n807_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT121), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n809_), .A2(G169gat), .A3(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT122), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n809_), .A2(KEYINPUT122), .A3(G169gat), .A4(new_n812_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(KEYINPUT62), .A3(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n808_), .A2(new_n319_), .A3(new_n463_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT62), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n813_), .A2(new_n814_), .A3(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n817_), .A2(new_n818_), .A3(new_n820_), .ZN(G1348gat));
  AOI21_X1  g620(.A(G176gat), .B1(new_n808_), .B2(new_n290_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n765_), .A2(new_n526_), .A3(new_n766_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT123), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT123), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n765_), .A2(new_n825_), .A3(new_n526_), .A4(new_n766_), .ZN(new_n826_));
  AOI211_X1 g625(.A(new_n333_), .B(new_n289_), .C1(new_n824_), .C2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n822_), .B1(new_n827_), .B2(new_n807_), .ZN(G1349gat));
  INV_X1    g627(.A(new_n458_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n808_), .A2(new_n577_), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n807_), .A2(new_n577_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n831_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n830_), .B1(new_n832_), .B2(new_n338_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT124), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT124), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n835_), .B(new_n830_), .C1(new_n832_), .C2(new_n338_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(G1350gat));
  NAND4_X1  g636(.A1(new_n808_), .A2(new_n345_), .A3(new_n341_), .A4(new_n590_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n808_), .A2(new_n627_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n839_), .B2(new_n344_), .ZN(G1351gat));
  NOR4_X1   g639(.A1(new_n757_), .A2(new_n758_), .A3(new_n787_), .A4(new_n674_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n514_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n843_), .A2(new_n320_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(new_n416_), .ZN(G1352gat));
  INV_X1    g644(.A(new_n843_), .ZN(new_n846_));
  AOI21_X1  g645(.A(G204gat), .B1(new_n846_), .B2(new_n290_), .ZN(new_n847_));
  INV_X1    g646(.A(G204gat), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n843_), .A2(new_n848_), .A3(new_n289_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n847_), .A2(new_n849_), .ZN(G1353gat));
  NOR2_X1   g649(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(KEYINPUT125), .ZN(new_n852_));
  NAND2_X1  g651(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n846_), .A2(new_n577_), .A3(new_n852_), .A4(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n852_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n841_), .A2(new_n577_), .A3(new_n842_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n853_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n855_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n854_), .A2(new_n858_), .ZN(G1354gat));
  NOR3_X1   g658(.A1(new_n757_), .A2(new_n758_), .A3(new_n787_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n860_), .A2(new_n842_), .A3(new_n590_), .A4(new_n648_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT126), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n841_), .A2(KEYINPUT126), .A3(new_n842_), .A4(new_n590_), .ZN(new_n864_));
  INV_X1    g663(.A(G218gat), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n863_), .A2(new_n864_), .A3(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n846_), .A2(G218gat), .A3(new_n627_), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1355gat));
endmodule


