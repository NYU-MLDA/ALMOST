//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 0 0 0 1 1 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 0 0 1 0 1 0 0 1 0 0 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n629_, new_n630_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n796_, new_n797_,
    new_n798_, new_n800_, new_n801_, new_n803_, new_n804_, new_n805_,
    new_n807_, new_n808_, new_n809_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n826_, new_n827_,
    new_n829_, new_n830_, new_n832_, new_n833_, new_n834_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n849_;
  XOR2_X1   g000(.A(KEYINPUT85), .B(G176gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT22), .B(G169gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205_));
  INV_X1    g004(.A(G183gat), .ZN(new_n206_));
  INV_X1    g005(.A(G190gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT23), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT84), .B(KEYINPUT23), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(new_n208_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n204_), .B(new_n205_), .C1(new_n214_), .C2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n209_), .A2(new_n211_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n217_), .B1(new_n218_), .B2(new_n209_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT25), .B(G183gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT26), .B(G190gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  OR2_X1    g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(KEYINPUT24), .A3(new_n205_), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n223_), .A2(KEYINPUT24), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n222_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n216_), .B1(new_n219_), .B2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT30), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G15gat), .B(G43gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G71gat), .B(G99gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G227gat), .A2(G233gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT86), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n231_), .B(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n228_), .B(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n235_), .B(KEYINPUT31), .Z(new_n236_));
  XNOR2_X1  g035(.A(G127gat), .B(G134gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G113gat), .B(G120gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n236_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n236_), .A2(new_n240_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G22gat), .B(G50gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT90), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(G197gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(G204gat), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n247_), .A2(G204gat), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT21), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G211gat), .B(G218gat), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n250_), .B1(KEYINPUT92), .B2(new_n248_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n253_), .B1(KEYINPUT92), .B2(new_n248_), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n251_), .B(new_n252_), .C1(new_n254_), .C2(KEYINPUT21), .ZN(new_n255_));
  INV_X1    g054(.A(new_n252_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n254_), .A2(KEYINPUT21), .A3(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G141gat), .A2(G148gat), .ZN(new_n259_));
  NOR2_X1   g058(.A1(G141gat), .A2(G148gat), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n260_), .A2(KEYINPUT87), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(KEYINPUT87), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n259_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G155gat), .A2(G162gat), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n264_), .A2(KEYINPUT1), .ZN(new_n265_));
  NOR2_X1   g064(.A1(G155gat), .A2(G162gat), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n264_), .B1(new_n266_), .B2(KEYINPUT1), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT88), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n265_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  OAI211_X1 g068(.A(KEYINPUT88), .B(new_n264_), .C1(new_n266_), .C2(KEYINPUT1), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n263_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT89), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT3), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT2), .ZN(new_n275_));
  AOI22_X1  g074(.A1(new_n260_), .A2(new_n274_), .B1(new_n259_), .B2(new_n275_), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n273_), .B(new_n276_), .C1(new_n274_), .C2(new_n260_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n264_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n278_), .A2(new_n266_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n271_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT29), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n258_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n282_), .B(KEYINPUT91), .Z(new_n283_));
  INV_X1    g082(.A(G228gat), .ZN(new_n284_));
  INV_X1    g083(.A(G233gat), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n283_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G78gat), .B(G106gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n286_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n283_), .B(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n288_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n280_), .A2(new_n281_), .ZN(new_n294_));
  XOR2_X1   g093(.A(new_n294_), .B(KEYINPUT28), .Z(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n289_), .A2(new_n293_), .A3(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n296_), .B1(new_n289_), .B2(new_n293_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n246_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n287_), .A2(new_n288_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n291_), .A2(new_n292_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n295_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n289_), .A2(new_n293_), .A3(new_n296_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n302_), .A2(new_n245_), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n299_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT98), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n203_), .B(KEYINPUT95), .Z(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n202_), .ZN(new_n309_));
  OAI221_X1 g108(.A(new_n205_), .B1(new_n215_), .B2(new_n219_), .C1(new_n308_), .C2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n213_), .A2(new_n225_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT94), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n205_), .A2(KEYINPUT24), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT93), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(new_n223_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n222_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n310_), .B1(new_n312_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n258_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n318_), .B(KEYINPUT20), .C1(new_n227_), .C2(new_n258_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G226gat), .A2(G233gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT19), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G8gat), .B(G36gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT18), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G64gat), .B(G92gat), .ZN(new_n325_));
  XOR2_X1   g124(.A(new_n324_), .B(new_n325_), .Z(new_n326_));
  AND2_X1   g125(.A1(new_n227_), .A2(new_n258_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n327_), .A2(new_n321_), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n328_), .B(KEYINPUT20), .C1(new_n258_), .C2(new_n317_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n322_), .A2(new_n326_), .A3(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT97), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n317_), .A2(new_n258_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT20), .ZN(new_n333_));
  NOR3_X1   g132(.A1(new_n332_), .A2(KEYINPUT96), .A3(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT96), .B1(new_n332_), .B2(new_n333_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n327_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n321_), .B1(new_n334_), .B2(new_n337_), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n319_), .A2(new_n321_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n326_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT27), .B1(new_n331_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n330_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n326_), .B1(new_n322_), .B2(new_n329_), .ZN(new_n343_));
  OR3_X1    g142(.A1(new_n342_), .A2(KEYINPUT27), .A3(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n341_), .A2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n280_), .B(new_n239_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT4), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  OR3_X1    g147(.A1(new_n280_), .A2(KEYINPUT4), .A3(new_n239_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G225gat), .A2(G233gat), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  OAI22_X1  g151(.A1(new_n348_), .A2(new_n352_), .B1(new_n346_), .B2(new_n351_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G1gat), .B(G29gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT0), .ZN(new_n355_));
  INV_X1    g154(.A(G57gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(G85gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n353_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n353_), .A2(new_n359_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n305_), .A2(new_n306_), .A3(new_n345_), .A4(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n360_), .B(KEYINPUT33), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n342_), .A2(new_n343_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n349_), .A2(new_n350_), .ZN(new_n367_));
  OAI221_X1 g166(.A(new_n359_), .B1(new_n346_), .B2(new_n350_), .C1(new_n348_), .C2(new_n367_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n365_), .A2(new_n366_), .A3(new_n368_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n338_), .A2(KEYINPUT32), .A3(new_n326_), .A4(new_n339_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n322_), .A2(new_n329_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n326_), .A2(KEYINPUT32), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n363_), .B1(new_n370_), .B2(new_n373_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n299_), .B(new_n304_), .C1(new_n369_), .C2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n364_), .A2(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n362_), .B1(new_n299_), .B2(new_n304_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n306_), .B1(new_n377_), .B2(new_n345_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n243_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n345_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n380_), .A2(new_n305_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n243_), .A2(new_n362_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n379_), .A2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G29gat), .B(G36gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT75), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G43gat), .B(G50gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT15), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT69), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G99gat), .A2(G106gat), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  AND2_X1   g191(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n393_));
  NOR2_X1   g192(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n392_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT65), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT6), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(new_n391_), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n395_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT7), .ZN(new_n402_));
  INV_X1    g201(.A(G99gat), .ZN(new_n403_));
  INV_X1    g202(.A(G106gat), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n402_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n401_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(G92gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n358_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT67), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G85gat), .A2(G92gat), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n411_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n409_), .A2(KEYINPUT8), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT8), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n407_), .B1(new_n395_), .B2(new_n400_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n417_), .B1(new_n418_), .B2(new_n414_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n416_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT66), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n395_), .A2(new_n400_), .ZN(new_n422_));
  OR2_X1    g221(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(new_n404_), .A3(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n411_), .A2(KEYINPUT9), .A3(new_n413_), .ZN(new_n426_));
  OR2_X1    g225(.A1(new_n413_), .A2(KEYINPUT9), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n425_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n421_), .B1(new_n422_), .B2(new_n428_), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n426_), .A2(new_n427_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n430_), .A2(new_n401_), .A3(KEYINPUT66), .A4(new_n425_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n390_), .B1(new_n420_), .B2(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT8), .B1(new_n409_), .B2(new_n415_), .ZN(new_n434_));
  AOI211_X1 g233(.A(new_n417_), .B(new_n414_), .C1(new_n401_), .C2(new_n408_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n429_), .A2(new_n431_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n437_), .A3(KEYINPUT69), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n389_), .A2(new_n433_), .A3(new_n438_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n416_), .A2(new_n419_), .A3(new_n431_), .A4(new_n429_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n388_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G232gat), .A2(G233gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT34), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n439_), .B(new_n442_), .C1(KEYINPUT35), .C2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(KEYINPUT35), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G190gat), .B(G218gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT76), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G134gat), .B(G162gat), .ZN(new_n451_));
  XOR2_X1   g250(.A(new_n450_), .B(new_n451_), .Z(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(KEYINPUT36), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n448_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n452_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n455_), .A2(KEYINPUT36), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n447_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n454_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n384_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G230gat), .A2(G233gat), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n460_), .B(KEYINPUT64), .Z(new_n461_));
  INV_X1    g260(.A(G64gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(G57gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n356_), .A2(G64gat), .ZN(new_n464_));
  AOI21_X1  g263(.A(KEYINPUT11), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G71gat), .B(G78gat), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT68), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  AND2_X1   g266(.A1(G71gat), .A2(G78gat), .ZN(new_n468_));
  NOR2_X1   g267(.A1(G71gat), .A2(G78gat), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT68), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G57gat), .B(G64gat), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n470_), .B(new_n471_), .C1(new_n472_), .C2(KEYINPUT11), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(KEYINPUT11), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n467_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n474_), .B1(new_n467_), .B2(new_n473_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n440_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n440_), .A2(new_n477_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n461_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT12), .B1(new_n440_), .B2(new_n477_), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n481_), .A2(new_n479_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT12), .ZN(new_n483_));
  NOR3_X1   g282(.A1(new_n475_), .A2(new_n476_), .A3(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n438_), .A2(new_n433_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT70), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT70), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n438_), .A2(new_n433_), .A3(new_n487_), .A4(new_n484_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n482_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n480_), .B1(new_n489_), .B2(new_n461_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G120gat), .B(G148gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G176gat), .B(G204gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(KEYINPUT71), .B(KEYINPUT5), .Z(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n490_), .A2(new_n495_), .ZN(new_n496_));
  XOR2_X1   g295(.A(new_n495_), .B(KEYINPUT72), .Z(new_n497_));
  OAI21_X1  g296(.A(new_n496_), .B1(new_n490_), .B2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n498_), .B1(KEYINPUT73), .B2(KEYINPUT13), .ZN(new_n499_));
  OR3_X1    g298(.A1(new_n499_), .A2(KEYINPUT73), .A3(KEYINPUT13), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n499_), .B1(KEYINPUT73), .B2(KEYINPUT13), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n502_), .A2(KEYINPUT74), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n502_), .A2(KEYINPUT74), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G15gat), .B(G22gat), .ZN(new_n505_));
  INV_X1    g304(.A(G1gat), .ZN(new_n506_));
  INV_X1    g305(.A(G8gat), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT14), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n505_), .A2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G1gat), .B(G8gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(new_n388_), .B(new_n511_), .Z(new_n512_));
  NAND2_X1  g311(.A1(G229gat), .A2(G233gat), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  MUX2_X1   g313(.A(new_n388_), .B(new_n389_), .S(new_n511_), .Z(new_n515_));
  AOI21_X1  g314(.A(new_n514_), .B1(new_n515_), .B2(new_n513_), .ZN(new_n516_));
  XOR2_X1   g315(.A(G169gat), .B(G197gat), .Z(new_n517_));
  XOR2_X1   g316(.A(new_n517_), .B(KEYINPUT82), .Z(new_n518_));
  XOR2_X1   g317(.A(G113gat), .B(G141gat), .Z(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT81), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n518_), .B(new_n520_), .ZN(new_n521_));
  OR2_X1    g320(.A1(new_n516_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT83), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n516_), .A2(new_n521_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n522_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n516_), .A2(KEYINPUT83), .A3(new_n521_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NOR3_X1   g326(.A1(new_n503_), .A2(new_n504_), .A3(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G127gat), .B(G155gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT16), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT78), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G183gat), .B(G211gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(KEYINPUT79), .B1(new_n533_), .B2(KEYINPUT17), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G231gat), .A2(G233gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n511_), .B(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(new_n477_), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n534_), .A2(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n533_), .A2(KEYINPUT17), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n539_), .B1(new_n534_), .B2(new_n537_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n528_), .A2(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n459_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(G1gat), .B1(new_n544_), .B2(new_n363_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n384_), .A2(new_n528_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n458_), .A2(KEYINPUT37), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT37), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n453_), .B(KEYINPUT77), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n447_), .A2(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n548_), .B1(new_n550_), .B2(new_n457_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n547_), .A2(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n541_), .B(KEYINPUT80), .Z(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n546_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT99), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT38), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n363_), .A2(G1gat), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n557_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n558_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n545_), .B1(new_n560_), .B2(new_n561_), .ZN(G1324gat));
  NAND2_X1  g361(.A1(new_n543_), .A2(new_n380_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(G8gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT39), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n557_), .A2(new_n507_), .A3(new_n380_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(G1325gat));
  INV_X1    g368(.A(G15gat), .ZN(new_n570_));
  INV_X1    g369(.A(new_n243_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n557_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n570_), .B1(new_n543_), .B2(new_n571_), .ZN(new_n573_));
  XOR2_X1   g372(.A(KEYINPUT101), .B(KEYINPUT41), .Z(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n572_), .A2(new_n575_), .ZN(G1326gat));
  INV_X1    g375(.A(G22gat), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n577_), .B1(new_n543_), .B2(new_n305_), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n578_), .B(KEYINPUT42), .Z(new_n579_));
  NAND3_X1  g378(.A1(new_n557_), .A2(new_n577_), .A3(new_n305_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(G1327gat));
  INV_X1    g380(.A(new_n553_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n458_), .A2(new_n582_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n546_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(G29gat), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(new_n585_), .A3(new_n362_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT102), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT43), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n588_), .B1(new_n384_), .B2(new_n552_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n552_), .ZN(new_n590_));
  AOI211_X1 g389(.A(KEYINPUT43), .B(new_n590_), .C1(new_n379_), .C2(new_n383_), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n528_), .B(new_n553_), .C1(new_n589_), .C2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT44), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n297_), .A2(new_n298_), .A3(new_n246_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n245_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n363_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(KEYINPUT98), .B1(new_n597_), .B2(new_n380_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n598_), .A2(new_n364_), .A3(new_n375_), .ZN(new_n599_));
  AOI22_X1  g398(.A1(new_n599_), .A2(new_n243_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n600_));
  OAI21_X1  g399(.A(KEYINPUT43), .B1(new_n600_), .B2(new_n590_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n384_), .A2(new_n588_), .A3(new_n552_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n603_), .A2(KEYINPUT44), .A3(new_n528_), .A4(new_n553_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n594_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(new_n362_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n587_), .B1(new_n606_), .B2(G29gat), .ZN(new_n607_));
  AOI211_X1 g406(.A(KEYINPUT102), .B(new_n585_), .C1(new_n605_), .C2(new_n362_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n586_), .B1(new_n607_), .B2(new_n608_), .ZN(G1328gat));
  INV_X1    g408(.A(G36gat), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n584_), .A2(new_n610_), .A3(new_n380_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT45), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n594_), .A2(new_n604_), .A3(new_n380_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT103), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(G36gat), .B1(new_n613_), .B2(new_n614_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n612_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  OAI221_X1 g418(.A(new_n612_), .B1(KEYINPUT104), .B2(KEYINPUT46), .C1(new_n615_), .C2(new_n616_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(G1329gat));
  NAND3_X1  g420(.A1(new_n594_), .A2(new_n604_), .A3(new_n571_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(G43gat), .ZN(new_n623_));
  INV_X1    g422(.A(G43gat), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n584_), .A2(new_n624_), .A3(new_n571_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(G1330gat));
  AOI21_X1  g427(.A(G50gat), .B1(new_n584_), .B2(new_n305_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n305_), .A2(G50gat), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n605_), .B2(new_n630_), .ZN(G1331gat));
  NOR2_X1   g430(.A1(new_n503_), .A2(new_n504_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n527_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n634_), .A2(new_n384_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(new_n554_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(G57gat), .B1(new_n637_), .B2(new_n362_), .ZN(new_n638_));
  NOR4_X1   g437(.A1(new_n459_), .A2(new_n633_), .A3(new_n632_), .A4(new_n553_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n362_), .A2(KEYINPUT106), .A3(G57gat), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n640_), .B1(KEYINPUT106), .B2(G57gat), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n638_), .B1(new_n639_), .B2(new_n641_), .ZN(G1332gat));
  NAND3_X1  g441(.A1(new_n637_), .A2(new_n462_), .A3(new_n380_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n639_), .A2(new_n380_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(G64gat), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n645_), .A2(KEYINPUT48), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(KEYINPUT48), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n643_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT107), .ZN(G1333gat));
  INV_X1    g448(.A(G71gat), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n650_), .B1(new_n639_), .B2(new_n571_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT49), .Z(new_n652_));
  NAND3_X1  g451(.A1(new_n637_), .A2(new_n650_), .A3(new_n571_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1334gat));
  NAND2_X1  g453(.A1(new_n639_), .A2(new_n305_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(G78gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT50), .ZN(new_n657_));
  INV_X1    g456(.A(new_n305_), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n658_), .A2(G78gat), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n657_), .B1(new_n636_), .B2(new_n659_), .ZN(G1335gat));
  NAND3_X1  g459(.A1(new_n603_), .A2(new_n553_), .A3(new_n634_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G85gat), .B1(new_n661_), .B2(new_n363_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n635_), .A2(new_n583_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n664_), .A2(new_n358_), .A3(new_n362_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n662_), .A2(new_n665_), .ZN(G1336gat));
  OAI21_X1  g465(.A(G92gat), .B1(new_n661_), .B2(new_n345_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n664_), .A2(new_n410_), .A3(new_n380_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1337gat));
  OAI21_X1  g468(.A(G99gat), .B1(new_n661_), .B2(new_n243_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n571_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n670_), .B1(new_n663_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT51), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n673_), .A2(KEYINPUT108), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n672_), .B(new_n674_), .ZN(G1338gat));
  INV_X1    g474(.A(KEYINPUT52), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n603_), .A2(new_n305_), .A3(new_n553_), .A4(new_n634_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n677_), .A2(new_n678_), .A3(G106gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n678_), .B1(new_n677_), .B2(G106gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n676_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n677_), .A2(G106gat), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT109), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n677_), .A2(new_n678_), .A3(G106gat), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n683_), .A2(KEYINPUT52), .A3(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n664_), .A2(new_n404_), .A3(new_n305_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n681_), .A2(new_n685_), .A3(new_n686_), .ZN(new_n687_));
  XOR2_X1   g486(.A(KEYINPUT110), .B(KEYINPUT53), .Z(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n688_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n681_), .A2(new_n685_), .A3(new_n686_), .A4(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(G1339gat));
  INV_X1    g491(.A(KEYINPUT118), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n582_), .A2(new_n527_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT111), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n695_), .A2(new_n590_), .A3(new_n500_), .A4(new_n501_), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT54), .Z(new_n697_));
  NAND2_X1  g496(.A1(new_n512_), .A2(new_n513_), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n521_), .B(new_n698_), .C1(new_n515_), .C2(new_n513_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n522_), .A2(new_n496_), .A3(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT55), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n486_), .A2(new_n488_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n482_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n461_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n701_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n489_), .A2(KEYINPUT55), .A3(new_n461_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n704_), .A2(new_n705_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n706_), .A2(new_n707_), .A3(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n497_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT56), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n709_), .A2(KEYINPUT56), .A3(new_n710_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n700_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT58), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT117), .ZN(new_n717_));
  XOR2_X1   g516(.A(KEYINPUT116), .B(KEYINPUT58), .Z(new_n718_));
  OAI21_X1  g517(.A(new_n552_), .B1(new_n715_), .B2(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n527_), .B1(new_n490_), .B2(new_n495_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT112), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n489_), .A2(KEYINPUT55), .A3(new_n461_), .ZN(new_n724_));
  AOI21_X1  g523(.A(KEYINPUT55), .B1(new_n489_), .B2(new_n461_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n489_), .A2(new_n461_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n724_), .A2(new_n725_), .A3(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n723_), .B1(new_n727_), .B2(new_n497_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT114), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n709_), .A2(KEYINPUT112), .A3(new_n710_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(KEYINPUT113), .B(KEYINPUT56), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n728_), .A2(new_n729_), .A3(new_n730_), .A4(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n714_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n731_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n734_), .B1(new_n711_), .B2(new_n723_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n729_), .B1(new_n735_), .B2(new_n730_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n722_), .B1(new_n733_), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT115), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT115), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n739_), .B(new_n722_), .C1(new_n733_), .C2(new_n736_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n498_), .A2(new_n522_), .A3(new_n699_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n738_), .A2(new_n740_), .A3(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT57), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n742_), .A2(new_n743_), .A3(new_n458_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n742_), .B2(new_n458_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n721_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n541_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n697_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n381_), .A2(new_n362_), .A3(new_n571_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n693_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n697_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n742_), .A2(new_n458_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT57), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n742_), .A2(new_n743_), .A3(new_n458_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n720_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n755_), .B2(new_n541_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n749_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(KEYINPUT118), .A3(new_n757_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n750_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(G113gat), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n759_), .A2(new_n760_), .A3(new_n633_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT119), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT59), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n763_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n697_), .B1(new_n746_), .B2(new_n553_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n749_), .A2(KEYINPUT59), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n765_), .A2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n762_), .B1(new_n764_), .B2(new_n768_), .ZN(new_n769_));
  OR2_X1    g568(.A1(new_n765_), .A2(new_n767_), .ZN(new_n770_));
  OAI21_X1  g569(.A(KEYINPUT59), .B1(new_n748_), .B2(new_n749_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n770_), .A2(new_n771_), .A3(KEYINPUT119), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n769_), .A2(new_n772_), .A3(new_n633_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n761_), .B1(new_n773_), .B2(new_n760_), .ZN(G1340gat));
  INV_X1    g573(.A(new_n632_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT60), .ZN(new_n776_));
  INV_X1    g575(.A(G120gat), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n775_), .A2(new_n776_), .A3(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n778_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n759_), .A2(new_n779_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n764_), .A2(new_n768_), .A3(new_n632_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n777_), .B2(new_n781_), .ZN(G1341gat));
  INV_X1    g581(.A(G127gat), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n747_), .A2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n769_), .A2(new_n772_), .A3(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n750_), .A2(new_n758_), .A3(new_n582_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n783_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n785_), .A2(KEYINPUT120), .A3(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT120), .B1(new_n785_), .B2(new_n787_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(G1342gat));
  INV_X1    g589(.A(G134gat), .ZN(new_n791_));
  INV_X1    g590(.A(new_n458_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n759_), .A2(new_n791_), .A3(new_n792_), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n769_), .A2(new_n772_), .A3(new_n552_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(new_n794_), .B2(new_n791_), .ZN(G1343gat));
  NAND4_X1  g594(.A1(new_n305_), .A2(new_n362_), .A3(new_n345_), .A4(new_n243_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n748_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n633_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n775_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(KEYINPUT121), .B(G148gat), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n800_), .B(new_n801_), .ZN(G1345gat));
  NAND2_X1  g601(.A1(new_n797_), .A2(new_n582_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(KEYINPUT122), .ZN(new_n804_));
  XOR2_X1   g603(.A(KEYINPUT61), .B(G155gat), .Z(new_n805_));
  XNOR2_X1  g604(.A(new_n804_), .B(new_n805_), .ZN(G1346gat));
  NAND2_X1  g605(.A1(new_n797_), .A2(new_n552_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n458_), .A2(G162gat), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n807_), .A2(G162gat), .B1(new_n797_), .B2(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT123), .ZN(G1347gat));
  NAND2_X1  g609(.A1(new_n380_), .A2(new_n382_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n765_), .A2(new_n305_), .A3(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n633_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(new_n308_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(G169gat), .ZN(new_n815_));
  XNOR2_X1  g614(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n814_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n815_), .B2(new_n816_), .ZN(G1348gat));
  NAND2_X1  g617(.A1(new_n756_), .A2(new_n658_), .ZN(new_n819_));
  INV_X1    g618(.A(G176gat), .ZN(new_n820_));
  NOR4_X1   g619(.A1(new_n819_), .A2(new_n820_), .A3(new_n632_), .A4(new_n811_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n309_), .B1(new_n812_), .B2(new_n775_), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n822_), .A2(KEYINPUT125), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(KEYINPUT125), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n821_), .B1(new_n823_), .B2(new_n824_), .ZN(G1349gat));
  OR3_X1    g624(.A1(new_n819_), .A2(new_n553_), .A3(new_n811_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n747_), .A2(new_n220_), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n826_), .A2(new_n206_), .B1(new_n812_), .B2(new_n827_), .ZN(G1350gat));
  NAND3_X1  g627(.A1(new_n812_), .A2(new_n792_), .A3(new_n221_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n812_), .A2(new_n552_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n207_), .ZN(G1351gat));
  NAND3_X1  g630(.A1(new_n377_), .A2(new_n380_), .A3(new_n243_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n748_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n633_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g634(.A(KEYINPUT126), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n632_), .B1(new_n836_), .B2(G204gat), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n833_), .A2(new_n837_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(KEYINPUT127), .ZN(new_n839_));
  OR2_X1    g638(.A1(new_n836_), .A2(G204gat), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n839_), .B(new_n840_), .ZN(G1353gat));
  INV_X1    g640(.A(KEYINPUT63), .ZN(new_n842_));
  INV_X1    g641(.A(G211gat), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n833_), .B(new_n541_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n843_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(G1354gat));
  INV_X1    g645(.A(G218gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n833_), .A2(new_n847_), .A3(new_n792_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n748_), .A2(new_n590_), .A3(new_n832_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(new_n847_), .ZN(G1355gat));
endmodule


