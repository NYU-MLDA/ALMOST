//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n869_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n917_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n928_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  XOR2_X1   g001(.A(G57gat), .B(G64gat), .Z(new_n203_));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(G71gat), .B(G78gat), .Z(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT68), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT68), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n205_), .A2(new_n209_), .A3(new_n206_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n203_), .A2(new_n204_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n208_), .A2(new_n212_), .A3(new_n210_), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G85gat), .Z(new_n217_));
  INV_X1    g016(.A(KEYINPUT9), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(new_n218_), .A3(G92gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G85gat), .B(G92gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n219_), .B1(new_n218_), .B2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT66), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT10), .B(G99gat), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n223_), .A2(G106gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G99gat), .A2(G106gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT6), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n229_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n219_), .B(new_n231_), .C1(new_n218_), .C2(new_n220_), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n222_), .A2(new_n226_), .A3(new_n230_), .A4(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(G99gat), .A2(G106gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT7), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n220_), .B1(new_n235_), .B2(new_n228_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(KEYINPUT67), .A2(KEYINPUT8), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n233_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n239_), .B1(new_n233_), .B2(new_n238_), .ZN(new_n242_));
  OAI211_X1 g041(.A(KEYINPUT12), .B(new_n216_), .C1(new_n241_), .C2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G230gat), .A2(G233gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n233_), .A2(new_n238_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n216_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT12), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n245_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n214_), .A2(new_n215_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n243_), .A2(new_n244_), .A3(new_n248_), .A4(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n246_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n216_), .A2(new_n245_), .ZN(new_n254_));
  OAI211_X1 g053(.A(G230gat), .B(G233gat), .C1(new_n253_), .C2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G120gat), .B(G148gat), .ZN(new_n256_));
  INV_X1    g055(.A(G204gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT5), .B(G176gat), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n258_), .B(new_n259_), .Z(new_n260_));
  NAND3_X1  g059(.A1(new_n252_), .A2(new_n255_), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n260_), .B1(new_n252_), .B2(new_n255_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n202_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n252_), .A2(new_n255_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n260_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n267_), .A2(KEYINPUT13), .A3(new_n261_), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n264_), .A2(new_n268_), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n269_), .A2(KEYINPUT70), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(KEYINPUT70), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G29gat), .B(G36gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(G50gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT71), .B(G43gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(G50gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n273_), .B(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n275_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n276_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G15gat), .B(G22gat), .ZN(new_n282_));
  INV_X1    g081(.A(G1gat), .ZN(new_n283_));
  INV_X1    g082(.A(G8gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT14), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G1gat), .B(G8gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n281_), .A2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n281_), .A2(new_n288_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G229gat), .A2(G233gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT76), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  AND3_X1   g092(.A1(new_n276_), .A2(new_n280_), .A3(KEYINPUT15), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT15), .B1(new_n276_), .B2(new_n280_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n288_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n290_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n296_), .A2(new_n292_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT76), .ZN(new_n299_));
  INV_X1    g098(.A(new_n292_), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n299_), .B(new_n300_), .C1(new_n289_), .C2(new_n290_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G113gat), .B(G141gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G169gat), .B(G197gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n293_), .A2(new_n298_), .A3(new_n301_), .A4(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n293_), .A2(new_n298_), .A3(new_n301_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT77), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT77), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n293_), .A2(new_n310_), .A3(new_n298_), .A4(new_n301_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(new_n311_), .A3(new_n304_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT78), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n307_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n309_), .A2(KEYINPUT78), .A3(new_n311_), .A4(new_n304_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n272_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT87), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT85), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G127gat), .A2(G134gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(G127gat), .A2(G134gat), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n319_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  OR2_X1    g122(.A1(G127gat), .A2(G134gat), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n324_), .A2(KEYINPUT85), .A3(new_n320_), .ZN(new_n325_));
  AND2_X1   g124(.A1(G113gat), .A2(G120gat), .ZN(new_n326_));
  NOR2_X1   g125(.A1(G113gat), .A2(G120gat), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT86), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(G113gat), .ZN(new_n329_));
  INV_X1    g128(.A(G120gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT86), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G113gat), .A2(G120gat), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n331_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  AND4_X1   g133(.A1(new_n323_), .A2(new_n325_), .A3(new_n328_), .A4(new_n334_), .ZN(new_n335_));
  AOI22_X1  g134(.A1(new_n323_), .A2(new_n325_), .B1(new_n328_), .B2(new_n334_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n318_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n323_), .A2(new_n325_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n328_), .A2(new_n334_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n318_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n337_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT31), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT84), .ZN(new_n344_));
  INV_X1    g143(.A(G43gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G227gat), .A2(G233gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT79), .B(G190gat), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n349_), .B1(new_n350_), .B2(KEYINPUT26), .ZN(new_n351_));
  XOR2_X1   g150(.A(KEYINPUT25), .B(G183gat), .Z(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(G169gat), .ZN(new_n354_));
  INV_X1    g153(.A(G176gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  OR2_X1    g155(.A1(new_n356_), .A2(KEYINPUT24), .ZN(new_n357_));
  INV_X1    g156(.A(G183gat), .ZN(new_n358_));
  INV_X1    g157(.A(G190gat), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT23), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT23), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n361_), .A2(G183gat), .A3(G190gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G169gat), .A2(G176gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT80), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n356_), .A2(KEYINPUT24), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n357_), .B(new_n363_), .C1(new_n365_), .C2(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n353_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n365_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n360_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT83), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n362_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n362_), .A2(new_n371_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n370_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n350_), .A2(G183gat), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n369_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n354_), .A2(KEYINPUT81), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n354_), .A2(KEYINPUT81), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT22), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT82), .ZN(new_n381_));
  OR2_X1    g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT22), .ZN(new_n383_));
  AOI21_X1  g182(.A(G176gat), .B1(new_n383_), .B2(G169gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n380_), .A2(new_n381_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n382_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n368_), .B1(new_n377_), .B2(new_n386_), .ZN(new_n387_));
  XOR2_X1   g186(.A(KEYINPUT30), .B(G15gat), .Z(new_n388_));
  XNOR2_X1  g187(.A(G71gat), .B(G99gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  XOR2_X1   g189(.A(new_n387_), .B(new_n390_), .Z(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n348_), .A2(new_n392_), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n346_), .A2(new_n347_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n346_), .A2(new_n347_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n394_), .A2(new_n395_), .A3(new_n391_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n393_), .A2(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(G141gat), .A2(G148gat), .ZN(new_n398_));
  AND2_X1   g197(.A1(G141gat), .A2(G148gat), .ZN(new_n399_));
  NOR2_X1   g198(.A1(G155gat), .A2(G162gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G155gat), .A2(G162gat), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n400_), .B1(KEYINPUT1), .B2(new_n401_), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n401_), .A2(KEYINPUT1), .ZN(new_n403_));
  AOI211_X1 g202(.A(new_n398_), .B(new_n399_), .C1(new_n402_), .C2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  OR2_X1    g204(.A1(KEYINPUT89), .A2(KEYINPUT2), .ZN(new_n406_));
  NAND2_X1  g205(.A1(KEYINPUT88), .A2(KEYINPUT3), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n406_), .A2(new_n399_), .B1(new_n398_), .B2(new_n407_), .ZN(new_n408_));
  OR2_X1    g207(.A1(G141gat), .A2(G148gat), .ZN(new_n409_));
  INV_X1    g208(.A(new_n407_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(KEYINPUT88), .A2(KEYINPUT3), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n409_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G141gat), .A2(G148gat), .ZN(new_n413_));
  AND2_X1   g212(.A1(KEYINPUT89), .A2(KEYINPUT2), .ZN(new_n414_));
  NOR2_X1   g213(.A1(KEYINPUT89), .A2(KEYINPUT2), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n413_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n408_), .A2(new_n412_), .A3(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT90), .ZN(new_n418_));
  XOR2_X1   g217(.A(G155gat), .B(G162gat), .Z(new_n419_));
  AND3_X1   g218(.A1(new_n417_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n418_), .B1(new_n417_), .B2(new_n419_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n405_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n422_), .A2(KEYINPUT29), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT28), .ZN(new_n424_));
  XOR2_X1   g223(.A(G22gat), .B(G50gat), .Z(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G78gat), .B(G106gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(KEYINPUT96), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G211gat), .B(G218gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G197gat), .B(G204gat), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT21), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n431_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT93), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT92), .ZN(new_n436_));
  INV_X1    g235(.A(G197gat), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n437_), .A3(G204gat), .ZN(new_n438_));
  AOI21_X1  g237(.A(KEYINPUT92), .B1(new_n257_), .B2(G197gat), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n257_), .A2(G197gat), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n433_), .B(new_n438_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n434_), .B1(new_n435_), .B2(new_n441_), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n441_), .A2(new_n435_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n431_), .A2(new_n433_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n438_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n444_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT94), .ZN(new_n449_));
  AOI22_X1  g248(.A1(new_n442_), .A2(new_n443_), .B1(new_n446_), .B2(new_n445_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT94), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n449_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G228gat), .A2(G233gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT91), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n456_), .B1(new_n422_), .B2(KEYINPUT29), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n453_), .A2(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n458_), .A2(KEYINPUT95), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(KEYINPUT95), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n450_), .B1(new_n422_), .B2(KEYINPUT29), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n462_), .A2(new_n455_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n430_), .B1(new_n461_), .B2(new_n464_), .ZN(new_n465_));
  AOI211_X1 g264(.A(new_n429_), .B(new_n463_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n427_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n460_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n458_), .A2(KEYINPUT95), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n464_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n429_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n461_), .A2(new_n430_), .A3(new_n464_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n426_), .A3(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n467_), .A2(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(G1gat), .B(G29gat), .Z(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(G85gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT0), .B(G57gat), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n476_), .B(new_n477_), .Z(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT100), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n338_), .A2(new_n339_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n323_), .A2(new_n325_), .A3(new_n328_), .A4(new_n334_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n340_), .B1(new_n483_), .B2(new_n318_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n422_), .A2(new_n484_), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n405_), .B(new_n483_), .C1(new_n420_), .C2(new_n421_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n480_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n480_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G225gat), .A2(G233gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT101), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n479_), .B1(new_n490_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT102), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT4), .B1(new_n487_), .B2(new_n489_), .ZN(new_n496_));
  AOI21_X1  g295(.A(KEYINPUT4), .B1(new_n422_), .B2(new_n484_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n495_), .B1(new_n499_), .B2(new_n491_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n491_), .ZN(new_n501_));
  AOI211_X1 g300(.A(KEYINPUT102), .B(new_n501_), .C1(new_n496_), .C2(new_n498_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n494_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT103), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n490_), .A2(new_n491_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n417_), .A2(new_n419_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT90), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n417_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n404_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n486_), .B1(new_n509_), .B2(new_n342_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT100), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n488_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n497_), .B1(new_n512_), .B2(KEYINPUT4), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n505_), .B(new_n479_), .C1(new_n513_), .C2(new_n492_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT33), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n492_), .B1(new_n496_), .B2(new_n498_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT33), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n517_), .A2(new_n518_), .A3(new_n505_), .A4(new_n479_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n515_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G226gat), .A2(G233gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT19), .ZN(new_n522_));
  INV_X1    g321(.A(new_n387_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n453_), .A2(new_n523_), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n360_), .A2(new_n362_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n354_), .A2(KEYINPUT22), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n384_), .A2(new_n527_), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n526_), .A2(new_n369_), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT97), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n526_), .A2(new_n369_), .A3(new_n528_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT97), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n356_), .A2(KEYINPUT24), .A3(new_n364_), .ZN(new_n534_));
  XOR2_X1   g333(.A(KEYINPUT26), .B(G190gat), .Z(new_n535_));
  OAI211_X1 g334(.A(new_n357_), .B(new_n534_), .C1(new_n352_), .C2(new_n535_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n536_), .A2(new_n374_), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n530_), .A2(new_n533_), .A3(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT20), .B1(new_n538_), .B2(new_n450_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n522_), .B1(new_n524_), .B2(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n387_), .B1(new_n449_), .B2(new_n452_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n522_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n530_), .A2(new_n533_), .A3(new_n537_), .ZN(new_n543_));
  OAI211_X1 g342(.A(KEYINPUT20), .B(new_n542_), .C1(new_n543_), .C2(new_n448_), .ZN(new_n544_));
  OAI21_X1  g343(.A(KEYINPUT98), .B1(new_n541_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n453_), .A2(new_n523_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n542_), .A2(KEYINPUT20), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n547_), .B1(new_n538_), .B2(new_n450_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT98), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n546_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n540_), .A2(new_n545_), .A3(new_n550_), .ZN(new_n551_));
  XOR2_X1   g350(.A(KEYINPUT99), .B(KEYINPUT18), .Z(new_n552_));
  XNOR2_X1  g351(.A(G8gat), .B(G36gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G64gat), .B(G92gat), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n554_), .B(new_n555_), .Z(new_n556_));
  NAND2_X1  g355(.A1(new_n551_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n556_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n540_), .A2(new_n545_), .A3(new_n550_), .A4(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT103), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n562_), .B(new_n494_), .C1(new_n500_), .C2(new_n502_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n504_), .A2(new_n520_), .A3(new_n561_), .A4(new_n563_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n558_), .A2(KEYINPUT32), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n551_), .A2(new_n565_), .ZN(new_n566_));
  OAI221_X1 g365(.A(KEYINPUT20), .B1(new_n538_), .B2(new_n450_), .C1(new_n453_), .C2(new_n523_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n567_), .A2(new_n522_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n537_), .A2(KEYINPUT104), .A3(new_n531_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT104), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n536_), .A2(new_n374_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n571_), .B1(new_n529_), .B2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n570_), .A2(new_n573_), .A3(new_n450_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(KEYINPUT20), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n575_), .A2(KEYINPUT105), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n541_), .B1(KEYINPUT105), .B2(new_n575_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n569_), .B1(new_n578_), .B2(new_n542_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n566_), .B1(new_n579_), .B2(new_n565_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n505_), .ZN(new_n581_));
  OAI211_X1 g380(.A(KEYINPUT106), .B(new_n478_), .C1(new_n516_), .C2(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n478_), .B1(new_n516_), .B2(new_n581_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT106), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n583_), .A2(new_n514_), .A3(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n580_), .A2(new_n582_), .A3(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n474_), .B1(new_n564_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT27), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n559_), .A2(KEYINPUT27), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n542_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n556_), .B1(new_n590_), .B2(new_n568_), .ZN(new_n591_));
  AOI22_X1  g390(.A1(new_n588_), .A2(new_n560_), .B1(new_n589_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n585_), .A2(new_n582_), .ZN(new_n593_));
  AND3_X1   g392(.A1(new_n474_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n397_), .B1(new_n587_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n397_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n592_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n597_), .A2(new_n474_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n596_), .A2(new_n598_), .A3(new_n593_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n317_), .B1(new_n595_), .B2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G232gat), .A2(G233gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT34), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT35), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  OAI22_X1  g405(.A1(new_n245_), .A2(new_n281_), .B1(KEYINPUT35), .B2(new_n602_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n241_), .A2(new_n242_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n294_), .A2(new_n295_), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n606_), .B(new_n608_), .C1(new_n609_), .C2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n245_), .A2(KEYINPUT69), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n610_), .B1(new_n612_), .B2(new_n240_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n605_), .B1(new_n613_), .B2(new_n607_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT74), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(G134gat), .B(G162gat), .Z(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT72), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G190gat), .B(G218gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT36), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n611_), .A2(new_n614_), .A3(KEYINPUT74), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n617_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT37), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT36), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n621_), .A2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT73), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n611_), .A2(new_n614_), .A3(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n624_), .A2(new_n625_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT75), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n615_), .A2(new_n622_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n629_), .ZN(new_n633_));
  OAI21_X1  g432(.A(KEYINPUT37), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n630_), .A2(new_n631_), .A3(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n631_), .B1(new_n630_), .B2(new_n634_), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(G231gat), .A2(G233gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n288_), .B(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n250_), .B(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(G127gat), .B(G155gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(G211gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(KEYINPUT16), .B(G183gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT17), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n640_), .A2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n644_), .B(KEYINPUT17), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n646_), .B1(new_n640_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n637_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n600_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n593_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n653_), .A2(new_n283_), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT38), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n624_), .A2(new_n629_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n659_), .A2(new_n650_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n600_), .A2(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G1gat), .B1(new_n661_), .B2(new_n593_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n655_), .A2(new_n656_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n657_), .A2(new_n662_), .A3(new_n663_), .ZN(G1324gat));
  NAND3_X1  g463(.A1(new_n653_), .A2(new_n284_), .A3(new_n597_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G8gat), .B1(new_n661_), .B2(new_n592_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n666_), .A2(KEYINPUT39), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(KEYINPUT39), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n665_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT40), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  OAI211_X1 g470(.A(KEYINPUT40), .B(new_n665_), .C1(new_n667_), .C2(new_n668_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1325gat));
  OAI21_X1  g472(.A(G15gat), .B1(new_n661_), .B2(new_n397_), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n674_), .A2(KEYINPUT41), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(KEYINPUT41), .ZN(new_n676_));
  OR3_X1    g475(.A1(new_n652_), .A2(G15gat), .A3(new_n397_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n675_), .A2(new_n676_), .A3(new_n677_), .ZN(G1326gat));
  INV_X1    g477(.A(new_n474_), .ZN(new_n679_));
  OAI21_X1  g478(.A(G22gat), .B1(new_n661_), .B2(new_n679_), .ZN(new_n680_));
  XOR2_X1   g479(.A(KEYINPUT107), .B(KEYINPUT42), .Z(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n679_), .A2(G22gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n682_), .B1(new_n652_), .B2(new_n683_), .ZN(G1327gat));
  NOR2_X1   g483(.A1(new_n658_), .A2(new_n649_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n600_), .A2(new_n685_), .ZN(new_n686_));
  OR3_X1    g485(.A1(new_n686_), .A2(G29gat), .A3(new_n593_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n650_), .B1(KEYINPUT108), .B2(KEYINPUT44), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n317_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n595_), .A2(new_n599_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n691_), .B2(new_n637_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n635_), .A2(new_n636_), .ZN(new_n693_));
  AOI211_X1 g492(.A(KEYINPUT43), .B(new_n693_), .C1(new_n595_), .C2(new_n599_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n689_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT108), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n695_), .A2(new_n698_), .ZN(new_n699_));
  OAI221_X1 g498(.A(new_n689_), .B1(new_n696_), .B2(new_n697_), .C1(new_n692_), .C2(new_n694_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n593_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n701_), .A2(KEYINPUT109), .ZN(new_n702_));
  OAI21_X1  g501(.A(G29gat), .B1(new_n701_), .B2(KEYINPUT109), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n687_), .B1(new_n702_), .B2(new_n703_), .ZN(G1328gat));
  INV_X1    g503(.A(G36gat), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n600_), .A2(new_n705_), .A3(new_n597_), .A4(new_n685_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT45), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n592_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n707_), .B1(new_n708_), .B2(new_n705_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT46), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  OAI211_X1 g510(.A(KEYINPUT46), .B(new_n707_), .C1(new_n708_), .C2(new_n705_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1329gat));
  NAND3_X1  g512(.A1(new_n600_), .A2(new_n596_), .A3(new_n685_), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n714_), .A2(KEYINPUT110), .A3(new_n345_), .ZN(new_n715_));
  AOI21_X1  g514(.A(KEYINPUT110), .B1(new_n714_), .B2(new_n345_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n596_), .A2(G43gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT47), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT47), .B1(new_n717_), .B2(new_n719_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1330gat));
  AOI21_X1  g523(.A(new_n679_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n474_), .A2(new_n277_), .ZN(new_n726_));
  OAI22_X1  g525(.A1(new_n725_), .A2(new_n277_), .B1(new_n686_), .B2(new_n726_), .ZN(G1331gat));
  AOI211_X1 g526(.A(new_n316_), .B(new_n272_), .C1(new_n595_), .C2(new_n599_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n660_), .ZN(new_n729_));
  INV_X1    g528(.A(G57gat), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n729_), .A2(new_n730_), .A3(new_n593_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n728_), .A2(new_n651_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(new_n654_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n731_), .B1(new_n730_), .B2(new_n734_), .ZN(G1332gat));
  OAI21_X1  g534(.A(G64gat), .B1(new_n729_), .B2(new_n592_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT48), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n592_), .A2(G64gat), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT111), .Z(new_n739_));
  OAI21_X1  g538(.A(new_n737_), .B1(new_n732_), .B2(new_n739_), .ZN(G1333gat));
  NAND3_X1  g539(.A1(new_n728_), .A2(new_n596_), .A3(new_n660_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT49), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n741_), .A2(new_n742_), .A3(G71gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n741_), .B2(G71gat), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n397_), .A2(G71gat), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT112), .Z(new_n746_));
  OAI22_X1  g545(.A1(new_n743_), .A2(new_n744_), .B1(new_n732_), .B2(new_n746_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT113), .ZN(G1334gat));
  OAI21_X1  g547(.A(G78gat), .B1(new_n729_), .B2(new_n679_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT50), .ZN(new_n750_));
  OR2_X1    g549(.A1(new_n679_), .A2(G78gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n732_), .B2(new_n751_), .ZN(G1335gat));
  NAND2_X1  g551(.A1(new_n728_), .A2(new_n685_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(G85gat), .B1(new_n754_), .B2(new_n654_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n272_), .A2(new_n316_), .A3(new_n649_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n756_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n654_), .A2(new_n217_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(G1336gat));
  AOI21_X1  g559(.A(G92gat), .B1(new_n754_), .B2(new_n597_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n597_), .A2(G92gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n758_), .B2(new_n762_), .ZN(G1337gat));
  OAI21_X1  g562(.A(G99gat), .B1(new_n757_), .B2(new_n397_), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n397_), .A2(new_n223_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n753_), .B2(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT51), .ZN(G1338gat));
  OR3_X1    g566(.A1(new_n753_), .A2(G106gat), .A3(new_n679_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n474_), .B(new_n756_), .C1(new_n692_), .C2(new_n694_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n769_), .A2(new_n770_), .A3(G106gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n769_), .B2(G106gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT53), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n775_), .B(new_n768_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1339gat));
  NAND3_X1  g576(.A1(new_n296_), .A2(new_n300_), .A3(new_n297_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n778_), .B(new_n304_), .C1(new_n300_), .C2(new_n291_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n306_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n261_), .A2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT116), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n254_), .B1(new_n247_), .B2(new_n246_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n244_), .B1(new_n783_), .B2(new_n243_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n252_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n783_), .A2(KEYINPUT55), .A3(new_n244_), .A4(new_n243_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n266_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT56), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n788_), .A2(KEYINPUT56), .A3(new_n266_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n782_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT117), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT58), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT58), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT56), .B1(new_n788_), .B2(new_n266_), .ZN(new_n797_));
  AOI211_X1 g596(.A(new_n790_), .B(new_n260_), .C1(new_n786_), .C2(new_n787_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  OAI211_X1 g598(.A(KEYINPUT117), .B(new_n796_), .C1(new_n799_), .C2(new_n782_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n795_), .A2(new_n637_), .A3(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n262_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n802_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n780_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n658_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n805_), .A2(KEYINPUT57), .A3(new_n658_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n801_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n264_), .A2(new_n268_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n312_), .A2(new_n313_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n813_), .A2(new_n315_), .A3(new_n306_), .A4(new_n649_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n812_), .B1(KEYINPUT114), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n314_), .A2(new_n816_), .A3(new_n315_), .A4(new_n649_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n811_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n814_), .A2(KEYINPUT114), .ZN(new_n819_));
  AND4_X1   g618(.A1(new_n811_), .A2(new_n819_), .A3(new_n269_), .A4(new_n817_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n693_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT54), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n823_), .B(new_n693_), .C1(new_n818_), .C2(new_n820_), .ZN(new_n824_));
  AOI22_X1  g623(.A1(new_n810_), .A2(new_n650_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n598_), .A2(new_n654_), .A3(new_n596_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(G113gat), .B1(new_n827_), .B2(new_n316_), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT59), .B1(new_n825_), .B2(new_n826_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT59), .ZN(new_n830_));
  INV_X1    g629(.A(new_n826_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n822_), .A2(new_n824_), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT57), .B1(new_n805_), .B2(new_n658_), .ZN(new_n833_));
  AOI211_X1 g632(.A(new_n807_), .B(new_n659_), .C1(new_n803_), .C2(new_n804_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n649_), .B1(new_n835_), .B2(new_n801_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n830_), .B(new_n831_), .C1(new_n832_), .C2(new_n836_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n829_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n329_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n828_), .B1(new_n838_), .B2(new_n839_), .ZN(G1340gat));
  INV_X1    g639(.A(new_n272_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n829_), .A2(new_n837_), .A3(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(G120gat), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n330_), .B1(new_n272_), .B2(KEYINPUT60), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n827_), .B(new_n844_), .C1(KEYINPUT60), .C2(new_n330_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(G1341gat));
  NOR2_X1   g645(.A1(new_n650_), .A2(KEYINPUT118), .ZN(new_n847_));
  MUX2_X1   g646(.A(KEYINPUT118), .B(new_n847_), .S(G127gat), .Z(new_n848_));
  NAND3_X1  g647(.A1(new_n829_), .A2(new_n837_), .A3(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n810_), .A2(new_n650_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n822_), .A2(new_n824_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n852_), .A2(new_n649_), .A3(new_n831_), .ZN(new_n853_));
  INV_X1    g652(.A(G127gat), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n849_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n849_), .A2(new_n855_), .A3(KEYINPUT119), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(G1342gat));
  AOI21_X1  g659(.A(G134gat), .B1(new_n827_), .B2(new_n659_), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n637_), .A2(G134gat), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n861_), .B1(new_n838_), .B2(new_n862_), .ZN(G1343gat));
  NAND4_X1  g662(.A1(new_n397_), .A2(new_n474_), .A3(new_n654_), .A4(new_n592_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(KEYINPUT120), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n852_), .A2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n316_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n841_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g669(.A1(new_n852_), .A2(new_n649_), .A3(new_n865_), .ZN(new_n871_));
  XOR2_X1   g670(.A(KEYINPUT121), .B(KEYINPUT122), .Z(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n872_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n852_), .A2(new_n649_), .A3(new_n865_), .A4(new_n874_), .ZN(new_n875_));
  XOR2_X1   g674(.A(KEYINPUT61), .B(G155gat), .Z(new_n876_));
  AND3_X1   g675(.A1(new_n873_), .A2(new_n875_), .A3(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n876_), .B1(new_n873_), .B2(new_n875_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(G1346gat));
  AOI21_X1  g678(.A(G162gat), .B1(new_n866_), .B2(new_n659_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n637_), .A2(G162gat), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n866_), .B2(new_n881_), .ZN(G1347gat));
  NOR2_X1   g681(.A1(new_n825_), .A2(new_n474_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n383_), .A2(G169gat), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n397_), .A2(new_n654_), .A3(new_n592_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n316_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NAND4_X1  g686(.A1(new_n883_), .A2(new_n884_), .A3(new_n527_), .A4(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n889_));
  XOR2_X1   g688(.A(new_n886_), .B(KEYINPUT123), .Z(new_n890_));
  NAND2_X1  g689(.A1(new_n883_), .A2(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n889_), .B1(new_n891_), .B2(G169gat), .ZN(new_n892_));
  AOI211_X1 g691(.A(KEYINPUT62), .B(new_n354_), .C1(new_n883_), .C2(new_n890_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n888_), .B1(new_n892_), .B2(new_n893_), .ZN(G1348gat));
  NAND3_X1  g693(.A1(new_n852_), .A2(new_n679_), .A3(new_n885_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n895_), .A2(new_n272_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(new_n355_), .ZN(G1349gat));
  NAND3_X1  g696(.A1(new_n883_), .A2(new_n649_), .A3(new_n885_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(G183gat), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n899_), .B1(new_n352_), .B2(new_n898_), .ZN(G1350gat));
  OAI21_X1  g699(.A(G190gat), .B1(new_n895_), .B2(new_n693_), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n658_), .A2(new_n535_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n895_), .B2(new_n902_), .ZN(G1351gat));
  NOR2_X1   g702(.A1(new_n679_), .A2(new_n654_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n904_), .A2(new_n597_), .A3(new_n397_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  OAI211_X1 g705(.A(new_n316_), .B(new_n906_), .C1(new_n832_), .C2(new_n836_), .ZN(new_n907_));
  OAI21_X1  g706(.A(KEYINPUT124), .B1(new_n907_), .B2(new_n437_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n825_), .A2(new_n905_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT124), .ZN(new_n910_));
  NAND4_X1  g709(.A1(new_n909_), .A2(new_n910_), .A3(G197gat), .A4(new_n316_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n908_), .A2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT125), .ZN(new_n913_));
  AND3_X1   g712(.A1(new_n907_), .A2(new_n913_), .A3(new_n437_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n913_), .B1(new_n907_), .B2(new_n437_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n912_), .A2(new_n914_), .A3(new_n915_), .ZN(G1352gat));
  NAND2_X1  g715(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n917_));
  XNOR2_X1  g716(.A(KEYINPUT126), .B(G204gat), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n909_), .A2(new_n841_), .ZN(new_n919_));
  MUX2_X1   g718(.A(new_n917_), .B(new_n918_), .S(new_n919_), .Z(G1353gat));
  NAND2_X1  g719(.A1(new_n909_), .A2(new_n649_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n922_));
  AND2_X1   g721(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n921_), .A2(new_n922_), .A3(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n924_), .B1(new_n921_), .B2(new_n922_), .ZN(G1354gat));
  AOI21_X1  g724(.A(G218gat), .B1(new_n909_), .B2(new_n659_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n637_), .A2(G218gat), .ZN(new_n927_));
  XOR2_X1   g726(.A(new_n927_), .B(KEYINPUT127), .Z(new_n928_));
  AOI21_X1  g727(.A(new_n926_), .B1(new_n909_), .B2(new_n928_), .ZN(G1355gat));
endmodule


