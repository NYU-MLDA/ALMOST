//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n800_, new_n801_, new_n803_,
    new_n804_, new_n805_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n913_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n947_,
    new_n948_, new_n950_, new_n951_, new_n952_, new_n954_, new_n955_,
    new_n957_, new_n959_, new_n960_, new_n961_, new_n962_, new_n964_,
    new_n965_, new_n966_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G64gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(G92gat), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT80), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT80), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(G183gat), .A3(G190gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(KEYINPUT79), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT79), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT23), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n215_), .A3(new_n207_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n212_), .A2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT22), .B(G169gat), .ZN(new_n222_));
  INV_X1    g021(.A(G176gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  AND3_X1   g023(.A1(new_n220_), .A2(new_n221_), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT95), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT82), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT79), .B(KEYINPUT23), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n227_), .B1(new_n228_), .B2(new_n207_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n208_), .A2(new_n210_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT23), .ZN(new_n231_));
  INV_X1    g030(.A(new_n207_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n214_), .A2(KEYINPUT23), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n211_), .A2(KEYINPUT79), .ZN(new_n234_));
  OAI211_X1 g033(.A(KEYINPUT82), .B(new_n232_), .C1(new_n233_), .C2(new_n234_), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n229_), .A2(new_n231_), .A3(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT24), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n239_), .A2(KEYINPUT94), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(KEYINPUT94), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n221_), .B(new_n238_), .C1(new_n240_), .C2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT26), .B(G190gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT25), .B(G183gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT94), .B(KEYINPUT24), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(new_n237_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n242_), .A2(new_n245_), .A3(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n226_), .B1(new_n236_), .B2(new_n248_), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n242_), .A2(new_n245_), .A3(new_n247_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n229_), .A2(new_n231_), .A3(new_n235_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(KEYINPUT95), .A3(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n225_), .B1(new_n249_), .B2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G211gat), .B(G218gat), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(G197gat), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n256_), .A2(G204gat), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n257_), .A2(KEYINPUT91), .ZN(new_n258_));
  AND2_X1   g057(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n259_));
  NOR2_X1   g058(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(G204gat), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n257_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n258_), .B1(new_n263_), .B2(KEYINPUT91), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT21), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n255_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  OR2_X1    g065(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(G204gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n271_), .B(KEYINPUT21), .C1(new_n256_), .C2(new_n270_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n254_), .A2(KEYINPUT92), .ZN(new_n273_));
  OR2_X1    g072(.A1(G211gat), .A2(G218gat), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT92), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G211gat), .A2(G218gat), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n273_), .A2(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n270_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT91), .B1(new_n279_), .B2(new_n257_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n258_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n278_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  AOI22_X1  g081(.A1(new_n266_), .A2(new_n272_), .B1(KEYINPUT21), .B2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT96), .B1(new_n253_), .B2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n220_), .A2(new_n221_), .A3(new_n224_), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n250_), .A2(KEYINPUT95), .A3(new_n251_), .ZN(new_n286_));
  AOI21_X1  g085(.A(KEYINPUT95), .B1(new_n250_), .B2(new_n251_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n285_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT96), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n280_), .A2(new_n281_), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n272_), .B(new_n254_), .C1(new_n290_), .C2(KEYINPUT21), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n282_), .A2(KEYINPUT21), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n288_), .A2(new_n289_), .A3(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n284_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(KEYINPUT81), .A2(G169gat), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n296_), .A2(KEYINPUT22), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n223_), .B1(new_n296_), .B2(KEYINPUT22), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n221_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n300_), .B1(new_n236_), .B2(new_n218_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(KEYINPUT78), .A2(G183gat), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n302_), .A2(KEYINPUT25), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(KEYINPUT25), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n303_), .A2(new_n243_), .A3(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n238_), .A2(KEYINPUT24), .A3(new_n221_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n237_), .A2(new_n239_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n217_), .A2(new_n305_), .A3(new_n306_), .A4(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n301_), .A2(KEYINPUT83), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT83), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n299_), .B1(new_n251_), .B2(new_n219_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n308_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n310_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n309_), .A2(new_n283_), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT20), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G226gat), .A2(G233gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT19), .ZN(new_n317_));
  NOR3_X1   g116(.A1(new_n295_), .A2(new_n315_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n317_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n250_), .A2(new_n251_), .ZN(new_n320_));
  AND4_X1   g119(.A1(new_n291_), .A2(new_n292_), .A3(new_n285_), .A4(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n309_), .A2(new_n313_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n321_), .B1(new_n322_), .B2(new_n293_), .ZN(new_n323_));
  XOR2_X1   g122(.A(KEYINPUT99), .B(KEYINPUT20), .Z(new_n324_));
  AOI21_X1  g123(.A(new_n319_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n206_), .B1(new_n318_), .B2(new_n325_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n284_), .A2(new_n294_), .A3(KEYINPUT20), .A4(new_n314_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n317_), .ZN(new_n328_));
  AOI21_X1  g127(.A(KEYINPUT83), .B1(new_n301_), .B2(new_n308_), .ZN(new_n329_));
  NOR3_X1   g128(.A1(new_n311_), .A2(new_n312_), .A3(new_n310_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n293_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n253_), .A2(new_n283_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n331_), .A2(KEYINPUT20), .A3(new_n319_), .A4(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n328_), .A2(new_n205_), .A3(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n326_), .A2(KEYINPUT27), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT101), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT27), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n283_), .A2(new_n285_), .A3(new_n320_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n331_), .A2(new_n324_), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(new_n317_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n341_), .B1(new_n317_), .B2(new_n327_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n338_), .B1(new_n342_), .B2(new_n206_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n343_), .A2(KEYINPUT101), .A3(new_n334_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n337_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n328_), .A2(new_n333_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(new_n206_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n334_), .ZN(new_n348_));
  XOR2_X1   g147(.A(KEYINPUT102), .B(KEYINPUT27), .Z(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n345_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT100), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT88), .ZN(new_n353_));
  INV_X1    g152(.A(G141gat), .ZN(new_n354_));
  INV_X1    g153(.A(G148gat), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n353_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT2), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G141gat), .A2(G148gat), .ZN(new_n358_));
  AOI22_X1  g157(.A1(new_n356_), .A2(KEYINPUT3), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n359_), .B(new_n360_), .C1(KEYINPUT3), .C2(new_n356_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G155gat), .A2(G162gat), .ZN(new_n362_));
  INV_X1    g161(.A(G155gat), .ZN(new_n363_));
  INV_X1    g162(.A(G162gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n361_), .A2(new_n362_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n354_), .A2(new_n355_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n362_), .A2(KEYINPUT1), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT87), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n362_), .A2(KEYINPUT87), .A3(KEYINPUT1), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(new_n371_), .A3(new_n365_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n362_), .A2(KEYINPUT1), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n367_), .B(new_n358_), .C1(new_n372_), .C2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n366_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT86), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G127gat), .B(G134gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G113gat), .B(G120gat), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n376_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n377_), .B(new_n378_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n379_), .B1(new_n380_), .B2(new_n376_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n375_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G225gat), .A2(G233gat), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n366_), .A2(new_n380_), .A3(new_n374_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n382_), .A2(new_n384_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT4), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT4), .B1(new_n375_), .B2(new_n381_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n383_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n386_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G1gat), .B(G29gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(G85gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT0), .ZN(new_n396_));
  INV_X1    g195(.A(G57gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n352_), .B1(new_n393_), .B2(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n389_), .B1(new_n387_), .B2(KEYINPUT4), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n385_), .B(new_n398_), .C1(new_n400_), .C2(new_n383_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n385_), .B1(new_n400_), .B2(new_n383_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n398_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(KEYINPUT100), .A3(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n399_), .A2(new_n401_), .A3(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G15gat), .B(G43gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT84), .B(KEYINPUT85), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n322_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n381_), .B(KEYINPUT30), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n411_), .ZN(new_n413_));
  XOR2_X1   g212(.A(G71gat), .B(G99gat), .Z(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT31), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G227gat), .A2(G233gat), .ZN(new_n416_));
  XOR2_X1   g215(.A(new_n415_), .B(new_n416_), .Z(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n412_), .A2(new_n413_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n418_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n409_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n421_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n423_), .A2(new_n408_), .A3(new_n419_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT29), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n366_), .A2(new_n426_), .A3(new_n374_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT93), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n283_), .B1(KEYINPUT29), .B2(new_n375_), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n429_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G22gat), .B(G50gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G228gat), .A2(G233gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n436_));
  XOR2_X1   g235(.A(new_n435_), .B(new_n436_), .Z(new_n437_));
  XOR2_X1   g236(.A(G78gat), .B(G106gat), .Z(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n432_), .A2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n430_), .A2(new_n431_), .A3(new_n439_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n425_), .A2(new_n443_), .ZN(new_n444_));
  NOR3_X1   g243(.A1(new_n351_), .A2(new_n405_), .A3(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n405_), .A2(new_n443_), .ZN(new_n446_));
  AOI21_X1  g245(.A(KEYINPUT101), .B1(new_n343_), .B2(new_n334_), .ZN(new_n447_));
  AND4_X1   g246(.A1(KEYINPUT101), .A2(new_n326_), .A3(KEYINPUT27), .A4(new_n334_), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n350_), .B(new_n446_), .C1(new_n447_), .C2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT103), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n342_), .A2(new_n451_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n405_), .B(new_n452_), .C1(new_n346_), .C2(new_n451_), .ZN(new_n453_));
  OR2_X1    g252(.A1(new_n387_), .A2(KEYINPUT97), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n387_), .A2(KEYINPUT97), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(new_n392_), .A3(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n403_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT98), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n391_), .A2(new_n383_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT98), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n456_), .A2(new_n460_), .A3(new_n403_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n458_), .A2(new_n459_), .A3(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n401_), .B(KEYINPUT33), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n462_), .A2(new_n334_), .A3(new_n463_), .A4(new_n347_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n453_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(new_n443_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT103), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n345_), .A2(new_n467_), .A3(new_n350_), .A4(new_n446_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n450_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n425_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n445_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G176gat), .B(G204gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G120gat), .B(G148gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n474_), .B(new_n475_), .Z(new_n476_));
  NAND2_X1  g275(.A1(G85gat), .A2(G92gat), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(G85gat), .A2(G92gat), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(G99gat), .A2(G106gat), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT7), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n480_), .B1(new_n483_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT8), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n481_), .B(KEYINPUT7), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT65), .ZN(new_n491_));
  INV_X1    g290(.A(new_n486_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n491_), .B1(new_n492_), .B2(new_n484_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n485_), .A2(KEYINPUT65), .A3(new_n486_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n490_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  NOR3_X1   g294(.A1(new_n478_), .A2(new_n479_), .A3(KEYINPUT8), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n489_), .A2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n499_));
  OAI22_X1  g298(.A1(new_n499_), .A2(KEYINPUT64), .B1(G85gat), .B2(G92gat), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT9), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n477_), .A2(KEYINPUT64), .A3(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n477_), .A2(new_n501_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n500_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n494_), .A2(new_n493_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(KEYINPUT10), .B(G99gat), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n506_), .A2(G106gat), .ZN(new_n507_));
  OR3_X1    g306(.A1(new_n504_), .A2(new_n505_), .A3(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n498_), .A2(new_n508_), .A3(KEYINPUT66), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT66), .ZN(new_n510_));
  AOI22_X1  g309(.A1(KEYINPUT8), .A2(new_n488_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n511_));
  NOR3_X1   g310(.A1(new_n504_), .A2(new_n505_), .A3(new_n507_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n510_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(G71gat), .B(G78gat), .Z(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G57gat), .B(G64gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT11), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n516_), .A2(KEYINPUT11), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n514_), .A2(KEYINPUT11), .A3(new_n516_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n509_), .A2(new_n513_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT12), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n521_), .ZN(new_n525_));
  AOI211_X1 g324(.A(new_n523_), .B(new_n525_), .C1(new_n498_), .C2(new_n508_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT67), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n521_), .B1(new_n509_), .B2(new_n513_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G230gat), .A2(G233gat), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n529_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n509_), .A2(new_n513_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n525_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n535_), .A2(KEYINPUT67), .A3(new_n531_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n528_), .B1(new_n533_), .B2(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n531_), .B1(new_n535_), .B2(new_n522_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n476_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT69), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n526_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n541_));
  AOI21_X1  g340(.A(KEYINPUT67), .B1(new_n535_), .B2(new_n531_), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n530_), .A2(new_n529_), .A3(new_n532_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n541_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n538_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n476_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n544_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n539_), .A2(new_n540_), .A3(new_n547_), .ZN(new_n548_));
  OAI211_X1 g347(.A(KEYINPUT69), .B(new_n476_), .C1(new_n537_), .C2(new_n538_), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n548_), .A2(KEYINPUT13), .A3(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT13), .B1(new_n548_), .B2(new_n549_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT70), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT70), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n554_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G113gat), .B(G141gat), .ZN(new_n557_));
  INV_X1    g356(.A(G169gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(new_n256_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G15gat), .B(G22gat), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G1gat), .A2(G8gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT14), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G1gat), .B(G8gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT15), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G29gat), .B(G36gat), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n569_), .A2(G43gat), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(G43gat), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n570_), .A2(G50gat), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(G50gat), .B1(new_n570_), .B2(new_n571_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n568_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n574_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n576_), .A2(new_n572_), .A3(KEYINPUT15), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n567_), .B1(new_n575_), .B2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G229gat), .A2(G233gat), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n567_), .A2(new_n572_), .A3(new_n576_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n578_), .A2(new_n580_), .A3(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n576_), .A2(new_n572_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(new_n566_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n579_), .B1(new_n585_), .B2(new_n581_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n560_), .B1(new_n583_), .B2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n575_), .A2(new_n577_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(new_n566_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n589_), .A2(new_n579_), .A3(new_n581_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n586_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n560_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n590_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n587_), .A2(new_n593_), .A3(KEYINPUT76), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT76), .ZN(new_n595_));
  OAI211_X1 g394(.A(new_n595_), .B(new_n560_), .C1(new_n583_), .C2(new_n586_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT77), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n471_), .A2(new_n556_), .A3(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n584_), .B1(new_n509_), .B2(new_n513_), .ZN(new_n601_));
  AOI22_X1  g400(.A1(new_n575_), .A2(new_n577_), .B1(new_n498_), .B2(new_n508_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G232gat), .A2(G233gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT34), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT35), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n604_), .A2(KEYINPUT35), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NOR4_X1   g408(.A1(new_n601_), .A2(new_n602_), .A3(KEYINPUT72), .A4(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n606_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT72), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n601_), .A2(new_n602_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(new_n608_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n610_), .B1(new_n613_), .B2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G190gat), .B(G218gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(G134gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(new_n364_), .ZN(new_n619_));
  XOR2_X1   g418(.A(KEYINPUT71), .B(KEYINPUT36), .Z(new_n620_));
  NAND3_X1  g419(.A1(new_n616_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT37), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n619_), .B(KEYINPUT36), .ZN(new_n623_));
  AOI22_X1  g422(.A1(new_n611_), .A2(new_n612_), .B1(new_n614_), .B2(new_n608_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n623_), .B1(new_n624_), .B2(new_n610_), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n621_), .A2(new_n622_), .A3(new_n625_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n623_), .B(KEYINPUT73), .Z(new_n627_));
  OAI21_X1  g426(.A(new_n627_), .B1(new_n624_), .B2(new_n610_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(KEYINPUT74), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT74), .ZN(new_n630_));
  OAI211_X1 g429(.A(new_n630_), .B(new_n627_), .C1(new_n624_), .C2(new_n610_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n629_), .A2(new_n621_), .A3(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n626_), .B1(KEYINPUT37), .B2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(G127gat), .B(G155gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT16), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(G183gat), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(G211gat), .Z(new_n637_));
  INV_X1    g436(.A(KEYINPUT17), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n566_), .B(new_n521_), .ZN(new_n640_));
  AND2_X1   g439(.A1(G231gat), .A2(G233gat), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n640_), .B(new_n641_), .Z(new_n642_));
  NAND2_X1  g441(.A1(new_n639_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT75), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n637_), .A2(new_n638_), .ZN(new_n646_));
  OR3_X1    g445(.A1(new_n642_), .A2(new_n646_), .A3(new_n639_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n633_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n600_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n405_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n650_), .A2(G1gat), .A3(new_n651_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT38), .Z(new_n653_));
  NAND2_X1  g452(.A1(new_n621_), .A2(new_n625_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n471_), .A2(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n556_), .A2(new_n597_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n648_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n656_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G1gat), .B1(new_n659_), .B2(new_n651_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n653_), .A2(new_n660_), .ZN(G1324gat));
  INV_X1    g460(.A(new_n351_), .ZN(new_n662_));
  OR3_X1    g461(.A1(new_n650_), .A2(G8gat), .A3(new_n662_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n656_), .A2(new_n657_), .A3(new_n658_), .A4(new_n351_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT39), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n664_), .A2(new_n665_), .A3(G8gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n664_), .B2(G8gat), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n663_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(KEYINPUT104), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT104), .ZN(new_n670_));
  OAI211_X1 g469(.A(new_n663_), .B(new_n670_), .C1(new_n666_), .C2(new_n667_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT40), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n669_), .A2(KEYINPUT40), .A3(new_n671_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1325gat));
  OAI21_X1  g475(.A(G15gat), .B1(new_n659_), .B2(new_n470_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT41), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n650_), .A2(G15gat), .A3(new_n470_), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1326gat));
  OAI21_X1  g479(.A(G22gat), .B1(new_n659_), .B2(new_n443_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT42), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n443_), .A2(G22gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n682_), .B1(new_n650_), .B2(new_n683_), .ZN(G1327gat));
  NAND2_X1  g483(.A1(new_n469_), .A2(new_n470_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n445_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n632_), .A2(KEYINPUT37), .ZN(new_n688_));
  INV_X1    g487(.A(new_n626_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n690_), .A2(KEYINPUT43), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n687_), .A2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n690_), .B(KEYINPUT105), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT43), .B1(new_n471_), .B2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n556_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n594_), .A2(new_n596_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n696_), .A2(new_n648_), .A3(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n695_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n695_), .A2(KEYINPUT44), .A3(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G29gat), .B1(new_n704_), .B2(new_n651_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n599_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n658_), .A2(new_n654_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n687_), .A2(new_n696_), .A3(new_n706_), .A4(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT106), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n600_), .A2(KEYINPUT106), .A3(new_n707_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  OR3_X1    g511(.A1(new_n712_), .A2(G29gat), .A3(new_n651_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n705_), .A2(new_n713_), .ZN(G1328gat));
  INV_X1    g513(.A(KEYINPUT46), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT107), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n715_), .A2(KEYINPUT107), .ZN(new_n717_));
  INV_X1    g516(.A(G36gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT44), .B1(new_n695_), .B2(new_n699_), .ZN(new_n719_));
  AOI211_X1 g518(.A(new_n701_), .B(new_n698_), .C1(new_n692_), .C2(new_n694_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n718_), .B1(new_n721_), .B2(new_n351_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n662_), .A2(G36gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n710_), .A2(new_n711_), .A3(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT45), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n710_), .A2(new_n711_), .A3(KEYINPUT45), .A4(new_n723_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n716_), .B(new_n717_), .C1(new_n722_), .C2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n728_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n702_), .A2(new_n351_), .A3(new_n703_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(G36gat), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n730_), .A2(new_n732_), .A3(KEYINPUT107), .A4(new_n715_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n729_), .A2(new_n733_), .ZN(G1329gat));
  NAND3_X1  g533(.A1(new_n710_), .A2(new_n711_), .A3(new_n425_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n736_));
  INV_X1    g535(.A(G43gat), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n735_), .A2(new_n736_), .A3(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n736_), .B1(new_n735_), .B2(new_n737_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n425_), .A2(G43gat), .ZN(new_n740_));
  OAI22_X1  g539(.A1(new_n738_), .A2(new_n739_), .B1(new_n704_), .B2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT47), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT47), .ZN(new_n743_));
  OAI221_X1 g542(.A(new_n743_), .B1(new_n704_), .B2(new_n740_), .C1(new_n738_), .C2(new_n739_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1330gat));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n746_), .B1(new_n704_), .B2(new_n443_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n443_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n721_), .A2(KEYINPUT109), .A3(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n747_), .A2(G50gat), .A3(new_n749_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n443_), .A2(G50gat), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT110), .Z(new_n752_));
  OAI21_X1  g551(.A(new_n750_), .B1(new_n712_), .B2(new_n752_), .ZN(G1331gat));
  NAND2_X1  g552(.A1(new_n658_), .A2(new_n599_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n656_), .A2(new_n556_), .A3(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT112), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT112), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n656_), .A2(new_n758_), .A3(new_n556_), .A4(new_n755_), .ZN(new_n759_));
  AND4_X1   g558(.A1(G57gat), .A2(new_n757_), .A3(new_n405_), .A4(new_n759_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n471_), .A2(new_n696_), .A3(new_n697_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(new_n649_), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT111), .Z(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n405_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n760_), .B1(new_n764_), .B2(new_n397_), .ZN(G1332gat));
  NAND3_X1  g564(.A1(new_n757_), .A2(new_n351_), .A3(new_n759_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(G64gat), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n767_), .A2(KEYINPUT48), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(KEYINPUT48), .ZN(new_n769_));
  INV_X1    g568(.A(new_n763_), .ZN(new_n770_));
  OR2_X1    g569(.A1(new_n662_), .A2(G64gat), .ZN(new_n771_));
  OAI22_X1  g570(.A1(new_n768_), .A2(new_n769_), .B1(new_n770_), .B2(new_n771_), .ZN(G1333gat));
  NOR2_X1   g571(.A1(new_n470_), .A2(G71gat), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n763_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n757_), .A2(new_n425_), .A3(new_n759_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT49), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n775_), .A2(new_n776_), .A3(G71gat), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n775_), .B2(G71gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n774_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT113), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n774_), .B(new_n781_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(G1334gat));
  OR2_X1    g582(.A1(new_n443_), .A2(G78gat), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n757_), .A2(new_n748_), .A3(new_n759_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT50), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n785_), .A2(new_n786_), .A3(G78gat), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n785_), .B2(G78gat), .ZN(new_n788_));
  OAI22_X1  g587(.A1(new_n770_), .A2(new_n784_), .B1(new_n787_), .B2(new_n788_), .ZN(G1335gat));
  AND2_X1   g588(.A1(new_n761_), .A2(new_n707_), .ZN(new_n790_));
  AOI21_X1  g589(.A(G85gat), .B1(new_n790_), .B2(new_n405_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n556_), .A2(new_n648_), .A3(new_n597_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n792_), .B(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n695_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT115), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n405_), .A2(G85gat), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT116), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n791_), .B1(new_n796_), .B2(new_n798_), .ZN(G1336gat));
  AOI21_X1  g598(.A(G92gat), .B1(new_n790_), .B2(new_n351_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n796_), .A2(new_n351_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n801_), .B2(G92gat), .ZN(G1337gat));
  NAND3_X1  g601(.A1(new_n794_), .A2(new_n425_), .A3(new_n695_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n470_), .A2(new_n506_), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n803_), .A2(G99gat), .B1(new_n790_), .B2(new_n804_), .ZN(new_n805_));
  XOR2_X1   g604(.A(new_n805_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g605(.A(G106gat), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n790_), .A2(new_n807_), .A3(new_n748_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n794_), .A2(new_n748_), .A3(new_n695_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n809_), .A2(new_n810_), .A3(G106gat), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n810_), .B1(new_n809_), .B2(G106gat), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n808_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n548_), .A2(new_n549_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n585_), .A2(new_n581_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n578_), .A2(new_n582_), .ZN(new_n818_));
  MUX2_X1   g617(.A(new_n817_), .B(new_n818_), .S(new_n580_), .Z(new_n819_));
  OAI21_X1  g618(.A(new_n593_), .B1(new_n819_), .B2(new_n592_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n816_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n544_), .A2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n532_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n824_));
  OAI211_X1 g623(.A(KEYINPUT55), .B(new_n541_), .C1(new_n542_), .C2(new_n543_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n823_), .A2(new_n824_), .A3(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n826_), .A2(KEYINPUT118), .A3(new_n476_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT119), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT56), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n826_), .A2(new_n476_), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT118), .B1(new_n830_), .B2(KEYINPUT119), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n537_), .A2(new_n538_), .A3(new_n476_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(new_n597_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n697_), .A2(new_n547_), .A3(KEYINPUT117), .ZN(new_n837_));
  AOI22_X1  g636(.A1(new_n832_), .A2(new_n833_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n821_), .B1(new_n831_), .B2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n815_), .B1(new_n839_), .B2(new_n655_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n832_), .A2(new_n833_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n836_), .A2(new_n837_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(KEYINPUT56), .B1(new_n827_), .B2(new_n828_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  OAI211_X1 g644(.A(KEYINPUT57), .B(new_n654_), .C1(new_n845_), .C2(new_n821_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT120), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n830_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n832_), .A2(new_n847_), .A3(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n835_), .A2(new_n820_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n826_), .A2(new_n848_), .A3(new_n830_), .A4(new_n476_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n850_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT58), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n850_), .A2(KEYINPUT58), .A3(new_n851_), .A4(new_n852_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(new_n633_), .A3(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n840_), .A2(new_n846_), .A3(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n648_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(KEYINPUT121), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n861_));
  INV_X1    g660(.A(new_n551_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n548_), .A2(KEYINPUT13), .A3(new_n549_), .ZN(new_n863_));
  AOI22_X1  g662(.A1(new_n862_), .A2(new_n863_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n861_), .B1(new_n864_), .B2(new_n755_), .ZN(new_n865_));
  NOR4_X1   g664(.A1(new_n552_), .A2(new_n633_), .A3(new_n754_), .A4(KEYINPUT54), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n858_), .A2(new_n869_), .A3(new_n648_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n860_), .A2(new_n868_), .A3(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n351_), .A2(new_n651_), .A3(new_n444_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n871_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT122), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n859_), .A2(new_n868_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n873_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(KEYINPUT59), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n871_), .A2(KEYINPUT122), .A3(new_n872_), .A4(new_n873_), .ZN(new_n880_));
  INV_X1    g679(.A(G113gat), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n599_), .A2(new_n881_), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n876_), .A2(new_n879_), .A3(new_n880_), .A4(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n881_), .B1(new_n878_), .B2(new_n597_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1340gat));
  NAND3_X1  g684(.A1(new_n876_), .A2(new_n879_), .A3(new_n880_), .ZN(new_n886_));
  OAI21_X1  g685(.A(G120gat), .B1(new_n886_), .B2(new_n696_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n878_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT60), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n889_), .B1(new_n696_), .B2(G120gat), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n888_), .B(new_n890_), .C1(new_n889_), .C2(G120gat), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n887_), .A2(new_n893_), .ZN(G1341gat));
  INV_X1    g693(.A(G127gat), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n648_), .A2(new_n895_), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n876_), .A2(new_n879_), .A3(new_n880_), .A4(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n895_), .B1(new_n878_), .B2(new_n648_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1342gat));
  INV_X1    g698(.A(G134gat), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n690_), .A2(new_n900_), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n876_), .A2(new_n879_), .A3(new_n880_), .A4(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n900_), .B1(new_n878_), .B2(new_n654_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1343gat));
  AOI21_X1  g703(.A(new_n867_), .B1(new_n858_), .B2(new_n648_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n351_), .A2(new_n651_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n425_), .A2(new_n443_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n905_), .A2(new_n907_), .A3(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n697_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g711(.A1(new_n910_), .A2(new_n556_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g713(.A1(new_n877_), .A2(new_n658_), .A3(new_n906_), .A4(new_n908_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(KEYINPUT124), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n910_), .A2(new_n917_), .A3(new_n658_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT61), .ZN(new_n919_));
  AND3_X1   g718(.A1(new_n916_), .A2(new_n918_), .A3(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n919_), .B1(new_n916_), .B2(new_n918_), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n920_), .A2(new_n921_), .A3(new_n363_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n915_), .A2(KEYINPUT124), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n917_), .B1(new_n910_), .B2(new_n658_), .ZN(new_n924_));
  OAI21_X1  g723(.A(KEYINPUT61), .B1(new_n923_), .B2(new_n924_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n916_), .A2(new_n918_), .A3(new_n919_), .ZN(new_n926_));
  AOI21_X1  g725(.A(G155gat), .B1(new_n925_), .B2(new_n926_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n922_), .A2(new_n927_), .ZN(G1346gat));
  AOI21_X1  g727(.A(G162gat), .B1(new_n910_), .B2(new_n655_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n693_), .A2(new_n364_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n929_), .B1(new_n910_), .B2(new_n930_), .ZN(G1347gat));
  NAND2_X1  g730(.A1(new_n351_), .A2(new_n651_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n932_), .A2(new_n444_), .ZN(new_n933_));
  AND2_X1   g732(.A1(new_n871_), .A2(new_n933_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n558_), .B1(new_n934_), .B2(new_n697_), .ZN(new_n935_));
  OR2_X1    g734(.A1(new_n935_), .A2(KEYINPUT62), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n934_), .A2(new_n222_), .A3(new_n697_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n935_), .A2(KEYINPUT62), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n936_), .A2(new_n937_), .A3(new_n938_), .ZN(G1348gat));
  NAND2_X1  g738(.A1(new_n934_), .A2(new_n556_), .ZN(new_n940_));
  AND3_X1   g739(.A1(new_n940_), .A2(KEYINPUT125), .A3(new_n223_), .ZN(new_n941_));
  AOI21_X1  g740(.A(KEYINPUT125), .B1(new_n940_), .B2(new_n223_), .ZN(new_n942_));
  NOR3_X1   g741(.A1(new_n905_), .A2(new_n444_), .A3(new_n932_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n943_), .A2(G176gat), .A3(new_n556_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(KEYINPUT126), .ZN(new_n945_));
  NOR3_X1   g744(.A1(new_n941_), .A2(new_n942_), .A3(new_n945_), .ZN(G1349gat));
  AOI21_X1  g745(.A(G183gat), .B1(new_n943_), .B2(new_n658_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n648_), .A2(new_n244_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n947_), .B1(new_n934_), .B2(new_n948_), .ZN(G1350gat));
  NAND2_X1  g748(.A1(new_n934_), .A2(new_n633_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n950_), .A2(G190gat), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n934_), .A2(new_n655_), .A3(new_n243_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n951_), .A2(new_n952_), .ZN(G1351gat));
  NOR3_X1   g752(.A1(new_n905_), .A2(new_n909_), .A3(new_n932_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n954_), .A2(new_n697_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n955_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g755(.A1(new_n954_), .A2(new_n556_), .ZN(new_n957_));
  XNOR2_X1  g756(.A(new_n957_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g757(.A1(new_n954_), .A2(new_n658_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n960_));
  AND2_X1   g759(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n961_));
  NOR3_X1   g760(.A1(new_n959_), .A2(new_n960_), .A3(new_n961_), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n962_), .B1(new_n959_), .B2(new_n960_), .ZN(G1354gat));
  NAND2_X1  g762(.A1(new_n954_), .A2(new_n655_), .ZN(new_n964_));
  XNOR2_X1  g763(.A(KEYINPUT127), .B(G218gat), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n690_), .A2(new_n965_), .ZN(new_n966_));
  AOI22_X1  g765(.A1(new_n964_), .A2(new_n965_), .B1(new_n954_), .B2(new_n966_), .ZN(G1355gat));
endmodule


