//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n900_, new_n902_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n935_, new_n936_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G226gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  XOR2_X1   g008(.A(G197gat), .B(G204gat), .Z(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT21), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G211gat), .B(G218gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G197gat), .B(G204gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT21), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n211_), .A2(new_n212_), .A3(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT87), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n212_), .A2(KEYINPUT88), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n212_), .A2(KEYINPUT88), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n218_), .A2(KEYINPUT21), .A3(new_n219_), .A4(new_n210_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n217_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  OR2_X1    g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n223_), .A2(KEYINPUT24), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(KEYINPUT24), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n224_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT26), .B(G190gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT25), .B(G183gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n228_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n233_), .A2(KEYINPUT83), .A3(KEYINPUT23), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT82), .B(KEYINPUT23), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n234_), .B1(new_n235_), .B2(new_n233_), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT83), .B1(new_n233_), .B2(KEYINPUT23), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n235_), .A2(new_n233_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n239_), .B1(KEYINPUT23), .B2(new_n233_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n240_), .B1(G183gat), .B2(G190gat), .ZN(new_n241_));
  NOR2_X1   g040(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(G169gat), .ZN(new_n243_));
  AOI22_X1  g042(.A1(new_n232_), .A2(new_n238_), .B1(new_n241_), .B2(new_n243_), .ZN(new_n244_));
  OR3_X1    g043(.A1(new_n222_), .A2(KEYINPUT95), .A3(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT95), .B1(new_n222_), .B2(new_n244_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n238_), .B1(G183gat), .B2(G190gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(new_n243_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT81), .ZN(new_n250_));
  INV_X1    g049(.A(G183gat), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n250_), .B1(new_n251_), .B2(KEYINPUT25), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n229_), .B(new_n252_), .C1(new_n230_), .C2(new_n250_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n228_), .A2(new_n240_), .A3(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n249_), .A2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(KEYINPUT20), .B1(new_n255_), .B2(new_n221_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n209_), .B1(new_n247_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n255_), .A2(new_n221_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n259_), .A2(KEYINPUT20), .A3(new_n209_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n222_), .A2(new_n244_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n206_), .B1(new_n258_), .B2(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n256_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n264_));
  OAI221_X1 g063(.A(new_n205_), .B1(new_n261_), .B2(new_n260_), .C1(new_n264_), .C2(new_n209_), .ZN(new_n265_));
  AOI21_X1  g064(.A(KEYINPUT27), .B1(new_n263_), .B2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n221_), .B(KEYINPUT90), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(new_n244_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT20), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT97), .ZN(new_n270_));
  AOI22_X1  g069(.A1(new_n269_), .A2(new_n270_), .B1(new_n221_), .B2(new_n255_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n268_), .A2(KEYINPUT97), .A3(KEYINPUT20), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n209_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n264_), .A2(new_n209_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n206_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n265_), .A2(KEYINPUT27), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n266_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(G141gat), .A2(G148gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT3), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G141gat), .A2(G148gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT2), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT86), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285_));
  NOR2_X1   g084(.A1(G155gat), .A2(G162gat), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n284_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n286_), .B1(KEYINPUT1), .B2(new_n285_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n289_), .B1(KEYINPUT1), .B2(new_n285_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n278_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n290_), .A2(new_n291_), .A3(new_n280_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n288_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT29), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G228gat), .A2(G233gat), .ZN(new_n295_));
  AND3_X1   g094(.A1(new_n294_), .A2(new_n295_), .A3(new_n221_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT89), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT90), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n221_), .B(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n293_), .A2(KEYINPUT89), .A3(KEYINPUT29), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n298_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n295_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n296_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G78gat), .B(G106gat), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT91), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(KEYINPUT91), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n304_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G22gat), .B(G50gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT28), .B1(new_n293_), .B2(KEYINPUT29), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NOR3_X1   g113(.A1(new_n293_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n312_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n315_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n317_), .A2(new_n313_), .A3(new_n311_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n319_), .B1(new_n304_), .B2(new_n308_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n310_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT93), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n316_), .A2(new_n318_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n306_), .A2(KEYINPUT92), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n323_), .B1(new_n304_), .B2(new_n325_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n304_), .A2(new_n325_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n322_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n304_), .A2(new_n325_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n304_), .A2(new_n325_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n329_), .A2(KEYINPUT93), .A3(new_n323_), .A4(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n321_), .B1(new_n328_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G225gat), .A2(G233gat), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G127gat), .B(G134gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G113gat), .B(G120gat), .ZN(new_n336_));
  OR2_X1    g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT84), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n335_), .A2(new_n336_), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n339_), .B(new_n340_), .Z(new_n341_));
  NAND2_X1  g140(.A1(new_n293_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n337_), .A2(new_n340_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n288_), .A2(new_n292_), .A3(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n342_), .A2(KEYINPUT4), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT4), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n293_), .A2(new_n346_), .A3(new_n341_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT96), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n347_), .A2(new_n348_), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n334_), .B(new_n345_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n342_), .A2(new_n344_), .A3(new_n333_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G1gat), .B(G29gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(G85gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT0), .B(G57gat), .ZN(new_n355_));
  XOR2_X1   g154(.A(new_n354_), .B(new_n355_), .Z(new_n356_));
  NAND3_X1  g155(.A1(new_n351_), .A2(new_n352_), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT98), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n351_), .A2(new_n352_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n356_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT98), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n351_), .A2(new_n362_), .A3(new_n352_), .A4(new_n356_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n358_), .A2(new_n361_), .A3(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G71gat), .B(G99gat), .ZN(new_n365_));
  INV_X1    g164(.A(G43gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n255_), .B(new_n367_), .Z(new_n368_));
  XOR2_X1   g167(.A(new_n341_), .B(KEYINPUT85), .Z(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G227gat), .A2(G233gat), .ZN(new_n371_));
  INV_X1    g170(.A(G15gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT30), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT31), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n370_), .B(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n364_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n277_), .A2(new_n332_), .A3(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n332_), .A2(new_n364_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n263_), .A2(new_n265_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT33), .ZN(new_n381_));
  OR2_X1    g180(.A1(new_n357_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n357_), .A2(new_n381_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n333_), .B(new_n345_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n342_), .A2(new_n344_), .A3(new_n334_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n384_), .A2(new_n360_), .A3(new_n385_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n380_), .A2(new_n382_), .A3(new_n383_), .A4(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n258_), .A2(new_n262_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n269_), .A2(new_n270_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n391_), .A2(new_n259_), .A3(new_n272_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n209_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n274_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n390_), .B1(new_n394_), .B2(new_n389_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n364_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n387_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n379_), .A2(new_n277_), .B1(new_n397_), .B2(new_n332_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n376_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n378_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT65), .ZN(new_n402_));
  OAI22_X1  g201(.A1(new_n402_), .A2(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT9), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n404_), .A2(KEYINPUT65), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(G85gat), .ZN(new_n407_));
  OR2_X1    g206(.A1(KEYINPUT66), .A2(G92gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(KEYINPUT66), .A2(G92gat), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n407_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n401_), .B1(new_n406_), .B2(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(KEYINPUT10), .B(G99gat), .Z(new_n412_));
  INV_X1    g211(.A(G106gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G99gat), .A2(G106gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT6), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT6), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(G99gat), .A3(G106gat), .ZN(new_n417_));
  AOI22_X1  g216(.A1(new_n412_), .A2(new_n413_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n411_), .A2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G85gat), .B(G92gat), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NOR3_X1   g221(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n415_), .A2(new_n417_), .ZN(new_n425_));
  AOI211_X1 g224(.A(KEYINPUT8), .B(new_n420_), .C1(new_n424_), .C2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT8), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT7), .ZN(new_n428_));
  INV_X1    g227(.A(G99gat), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(new_n429_), .A3(new_n413_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n416_), .B1(G99gat), .B2(G106gat), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n414_), .A2(KEYINPUT6), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n421_), .B(new_n430_), .C1(new_n431_), .C2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n420_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n427_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n419_), .B1(new_n426_), .B2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G57gat), .B(G64gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G71gat), .B(G78gat), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(KEYINPUT11), .ZN(new_n439_));
  INV_X1    g238(.A(new_n438_), .ZN(new_n440_));
  INV_X1    g239(.A(G64gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(G57gat), .ZN(new_n442_));
  INV_X1    g241(.A(G57gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(G64gat), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n444_), .A3(KEYINPUT11), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n440_), .A2(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n437_), .A2(KEYINPUT11), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n439_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n436_), .A2(new_n449_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n419_), .B(new_n448_), .C1(new_n426_), .C2(new_n435_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n450_), .A2(KEYINPUT12), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT12), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n436_), .A2(new_n453_), .A3(new_n449_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G230gat), .A2(G233gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT64), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n455_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n450_), .A2(new_n451_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT67), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n460_), .A2(new_n461_), .A3(new_n457_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n433_), .A2(new_n434_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT8), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n433_), .A2(new_n427_), .A3(new_n434_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n448_), .B1(new_n466_), .B2(new_n419_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n451_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n457_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT67), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G120gat), .B(G148gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT5), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G176gat), .B(G204gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n459_), .A2(new_n462_), .A3(new_n470_), .A4(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT68), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n461_), .B1(new_n460_), .B2(new_n457_), .ZN(new_n477_));
  AOI211_X1 g276(.A(KEYINPUT67), .B(new_n458_), .C1(new_n450_), .C2(new_n451_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT68), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n479_), .A2(new_n480_), .A3(new_n459_), .A4(new_n474_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n476_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n474_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n470_), .A2(new_n462_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n457_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n483_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n482_), .A2(KEYINPUT13), .A3(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(KEYINPUT13), .B1(new_n482_), .B2(new_n486_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT69), .ZN(new_n491_));
  INV_X1    g290(.A(new_n489_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(new_n487_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT69), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n491_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G229gat), .A2(G233gat), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT73), .B(G8gat), .ZN(new_n500_));
  INV_X1    g299(.A(G1gat), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT14), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G15gat), .B(G22gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G1gat), .B(G8gat), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n508_));
  INV_X1    g307(.A(G8gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT73), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT73), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(G8gat), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n501_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT14), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n505_), .B(new_n503_), .C1(new_n513_), .C2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n507_), .A2(new_n508_), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n508_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n515_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n505_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n517_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G43gat), .B(G50gat), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G29gat), .B(G36gat), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n523_), .A2(KEYINPUT70), .ZN(new_n524_));
  INV_X1    g323(.A(G36gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(G29gat), .ZN(new_n526_));
  INV_X1    g325(.A(G29gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(G36gat), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n526_), .A2(new_n528_), .A3(KEYINPUT70), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n522_), .B1(new_n524_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n526_), .A2(new_n528_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT70), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n523_), .A2(KEYINPUT70), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(new_n534_), .A3(new_n521_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n530_), .A2(new_n535_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n516_), .A2(new_n520_), .A3(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n536_), .B1(new_n516_), .B2(new_n520_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n499_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G113gat), .B(G141gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G169gat), .B(G197gat), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n540_), .B(new_n541_), .Z(new_n542_));
  NOR2_X1   g341(.A1(new_n542_), .A2(KEYINPUT80), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n536_), .ZN(new_n545_));
  NOR3_X1   g344(.A1(new_n518_), .A2(new_n519_), .A3(new_n517_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n508_), .B1(new_n507_), .B2(new_n515_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n545_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n530_), .A2(KEYINPUT15), .A3(new_n535_), .ZN(new_n549_));
  AOI21_X1  g348(.A(KEYINPUT15), .B1(new_n530_), .B2(new_n535_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n516_), .B(new_n520_), .C1(new_n549_), .C2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n548_), .A2(new_n551_), .A3(new_n498_), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n539_), .A2(new_n544_), .A3(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n544_), .B1(new_n539_), .B2(new_n552_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n497_), .A2(new_n555_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n400_), .A2(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n436_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n466_), .A2(new_n545_), .A3(new_n419_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT71), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G232gat), .A2(G233gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT34), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT35), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n558_), .A2(new_n559_), .A3(new_n560_), .A4(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n564_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n558_), .A2(new_n559_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n565_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n569_), .B1(new_n558_), .B2(KEYINPUT71), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n566_), .B1(new_n568_), .B2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G190gat), .B(G218gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G134gat), .B(G162gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n574_), .A2(KEYINPUT36), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n574_), .A2(KEYINPUT36), .ZN(new_n576_));
  OR3_X1    g375(.A1(new_n571_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n571_), .A2(KEYINPUT72), .A3(new_n575_), .ZN(new_n578_));
  AOI21_X1  g377(.A(KEYINPUT72), .B1(new_n571_), .B2(new_n575_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n577_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT37), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n577_), .B(KEYINPUT37), .C1(new_n579_), .C2(new_n578_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G127gat), .B(G155gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G183gat), .B(G211gat), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(KEYINPUT77), .B(KEYINPUT17), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n587_), .A2(new_n588_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n589_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT78), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT78), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n589_), .A2(new_n594_), .A3(new_n591_), .A4(new_n590_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n516_), .A2(new_n520_), .ZN(new_n597_));
  AND2_X1   g396(.A1(G231gat), .A2(G233gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n448_), .B(new_n598_), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n597_), .A2(new_n599_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n596_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n591_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n587_), .A2(new_n588_), .ZN(new_n604_));
  OAI21_X1  g403(.A(KEYINPUT17), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT17), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n589_), .A2(new_n606_), .A3(new_n591_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n597_), .A2(new_n599_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n597_), .A2(new_n599_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n608_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n602_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT79), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT79), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n602_), .A2(new_n611_), .A3(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n584_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n557_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(new_n501_), .A3(new_n364_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT38), .ZN(new_n622_));
  INV_X1    g421(.A(new_n378_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n397_), .A2(new_n332_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n328_), .A2(new_n331_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n321_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n627_), .A2(new_n277_), .A3(new_n396_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n624_), .A2(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n623_), .B1(new_n629_), .B2(new_n376_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n580_), .B(KEYINPUT100), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT101), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n632_), .A2(KEYINPUT101), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n556_), .B(KEYINPUT99), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n637_), .A2(new_n616_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n636_), .A2(new_n364_), .A3(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(G1gat), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n622_), .A2(new_n640_), .ZN(G1324gat));
  INV_X1    g440(.A(new_n277_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n620_), .A2(new_n642_), .A3(new_n500_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n642_), .B(new_n638_), .C1(new_n634_), .C2(new_n635_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT39), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n644_), .A2(new_n645_), .A3(G8gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n644_), .B2(G8gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n643_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT40), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  OAI211_X1 g449(.A(KEYINPUT40), .B(new_n643_), .C1(new_n646_), .C2(new_n647_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1325gat));
  NAND3_X1  g451(.A1(new_n620_), .A2(new_n372_), .A3(new_n399_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n636_), .A2(new_n399_), .A3(new_n638_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n654_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT41), .B1(new_n654_), .B2(G15gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n653_), .B1(new_n655_), .B2(new_n656_), .ZN(G1326gat));
  NOR2_X1   g456(.A1(new_n332_), .A2(G22gat), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT102), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n620_), .A2(new_n659_), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n627_), .B(new_n638_), .C1(new_n634_), .C2(new_n635_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n661_), .A2(new_n662_), .A3(G22gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n662_), .B1(new_n661_), .B2(G22gat), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n660_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT103), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  OAI211_X1 g466(.A(KEYINPUT103), .B(new_n660_), .C1(new_n663_), .C2(new_n664_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1327gat));
  INV_X1    g468(.A(new_n631_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n670_), .A2(new_n616_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n557_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n673_), .A2(new_n527_), .A3(new_n364_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n399_), .B1(new_n624_), .B2(new_n628_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n675_), .B(new_n584_), .C1(new_n676_), .C2(new_n623_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n400_), .A2(KEYINPUT104), .A3(new_n675_), .A4(new_n584_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n584_), .ZN(new_n681_));
  OAI21_X1  g480(.A(KEYINPUT43), .B1(new_n630_), .B2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n679_), .A2(new_n680_), .A3(new_n682_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n637_), .A2(new_n617_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n683_), .A2(new_n684_), .A3(KEYINPUT44), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT44), .B1(new_n683_), .B2(new_n684_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT105), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(new_n688_), .A3(new_n364_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G29gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n688_), .B1(new_n687_), .B2(new_n364_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n674_), .B1(new_n690_), .B2(new_n691_), .ZN(G1328gat));
  NAND4_X1  g491(.A1(new_n557_), .A2(new_n525_), .A3(new_n642_), .A4(new_n671_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT45), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n685_), .A2(new_n686_), .A3(new_n277_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n696_), .B1(new_n697_), .B2(new_n525_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n699_));
  NOR2_X1   g498(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT107), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n698_), .A2(new_n699_), .A3(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n701_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n683_), .A2(new_n684_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n683_), .A2(new_n684_), .A3(KEYINPUT44), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n706_), .A2(new_n642_), .A3(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n695_), .B1(new_n708_), .B2(G36gat), .ZN(new_n709_));
  INV_X1    g508(.A(new_n699_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n703_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n702_), .A2(new_n711_), .ZN(G1329gat));
  AOI21_X1  g511(.A(G43gat), .B1(new_n673_), .B2(new_n399_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n376_), .A2(new_n366_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n687_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT47), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n715_), .B(new_n716_), .ZN(G1330gat));
  AOI21_X1  g516(.A(G50gat), .B1(new_n673_), .B2(new_n627_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n627_), .A2(G50gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n687_), .B2(new_n719_), .ZN(G1331gat));
  NAND3_X1  g519(.A1(new_n555_), .A2(new_n613_), .A3(new_n615_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n496_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n636_), .A2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(G57gat), .B1(new_n723_), .B2(new_n396_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n555_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n630_), .A2(new_n725_), .A3(new_n496_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(new_n618_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n727_), .A2(new_n443_), .A3(new_n364_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n724_), .A2(new_n728_), .ZN(G1332gat));
  NAND3_X1  g528(.A1(new_n727_), .A2(new_n441_), .A3(new_n642_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n636_), .A2(new_n642_), .A3(new_n722_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT48), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n731_), .A2(new_n732_), .A3(G64gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n731_), .B2(G64gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n730_), .B1(new_n733_), .B2(new_n734_), .ZN(G1333gat));
  INV_X1    g534(.A(G71gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n727_), .A2(new_n736_), .A3(new_n399_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n636_), .A2(new_n399_), .A3(new_n722_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(KEYINPUT108), .B(KEYINPUT49), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n738_), .A2(G71gat), .A3(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n738_), .B2(G71gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n740_), .B2(new_n741_), .ZN(G1334gat));
  INV_X1    g541(.A(G78gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n727_), .A2(new_n743_), .A3(new_n627_), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n627_), .B(new_n722_), .C1(new_n634_), .C2(new_n635_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n745_), .A2(G78gat), .A3(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n745_), .B2(G78gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  OAI211_X1 g550(.A(KEYINPUT110), .B(new_n744_), .C1(new_n747_), .C2(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1335gat));
  NOR3_X1   g552(.A1(new_n496_), .A2(new_n616_), .A3(new_n725_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n683_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT111), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n755_), .B(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(G85gat), .B1(new_n757_), .B2(new_n396_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n726_), .A2(new_n671_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n759_), .A2(new_n407_), .A3(new_n364_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1336gat));
  AND2_X1   g560(.A1(new_n759_), .A2(new_n642_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n762_), .A2(G92gat), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n408_), .A2(new_n409_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n642_), .A2(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n763_), .B1(new_n757_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT112), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  OAI211_X1 g567(.A(KEYINPUT112), .B(new_n763_), .C1(new_n757_), .C2(new_n765_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(G1337gat));
  OAI21_X1  g569(.A(G99gat), .B1(new_n755_), .B2(new_n376_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n759_), .A2(new_n399_), .A3(new_n412_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g573(.A1(new_n759_), .A2(new_n413_), .A3(new_n627_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n683_), .A2(new_n627_), .A3(new_n754_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777_));
  AND4_X1   g576(.A1(KEYINPUT113), .A2(new_n776_), .A3(new_n777_), .A4(G106gat), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n413_), .B1(new_n779_), .B2(KEYINPUT52), .ZN(new_n780_));
  AOI22_X1  g579(.A1(new_n776_), .A2(new_n780_), .B1(KEYINPUT113), .B2(new_n777_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n775_), .B1(new_n778_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT53), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n784_), .B(new_n775_), .C1(new_n778_), .C2(new_n781_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(G1339gat));
  INV_X1    g585(.A(KEYINPUT121), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT59), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n616_), .A2(KEYINPUT114), .A3(new_n555_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n721_), .A2(new_n791_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n490_), .A2(new_n681_), .A3(new_n789_), .A4(new_n793_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n582_), .A2(new_n790_), .A3(new_n583_), .A4(new_n792_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT54), .B1(new_n493_), .B2(new_n795_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT57), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n498_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n548_), .A2(new_n551_), .A3(new_n499_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n542_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n542_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n802_), .B1(new_n539_), .B2(new_n552_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n801_), .A2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n482_), .B2(new_n486_), .ZN(new_n805_));
  AOI211_X1 g604(.A(KEYINPUT115), .B(new_n555_), .C1(new_n476_), .C2(new_n481_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT115), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n482_), .B2(new_n725_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n459_), .A2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n485_), .A2(KEYINPUT55), .ZN(new_n812_));
  OAI21_X1  g611(.A(KEYINPUT116), .B1(new_n455_), .B2(new_n458_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n452_), .A2(new_n814_), .A3(new_n457_), .A4(new_n454_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n811_), .A2(new_n812_), .A3(new_n813_), .A4(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n483_), .ZN(new_n817_));
  AOI21_X1  g616(.A(KEYINPUT56), .B1(new_n817_), .B2(KEYINPUT117), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT117), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT56), .ZN(new_n820_));
  AOI211_X1 g619(.A(new_n819_), .B(new_n820_), .C1(new_n816_), .C2(new_n483_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n818_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n805_), .B1(new_n809_), .B2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n798_), .B1(new_n823_), .B2(new_n631_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n485_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n480_), .B1(new_n825_), .B2(new_n474_), .ZN(new_n826_));
  NOR4_X1   g625(.A1(new_n484_), .A2(KEYINPUT68), .A3(new_n485_), .A4(new_n483_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n725_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT115), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n482_), .A2(new_n807_), .A3(new_n725_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n813_), .A2(new_n815_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT55), .B1(new_n455_), .B2(new_n458_), .ZN(new_n832_));
  AOI211_X1 g631(.A(new_n810_), .B(new_n457_), .C1(new_n452_), .C2(new_n454_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n474_), .B1(new_n831_), .B2(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n820_), .B1(new_n835_), .B2(new_n819_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n817_), .A2(KEYINPUT117), .A3(KEYINPUT56), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n829_), .A2(new_n830_), .A3(new_n836_), .A4(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n805_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n840_), .A2(KEYINPUT57), .A3(new_n670_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n835_), .A2(new_n820_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n817_), .A2(KEYINPUT56), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n804_), .B1(new_n476_), .B2(new_n481_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n842_), .A2(new_n843_), .A3(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT58), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(KEYINPUT118), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(KEYINPUT118), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n842_), .A2(new_n843_), .A3(new_n848_), .A4(new_n844_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n847_), .A2(new_n584_), .A3(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n824_), .A2(new_n841_), .A3(new_n850_), .ZN(new_n851_));
  AOI211_X1 g650(.A(KEYINPUT119), .B(new_n797_), .C1(new_n851_), .C2(new_n617_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n631_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n850_), .B1(new_n854_), .B2(KEYINPUT57), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n823_), .A2(new_n798_), .A3(new_n631_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n617_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n797_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n853_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n852_), .A2(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n642_), .A2(new_n627_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n396_), .A2(new_n376_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n788_), .B1(new_n860_), .B2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT120), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n856_), .B1(new_n855_), .B2(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n824_), .A2(KEYINPUT120), .A3(new_n850_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n616_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n788_), .B(new_n864_), .C1(new_n869_), .C2(new_n797_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n787_), .B1(new_n865_), .B2(new_n871_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n852_), .A2(new_n859_), .A3(new_n863_), .ZN(new_n873_));
  OAI211_X1 g672(.A(KEYINPUT121), .B(new_n870_), .C1(new_n873_), .C2(new_n788_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n872_), .A2(new_n725_), .A3(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(G113gat), .ZN(new_n876_));
  INV_X1    g675(.A(new_n873_), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n555_), .A2(G113gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n876_), .B1(new_n877_), .B2(new_n878_), .ZN(G1340gat));
  INV_X1    g678(.A(G120gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(new_n496_), .B2(KEYINPUT60), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n873_), .B(new_n881_), .C1(KEYINPUT60), .C2(new_n880_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n497_), .B(new_n870_), .C1(new_n873_), .C2(new_n788_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n882_), .B1(new_n884_), .B2(new_n880_), .ZN(G1341gat));
  NAND3_X1  g684(.A1(new_n872_), .A2(new_n616_), .A3(new_n874_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(G127gat), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n617_), .A2(G127gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n877_), .B2(new_n888_), .ZN(G1342gat));
  NAND3_X1  g688(.A1(new_n872_), .A2(new_n584_), .A3(new_n874_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(G134gat), .ZN(new_n891_));
  OR3_X1    g690(.A1(new_n877_), .A2(G134gat), .A3(new_n670_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(KEYINPUT122), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n891_), .A2(new_n895_), .A3(new_n892_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(G1343gat));
  NAND4_X1  g696(.A1(new_n627_), .A2(new_n277_), .A3(new_n364_), .A4(new_n376_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n852_), .A2(new_n859_), .A3(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n725_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n497_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g702(.A1(new_n899_), .A2(new_n616_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(KEYINPUT61), .B(G155gat), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n904_), .B(new_n905_), .ZN(G1346gat));
  INV_X1    g705(.A(G162gat), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n899_), .A2(new_n907_), .A3(new_n631_), .ZN(new_n908_));
  AND2_X1   g707(.A1(new_n899_), .A2(new_n584_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n909_), .B2(new_n907_), .ZN(G1347gat));
  NOR3_X1   g709(.A1(new_n277_), .A2(new_n364_), .A3(new_n376_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n725_), .ZN(new_n912_));
  XOR2_X1   g711(.A(new_n912_), .B(KEYINPUT123), .Z(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n332_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n869_), .A2(new_n797_), .ZN(new_n915_));
  OAI21_X1  g714(.A(G169gat), .B1(new_n914_), .B2(new_n915_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(KEYINPUT62), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n911_), .A2(new_n332_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n915_), .A2(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n921_));
  AND2_X1   g720(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n725_), .B1(new_n921_), .B2(new_n922_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n917_), .B1(new_n920_), .B2(new_n923_), .ZN(G1348gat));
  NAND3_X1  g723(.A1(new_n860_), .A2(new_n332_), .A3(new_n911_), .ZN(new_n925_));
  INV_X1    g724(.A(G176gat), .ZN(new_n926_));
  NOR3_X1   g725(.A1(new_n925_), .A2(new_n926_), .A3(new_n496_), .ZN(new_n927_));
  AOI21_X1  g726(.A(G176gat), .B1(new_n919_), .B2(new_n497_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n927_), .A2(new_n928_), .ZN(G1349gat));
  NOR3_X1   g728(.A1(new_n920_), .A2(new_n230_), .A3(new_n617_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n925_), .A2(new_n617_), .ZN(new_n931_));
  OR2_X1    g730(.A1(new_n931_), .A2(KEYINPUT124), .ZN(new_n932_));
  AOI21_X1  g731(.A(G183gat), .B1(new_n931_), .B2(KEYINPUT124), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n930_), .B1(new_n932_), .B2(new_n933_), .ZN(G1350gat));
  OAI21_X1  g733(.A(G190gat), .B1(new_n920_), .B2(new_n681_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n919_), .A2(new_n229_), .A3(new_n631_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(G1351gat));
  NAND3_X1  g736(.A1(new_n379_), .A2(new_n642_), .A3(new_n376_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n938_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n860_), .A2(new_n939_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n860_), .A2(KEYINPUT125), .A3(new_n939_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(new_n725_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(KEYINPUT126), .B(G197gat), .ZN(new_n946_));
  XOR2_X1   g745(.A(new_n945_), .B(new_n946_), .Z(G1352gat));
  NAND2_X1  g746(.A1(new_n944_), .A2(new_n497_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g748(.A(new_n617_), .B1(new_n942_), .B2(new_n943_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n951_));
  AND2_X1   g750(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n950_), .B1(new_n951_), .B2(new_n952_), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n953_), .B1(new_n950_), .B2(new_n951_), .ZN(G1354gat));
  INV_X1    g753(.A(KEYINPUT127), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n681_), .B1(new_n942_), .B2(new_n943_), .ZN(new_n956_));
  INV_X1    g755(.A(G218gat), .ZN(new_n957_));
  OR2_X1    g756(.A1(new_n956_), .A2(new_n957_), .ZN(new_n958_));
  NAND3_X1  g757(.A1(new_n944_), .A2(new_n957_), .A3(new_n631_), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n955_), .B1(new_n958_), .B2(new_n959_), .ZN(new_n960_));
  OAI211_X1 g759(.A(new_n959_), .B(new_n955_), .C1(new_n956_), .C2(new_n957_), .ZN(new_n961_));
  INV_X1    g760(.A(new_n961_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n960_), .A2(new_n962_), .ZN(G1355gat));
endmodule


