//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 0 0 1 0 0 0 1 0 1 0 1 1 0 1 0 1 0 1 0 0 1 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n891_, new_n892_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n907_, new_n909_, new_n910_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  AND2_X1   g001(.A1(new_n202_), .A2(KEYINPUT70), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(KEYINPUT70), .ZN(new_n204_));
  XOR2_X1   g003(.A(G43gat), .B(G50gat), .Z(new_n205_));
  OR3_X1    g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n205_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G15gat), .B(G22gat), .ZN(new_n209_));
  INV_X1    g008(.A(G1gat), .ZN(new_n210_));
  INV_X1    g009(.A(G8gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT14), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G1gat), .B(G8gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n208_), .B(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT76), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(G229gat), .A3(G233gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT15), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n208_), .B(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n215_), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G229gat), .A2(G233gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n208_), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n222_), .B(new_n223_), .C1(new_n215_), .C2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n218_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G113gat), .B(G141gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G169gat), .B(G197gat), .ZN(new_n228_));
  XOR2_X1   g027(.A(new_n227_), .B(new_n228_), .Z(new_n229_));
  OR2_X1    g028(.A1(new_n229_), .A2(KEYINPUT77), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n226_), .B(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G22gat), .B(G50gat), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT28), .ZN(new_n234_));
  AND2_X1   g033(.A1(G155gat), .A2(G162gat), .ZN(new_n235_));
  NOR2_X1   g034(.A1(G155gat), .A2(G162gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(G141gat), .A2(G148gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  AND2_X1   g042(.A1(G141gat), .A2(G148gat), .ZN(new_n244_));
  NOR3_X1   g043(.A1(new_n244_), .A2(KEYINPUT84), .A3(KEYINPUT2), .ZN(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT84), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n240_), .B(new_n243_), .C1(new_n245_), .C2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT83), .ZN(new_n250_));
  NOR3_X1   g049(.A1(new_n235_), .A2(new_n236_), .A3(KEYINPUT1), .ZN(new_n251_));
  INV_X1    g050(.A(G141gat), .ZN(new_n252_));
  INV_X1    g051(.A(G148gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G141gat), .A2(G148gat), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n254_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n250_), .B1(new_n251_), .B2(new_n257_), .ZN(new_n258_));
  OR2_X1    g057(.A1(G155gat), .A2(G162gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT1), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G155gat), .A2(G162gat), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n244_), .A2(new_n241_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n262_), .A2(new_n263_), .A3(KEYINPUT83), .A4(new_n255_), .ZN(new_n264_));
  AOI22_X1  g063(.A1(new_n237_), .A2(new_n249_), .B1(new_n258_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT29), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n234_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n258_), .A2(new_n264_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n246_), .B(KEYINPUT84), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n243_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n237_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  AND4_X1   g070(.A1(new_n234_), .A2(new_n268_), .A3(new_n271_), .A4(new_n266_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n233_), .B1(new_n267_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n268_), .A2(new_n271_), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT28), .B1(new_n274_), .B2(KEYINPUT29), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n265_), .A2(new_n234_), .A3(new_n266_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(new_n276_), .A3(new_n232_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n273_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G228gat), .A2(G233gat), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n266_), .B1(new_n268_), .B2(new_n271_), .ZN(new_n281_));
  OR2_X1    g080(.A1(G197gat), .A2(G204gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G197gat), .A2(G204gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT21), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n282_), .A2(KEYINPUT21), .A3(new_n283_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G211gat), .B(G218gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n286_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n287_), .A2(new_n288_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n280_), .B1(new_n281_), .B2(new_n292_), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n279_), .B(new_n291_), .C1(new_n265_), .C2(new_n266_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G78gat), .B(G106gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT85), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n293_), .A2(new_n294_), .A3(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n296_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n278_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT86), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT86), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n278_), .B(new_n301_), .C1(new_n297_), .C2(new_n298_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n278_), .A2(new_n297_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT87), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n293_), .A2(new_n294_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n305_), .B1(new_n306_), .B2(new_n295_), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n306_), .A2(new_n305_), .A3(new_n295_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n304_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n303_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT88), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n303_), .A2(new_n309_), .A3(KEYINPUT88), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT27), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT26), .B(G190gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT25), .B(G183gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G183gat), .A2(G190gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT23), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT23), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n321_), .A2(G183gat), .A3(G190gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(G169gat), .A2(G176gat), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT24), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n318_), .A2(new_n323_), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G169gat), .A2(G176gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT24), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n329_), .A2(KEYINPUT89), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT89), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n331_), .B1(new_n328_), .B2(KEYINPUT24), .ZN(new_n332_));
  NOR3_X1   g131(.A1(new_n330_), .A2(new_n324_), .A3(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT90), .B1(new_n327_), .B2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n332_), .A2(new_n324_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n335_), .B1(KEYINPUT89), .B2(new_n329_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT90), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n323_), .A2(new_n326_), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n336_), .A2(new_n337_), .A3(new_n318_), .A4(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT22), .B(G169gat), .ZN(new_n340_));
  INV_X1    g139(.A(G176gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n328_), .A2(KEYINPUT91), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n328_), .A2(KEYINPUT91), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n342_), .A2(new_n345_), .ZN(new_n346_));
  AND3_X1   g145(.A1(new_n319_), .A2(KEYINPUT80), .A3(KEYINPUT23), .ZN(new_n347_));
  AOI21_X1  g146(.A(KEYINPUT80), .B1(new_n319_), .B2(KEYINPUT23), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n322_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(G183gat), .A2(G190gat), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n346_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n334_), .A2(new_n339_), .A3(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n291_), .ZN(new_n355_));
  OR2_X1    g154(.A1(KEYINPUT78), .A2(G183gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(KEYINPUT78), .A2(G183gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n323_), .B1(new_n358_), .B2(G190gat), .ZN(new_n359_));
  INV_X1    g158(.A(G169gat), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT22), .B1(new_n360_), .B2(KEYINPUT81), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n360_), .A2(KEYINPUT22), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n341_), .B(new_n361_), .C1(new_n362_), .C2(KEYINPUT81), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n359_), .A2(new_n363_), .A3(new_n328_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT25), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n365_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n316_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n360_), .A2(new_n341_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n369_), .A2(KEYINPUT24), .A3(new_n328_), .ZN(new_n370_));
  AOI22_X1  g169(.A1(new_n370_), .A2(KEYINPUT79), .B1(new_n325_), .B2(new_n324_), .ZN(new_n371_));
  OR3_X1    g170(.A1(new_n329_), .A2(KEYINPUT79), .A3(new_n324_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n368_), .A2(new_n371_), .A3(new_n372_), .A4(new_n349_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n292_), .A2(new_n364_), .A3(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n355_), .A2(KEYINPUT20), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G226gat), .A2(G233gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT19), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT20), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n373_), .A2(new_n364_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n379_), .B1(new_n380_), .B2(new_n291_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n336_), .A2(new_n318_), .A3(new_n338_), .ZN(new_n382_));
  AOI22_X1  g181(.A1(new_n382_), .A2(KEYINPUT90), .B1(new_n352_), .B2(new_n346_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n383_), .A2(new_n292_), .A3(new_n339_), .ZN(new_n384_));
  AOI22_X1  g183(.A1(new_n375_), .A2(new_n377_), .B1(new_n381_), .B2(new_n384_), .ZN(new_n385_));
  XOR2_X1   g184(.A(G8gat), .B(G36gat), .Z(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G64gat), .B(G92gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n315_), .B1(new_n385_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT98), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n289_), .B(new_n290_), .C1(new_n327_), .C2(new_n333_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n345_), .A2(new_n342_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n395_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n393_), .B(KEYINPUT20), .C1(new_n394_), .C2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n380_), .A2(new_n291_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n292_), .A2(new_n353_), .A3(new_n382_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n393_), .B1(new_n400_), .B2(KEYINPUT20), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n377_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n355_), .A2(KEYINPUT20), .A3(new_n378_), .A4(new_n374_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(new_n390_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n392_), .A2(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n292_), .B1(new_n383_), .B2(new_n339_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n374_), .A2(KEYINPUT20), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n377_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n384_), .A2(new_n381_), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n409_), .A2(new_n391_), .A3(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n391_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n315_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n406_), .A2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n314_), .A2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G127gat), .B(G134gat), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G113gat), .B(G120gat), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n416_), .A2(new_n418_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n268_), .A2(new_n271_), .A3(new_n422_), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n420_), .A2(KEYINPUT82), .A3(new_n421_), .ZN(new_n424_));
  AOI21_X1  g223(.A(KEYINPUT82), .B1(new_n420_), .B2(new_n421_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  OAI211_X1 g225(.A(KEYINPUT4), .B(new_n423_), .C1(new_n426_), .C2(new_n265_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT93), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n274_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT93), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n429_), .A2(new_n430_), .A3(KEYINPUT4), .A4(new_n423_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G225gat), .A2(G233gat), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n434_), .B1(new_n429_), .B2(KEYINPUT4), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n432_), .A2(new_n436_), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n429_), .A2(new_n423_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n433_), .ZN(new_n439_));
  XOR2_X1   g238(.A(G1gat), .B(G29gat), .Z(new_n440_));
  XNOR2_X1  g239(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G57gat), .B(G85gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n437_), .A2(new_n439_), .A3(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n435_), .B1(new_n428_), .B2(new_n431_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n439_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n444_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n446_), .A2(new_n449_), .A3(KEYINPUT99), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT99), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n451_), .B(new_n444_), .C1(new_n447_), .C2(new_n448_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G227gat), .A2(G233gat), .ZN(new_n455_));
  XOR2_X1   g254(.A(new_n455_), .B(G15gat), .Z(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT30), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n380_), .B(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(new_n426_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G71gat), .B(G99gat), .ZN(new_n460_));
  INV_X1    g259(.A(G43gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT31), .ZN(new_n463_));
  OR2_X1    g262(.A1(new_n459_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n459_), .A2(new_n463_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n454_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n415_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n466_), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n406_), .A2(new_n413_), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n303_), .A2(KEYINPUT88), .A3(new_n309_), .ZN(new_n472_));
  AOI21_X1  g271(.A(KEYINPUT88), .B1(new_n303_), .B2(new_n309_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n453_), .B(new_n471_), .C1(new_n472_), .C2(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n472_), .A2(new_n473_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n391_), .A2(KEYINPUT32), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n409_), .A2(new_n410_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n476_), .B1(new_n477_), .B2(KEYINPUT97), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n409_), .A2(KEYINPUT97), .A3(new_n410_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n402_), .A2(KEYINPUT32), .A3(new_n391_), .A4(new_n403_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n478_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n450_), .A2(new_n481_), .A3(new_n452_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT33), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n446_), .A2(new_n483_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n432_), .B(new_n433_), .C1(KEYINPUT4), .C2(new_n429_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n429_), .A2(KEYINPUT95), .A3(new_n423_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n434_), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT95), .B1(new_n429_), .B2(new_n423_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n444_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT96), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT96), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n491_), .B(new_n444_), .C1(new_n487_), .C2(new_n488_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n485_), .A2(new_n490_), .A3(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n411_), .A2(new_n412_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n437_), .A2(KEYINPUT33), .A3(new_n439_), .A4(new_n445_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n484_), .A2(new_n493_), .A3(new_n494_), .A4(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n482_), .A2(new_n496_), .ZN(new_n497_));
  AOI22_X1  g296(.A1(new_n474_), .A2(KEYINPUT100), .B1(new_n475_), .B2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n414_), .B1(new_n452_), .B2(new_n450_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT100), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n314_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n470_), .B1(new_n498_), .B2(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n469_), .B1(new_n502_), .B2(KEYINPUT101), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n471_), .A2(new_n453_), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT100), .B1(new_n475_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n475_), .A2(new_n497_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(new_n501_), .A3(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT101), .B1(new_n507_), .B2(new_n466_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n231_), .B1(new_n503_), .B2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G190gat), .B(G218gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G134gat), .B(G162gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n513_), .B(KEYINPUT36), .Z(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G85gat), .B(G92gat), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT9), .ZN(new_n518_));
  XOR2_X1   g317(.A(KEYINPUT10), .B(G99gat), .Z(new_n519_));
  INV_X1    g318(.A(G106gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(G85gat), .ZN(new_n522_));
  INV_X1    g321(.A(G92gat), .ZN(new_n523_));
  OR3_X1    g322(.A1(new_n522_), .A2(new_n523_), .A3(KEYINPUT9), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G99gat), .A2(G106gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT6), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n518_), .A2(new_n521_), .A3(new_n524_), .A4(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT8), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT65), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n529_), .ZN(new_n530_));
  OR2_X1    g329(.A1(G99gat), .A2(G106gat), .ZN(new_n531_));
  NOR2_X1   g330(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n525_), .A2(KEYINPUT6), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n525_), .A2(KEYINPUT6), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(KEYINPUT65), .A3(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n530_), .A2(new_n533_), .A3(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n528_), .B1(new_n537_), .B2(new_n517_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT66), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  AOI211_X1 g340(.A(KEYINPUT8), .B(new_n516_), .C1(new_n533_), .C2(new_n526_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n543_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n527_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n220_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n546_), .B1(new_n208_), .B2(new_n545_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n547_), .A2(KEYINPUT35), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G232gat), .A2(G233gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n552_), .B1(new_n547_), .B2(KEYINPUT71), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n548_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n547_), .A2(KEYINPUT71), .A3(new_n552_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n515_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n555_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n557_), .B1(new_n548_), .B2(new_n553_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n513_), .A2(KEYINPUT36), .ZN(new_n559_));
  AOI22_X1  g358(.A1(new_n556_), .A2(KEYINPUT72), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n554_), .A2(new_n555_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n514_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT72), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(KEYINPUT37), .B1(new_n560_), .B2(new_n564_), .ZN(new_n565_));
  AND3_X1   g364(.A1(new_n554_), .A2(new_n555_), .A3(new_n559_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT37), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n566_), .A2(new_n556_), .A3(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(G127gat), .B(G155gat), .Z(new_n569_));
  XNOR2_X1  g368(.A(G183gat), .B(G211gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT17), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n573_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n576_), .A2(KEYINPUT17), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G231gat), .A2(G233gat), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n578_), .B(KEYINPUT73), .Z(new_n579_));
  XNOR2_X1  g378(.A(new_n215_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G57gat), .B(G64gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT11), .ZN(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT67), .B(G71gat), .ZN(new_n583_));
  INV_X1    g382(.A(G78gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n582_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n583_), .B(G78gat), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n581_), .A2(KEYINPUT11), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n586_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  AOI211_X1 g390(.A(new_n575_), .B(new_n577_), .C1(new_n580_), .C2(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n592_), .B1(new_n580_), .B2(new_n591_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n590_), .B(KEYINPUT68), .ZN(new_n594_));
  INV_X1    g393(.A(new_n580_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(KEYINPUT75), .B(KEYINPUT17), .Z(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(new_n597_), .A3(new_n576_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n593_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NOR3_X1   g399(.A1(new_n565_), .A2(new_n568_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT12), .ZN(new_n602_));
  INV_X1    g401(.A(new_n527_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n537_), .A2(new_n517_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT8), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n542_), .B1(new_n605_), .B2(KEYINPUT66), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n603_), .B1(new_n606_), .B2(new_n540_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n602_), .B1(new_n607_), .B2(new_n591_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(G230gat), .A2(G233gat), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n527_), .B(new_n591_), .C1(new_n541_), .C2(new_n544_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n545_), .A2(KEYINPUT12), .A3(new_n594_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n608_), .A2(new_n609_), .A3(new_n610_), .A4(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n545_), .B(new_n591_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n614_), .A2(new_n609_), .ZN(new_n615_));
  XOR2_X1   g414(.A(G120gat), .B(G148gat), .Z(new_n616_));
  XNOR2_X1  g415(.A(G176gat), .B(G204gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n613_), .A2(new_n615_), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n620_), .B1(new_n613_), .B2(new_n615_), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n622_), .A2(KEYINPUT13), .A3(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(KEYINPUT13), .B1(new_n622_), .B2(new_n623_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n510_), .A2(new_n601_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(new_n210_), .A3(new_n454_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT38), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n556_), .A2(KEYINPUT72), .ZN(new_n632_));
  AOI211_X1 g431(.A(new_n563_), .B(new_n515_), .C1(new_n554_), .C2(new_n555_), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n632_), .A2(new_n633_), .A3(new_n566_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n634_), .B1(new_n503_), .B2(new_n509_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n626_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n636_), .A2(new_n231_), .A3(new_n600_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(G1gat), .B1(new_n638_), .B2(new_n453_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n629_), .A2(new_n630_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n640_), .A2(KEYINPUT102), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n640_), .A2(KEYINPUT102), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n631_), .B(new_n639_), .C1(new_n641_), .C2(new_n642_), .ZN(G1324gat));
  NAND3_X1  g442(.A1(new_n628_), .A2(new_n211_), .A3(new_n414_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n635_), .A2(new_n414_), .A3(new_n637_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(new_n646_), .A3(G8gat), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n646_), .B1(new_n645_), .B2(G8gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n644_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n650_), .B(KEYINPUT40), .Z(G1325gat));
  NOR3_X1   g450(.A1(new_n627_), .A2(G15gat), .A3(new_n466_), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n652_), .A2(KEYINPUT103), .ZN(new_n653_));
  OAI21_X1  g452(.A(G15gat), .B1(new_n638_), .B2(new_n466_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT41), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n654_), .A2(KEYINPUT41), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n652_), .A2(KEYINPUT103), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n653_), .A2(new_n655_), .A3(new_n656_), .A4(new_n657_), .ZN(G1326gat));
  OAI21_X1  g457(.A(G22gat), .B1(new_n638_), .B2(new_n475_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT42), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n475_), .A2(G22gat), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n660_), .B1(new_n627_), .B2(new_n661_), .ZN(G1327gat));
  NAND2_X1  g461(.A1(new_n634_), .A2(new_n600_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n663_), .A2(new_n636_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n510_), .A2(new_n664_), .ZN(new_n665_));
  OR3_X1    g464(.A1(new_n665_), .A2(G29gat), .A3(new_n453_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667_));
  INV_X1    g466(.A(new_n231_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n626_), .A2(new_n668_), .A3(new_n600_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n560_), .A2(new_n564_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(new_n567_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n568_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n507_), .A2(KEYINPUT101), .A3(new_n466_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(new_n468_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n673_), .B1(new_n675_), .B2(new_n508_), .ZN(new_n676_));
  XOR2_X1   g475(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(KEYINPUT104), .A2(KEYINPUT43), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n673_), .B(new_n680_), .C1(new_n675_), .C2(new_n508_), .ZN(new_n681_));
  AOI211_X1 g480(.A(new_n667_), .B(new_n669_), .C1(new_n679_), .C2(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n565_), .A2(new_n568_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n683_), .B1(new_n503_), .B2(new_n509_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n681_), .B1(new_n684_), .B2(new_n677_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n669_), .ZN(new_n686_));
  AOI21_X1  g485(.A(KEYINPUT44), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n682_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT105), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n688_), .A2(new_n689_), .A3(new_n454_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(G29gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n689_), .B1(new_n688_), .B2(new_n454_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n666_), .B1(new_n691_), .B2(new_n692_), .ZN(G1328gat));
  INV_X1    g492(.A(KEYINPUT46), .ZN(new_n694_));
  INV_X1    g493(.A(G36gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n695_), .B1(new_n688_), .B2(new_n414_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n471_), .A2(G36gat), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n697_), .B1(new_n665_), .B2(new_n699_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n510_), .A2(KEYINPUT107), .A3(new_n664_), .A4(new_n698_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  XOR2_X1   g501(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n700_), .A2(new_n703_), .A3(new_n701_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n694_), .B1(new_n696_), .B2(new_n707_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n700_), .A2(new_n703_), .A3(new_n701_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n703_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n682_), .A2(new_n687_), .A3(new_n471_), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n711_), .B(KEYINPUT46), .C1(new_n695_), .C2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n708_), .A2(new_n713_), .ZN(G1329gat));
  OAI21_X1  g513(.A(new_n461_), .B1(new_n665_), .B2(new_n466_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT108), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  NOR4_X1   g516(.A1(new_n682_), .A2(new_n687_), .A3(new_n461_), .A4(new_n466_), .ZN(new_n718_));
  OAI21_X1  g517(.A(KEYINPUT47), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n688_), .A2(G43gat), .A3(new_n470_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT47), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n720_), .A2(new_n721_), .A3(new_n716_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n719_), .A2(new_n722_), .ZN(G1330gat));
  INV_X1    g522(.A(new_n665_), .ZN(new_n724_));
  AOI21_X1  g523(.A(G50gat), .B1(new_n724_), .B2(new_n314_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n314_), .A2(G50gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n688_), .B2(new_n726_), .ZN(G1331gat));
  NAND2_X1  g526(.A1(new_n601_), .A2(new_n636_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n728_), .B(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n668_), .B1(new_n503_), .B2(new_n509_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(G57gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(new_n733_), .A3(new_n454_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n635_), .A2(new_n231_), .A3(new_n599_), .A4(new_n636_), .ZN(new_n735_));
  OAI21_X1  g534(.A(G57gat), .B1(new_n735_), .B2(new_n453_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT110), .ZN(G1332gat));
  OAI21_X1  g537(.A(G64gat), .B1(new_n735_), .B2(new_n471_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT48), .ZN(new_n740_));
  INV_X1    g539(.A(G64gat), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n732_), .A2(new_n741_), .A3(new_n414_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(G1333gat));
  OAI21_X1  g542(.A(G71gat), .B1(new_n735_), .B2(new_n466_), .ZN(new_n744_));
  XOR2_X1   g543(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n745_));
  XNOR2_X1  g544(.A(new_n744_), .B(new_n745_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n466_), .A2(G71gat), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT112), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n732_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n746_), .A2(new_n749_), .ZN(G1334gat));
  OAI21_X1  g549(.A(G78gat), .B1(new_n735_), .B2(new_n475_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT50), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n732_), .A2(new_n584_), .A3(new_n314_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(G1335gat));
  NAND3_X1  g553(.A1(new_n636_), .A2(new_n231_), .A3(new_n600_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT113), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n685_), .A2(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(G85gat), .B1(new_n757_), .B2(new_n453_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n663_), .A2(new_n626_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n731_), .A2(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n760_), .A2(new_n522_), .A3(new_n454_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n758_), .A2(new_n761_), .ZN(G1336gat));
  OAI21_X1  g561(.A(G92gat), .B1(new_n757_), .B2(new_n471_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n760_), .A2(new_n523_), .A3(new_n414_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(G1337gat));
  NAND3_X1  g564(.A1(new_n685_), .A2(new_n470_), .A3(new_n756_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n470_), .A2(new_n519_), .ZN(new_n767_));
  AOI22_X1  g566(.A1(new_n766_), .A2(G99gat), .B1(new_n760_), .B2(new_n767_), .ZN(new_n768_));
  AND4_X1   g567(.A1(KEYINPUT114), .A2(new_n768_), .A3(KEYINPUT115), .A4(KEYINPUT51), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT51), .B1(new_n768_), .B2(KEYINPUT115), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n768_), .A2(KEYINPUT114), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n769_), .A2(new_n770_), .A3(new_n771_), .ZN(G1338gat));
  NAND3_X1  g571(.A1(new_n760_), .A2(new_n520_), .A3(new_n314_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n685_), .A2(new_n314_), .A3(new_n756_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n774_), .A2(new_n775_), .A3(G106gat), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n774_), .B2(G106gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT53), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n780_), .B(new_n773_), .C1(new_n776_), .C2(new_n777_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1339gat));
  XOR2_X1   g581(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n671_), .A2(new_n672_), .A3(new_n599_), .A4(new_n626_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n784_), .B1(new_n785_), .B2(new_n668_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n601_), .A2(new_n231_), .A3(new_n626_), .A4(new_n783_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n231_), .A2(new_n621_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT117), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT55), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n790_), .B1(new_n612_), .B2(new_n791_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n590_), .A2(KEYINPUT68), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n590_), .A2(KEYINPUT68), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT12), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n610_), .B1(new_n607_), .B2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT12), .B1(new_n545_), .B2(new_n590_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n798_), .A2(KEYINPUT117), .A3(KEYINPUT55), .A4(new_n609_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n608_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n609_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n791_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n792_), .B(new_n799_), .C1(new_n802_), .C2(new_n613_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n803_), .A2(KEYINPUT56), .A3(new_n620_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT56), .B1(new_n803_), .B2(new_n620_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n789_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n217_), .A2(new_n223_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n229_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT118), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n807_), .A2(KEYINPUT118), .A3(new_n808_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n223_), .B1(new_n208_), .B2(new_n221_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n222_), .A2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n811_), .A2(new_n812_), .A3(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n218_), .A2(new_n229_), .A3(new_n225_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n623_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n815_), .B(new_n816_), .C1(new_n817_), .C2(new_n621_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n634_), .B1(new_n806_), .B2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(KEYINPUT57), .B1(new_n819_), .B2(KEYINPUT119), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n822_));
  INV_X1    g621(.A(new_n818_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n803_), .A2(new_n620_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT56), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n803_), .A2(KEYINPUT56), .A3(new_n620_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n823_), .B1(new_n828_), .B2(new_n789_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n821_), .B(new_n822_), .C1(new_n829_), .C2(new_n634_), .ZN(new_n830_));
  OR2_X1    g629(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n827_), .A2(KEYINPUT120), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT120), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n803_), .A2(new_n833_), .A3(KEYINPUT56), .A4(new_n620_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n832_), .A2(new_n834_), .A3(new_n826_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n815_), .A2(new_n816_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n836_), .A2(new_n621_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n831_), .B1(new_n835_), .B2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n835_), .A2(new_n837_), .A3(new_n831_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n673_), .A2(new_n839_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n820_), .B(new_n830_), .C1(new_n838_), .C2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n788_), .B1(new_n841_), .B2(new_n600_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n415_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n843_), .A2(new_n466_), .A3(new_n453_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n842_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(G113gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(new_n847_), .A3(new_n668_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n820_), .A2(new_n830_), .ZN(new_n849_));
  OR2_X1    g648(.A1(new_n840_), .A2(new_n838_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n599_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  OAI211_X1 g650(.A(KEYINPUT59), .B(new_n844_), .C1(new_n851_), .C2(new_n788_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(new_n842_), .B2(new_n845_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n231_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n848_), .B1(new_n855_), .B2(new_n847_), .ZN(G1340gat));
  INV_X1    g655(.A(G120gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n626_), .B2(KEYINPUT60), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n846_), .B(new_n858_), .C1(KEYINPUT60), .C2(new_n857_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n626_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(new_n857_), .ZN(G1341gat));
  INV_X1    g660(.A(G127gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n846_), .A2(new_n862_), .A3(new_n599_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n600_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n862_), .ZN(G1342gat));
  INV_X1    g664(.A(G134gat), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n683_), .A2(new_n866_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(KEYINPUT122), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n841_), .A2(new_n600_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n788_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(KEYINPUT59), .B1(new_n871_), .B2(new_n844_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n842_), .A2(new_n853_), .A3(new_n845_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n868_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT123), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n846_), .A2(new_n634_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n866_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n874_), .A2(new_n875_), .A3(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n868_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n879_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n880_));
  AOI21_X1  g679(.A(G134gat), .B1(new_n846_), .B2(new_n634_), .ZN(new_n881_));
  OAI21_X1  g680(.A(KEYINPUT123), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n878_), .A2(new_n882_), .ZN(G1343gat));
  NAND4_X1  g682(.A1(new_n314_), .A2(new_n466_), .A3(new_n454_), .A4(new_n471_), .ZN(new_n884_));
  XOR2_X1   g683(.A(new_n884_), .B(KEYINPUT124), .Z(new_n885_));
  NAND2_X1  g684(.A1(new_n871_), .A2(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n886_), .A2(new_n231_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(new_n252_), .ZN(G1344gat));
  NOR2_X1   g687(.A1(new_n886_), .A2(new_n626_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(new_n253_), .ZN(G1345gat));
  NOR2_X1   g689(.A1(new_n886_), .A2(new_n600_), .ZN(new_n891_));
  XOR2_X1   g690(.A(KEYINPUT61), .B(G155gat), .Z(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(G1346gat));
  OAI21_X1  g692(.A(G162gat), .B1(new_n886_), .B2(new_n683_), .ZN(new_n894_));
  OR2_X1    g693(.A1(new_n670_), .A2(G162gat), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n886_), .B2(new_n895_), .ZN(G1347gat));
  INV_X1    g695(.A(KEYINPUT62), .ZN(new_n897_));
  NOR4_X1   g696(.A1(new_n314_), .A2(new_n466_), .A3(new_n454_), .A4(new_n471_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n871_), .A2(new_n898_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(new_n231_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n897_), .B1(new_n900_), .B2(new_n360_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n340_), .ZN(new_n902_));
  OAI211_X1 g701(.A(KEYINPUT62), .B(G169gat), .C1(new_n899_), .C2(new_n231_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n901_), .A2(new_n902_), .A3(new_n903_), .ZN(G1348gat));
  NOR2_X1   g703(.A1(new_n899_), .A2(new_n626_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(new_n341_), .ZN(G1349gat));
  NAND3_X1  g705(.A1(new_n871_), .A2(new_n599_), .A3(new_n898_), .ZN(new_n907_));
  MUX2_X1   g706(.A(new_n317_), .B(new_n358_), .S(new_n907_), .Z(G1350gat));
  OAI21_X1  g707(.A(G190gat), .B1(new_n899_), .B2(new_n683_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n634_), .A2(new_n316_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n909_), .B1(new_n899_), .B2(new_n910_), .ZN(G1351gat));
  NOR2_X1   g710(.A1(new_n471_), .A2(new_n470_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n912_), .A2(new_n314_), .A3(new_n453_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n842_), .A2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(new_n668_), .ZN(new_n915_));
  XOR2_X1   g714(.A(KEYINPUT125), .B(G197gat), .Z(new_n916_));
  XNOR2_X1  g715(.A(new_n915_), .B(new_n916_), .ZN(G1352gat));
  NAND2_X1  g716(.A1(new_n914_), .A2(new_n636_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g718(.A1(new_n914_), .A2(new_n599_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  AND2_X1   g720(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n920_), .A2(new_n921_), .A3(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n923_), .B1(new_n920_), .B2(new_n921_), .ZN(G1354gat));
  XOR2_X1   g723(.A(KEYINPUT126), .B(G218gat), .Z(new_n925_));
  NAND3_X1  g724(.A1(new_n914_), .A2(new_n673_), .A3(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n842_), .A2(new_n670_), .A3(new_n913_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n928_), .A2(new_n925_), .ZN(new_n929_));
  OAI21_X1  g728(.A(KEYINPUT127), .B1(new_n927_), .B2(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n926_), .B(new_n931_), .C1(new_n928_), .C2(new_n925_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n930_), .A2(new_n932_), .ZN(G1355gat));
endmodule


