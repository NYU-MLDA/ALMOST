//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 0 0 0 0 0 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 1 0 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 1 1 0 0 1 1 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n770_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n868_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n932_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT89), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G29gat), .B(G36gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G43gat), .B(G50gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT15), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G15gat), .B(G22gat), .ZN(new_n208_));
  INV_X1    g007(.A(G8gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G1gat), .B(G8gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n207_), .A2(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(new_n204_), .B(new_n205_), .Z(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT86), .ZN(new_n216_));
  XOR2_X1   g015(.A(new_n211_), .B(new_n212_), .Z(new_n217_));
  INV_X1    g016(.A(KEYINPUT86), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n206_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n216_), .A2(new_n217_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G229gat), .A2(G233gat), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n214_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT87), .ZN(new_n223_));
  INV_X1    g022(.A(new_n219_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n206_), .A2(new_n218_), .ZN(new_n225_));
  NOR3_X1   g024(.A1(new_n224_), .A2(new_n225_), .A3(new_n213_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n217_), .B1(new_n216_), .B2(new_n219_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n223_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n213_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(new_n220_), .A3(KEYINPUT87), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n221_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n222_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT88), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n203_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G113gat), .B(G141gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G169gat), .B(G197gat), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n236_), .B(new_n237_), .Z(new_n238_));
  AOI21_X1  g037(.A(KEYINPUT88), .B1(new_n238_), .B2(KEYINPUT89), .ZN(new_n239_));
  OAI22_X1  g038(.A1(new_n235_), .A2(new_n238_), .B1(new_n239_), .B2(new_n233_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT13), .ZN(new_n241_));
  NOR2_X1   g040(.A1(G85gat), .A2(G92gat), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  AND2_X1   g042(.A1(G85gat), .A2(G92gat), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n244_), .A2(new_n242_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n246_));
  AOI21_X1  g045(.A(KEYINPUT9), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT9), .ZN(new_n248_));
  NOR4_X1   g047(.A1(new_n244_), .A2(new_n242_), .A3(KEYINPUT68), .A4(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n243_), .B1(new_n247_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT6), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT70), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT70), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT6), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G99gat), .A2(G106gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n258_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n260_), .A2(new_n254_), .A3(new_n256_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT66), .B(G106gat), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT65), .ZN(new_n268_));
  NOR3_X1   g067(.A1(new_n266_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  OR2_X1    g068(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n270_));
  AOI21_X1  g069(.A(KEYINPUT65), .B1(new_n270_), .B2(new_n265_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n264_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n262_), .B1(new_n272_), .B2(KEYINPUT67), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT67), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n274_), .B(new_n264_), .C1(new_n269_), .C2(new_n271_), .ZN(new_n275_));
  OAI211_X1 g074(.A(KEYINPUT69), .B(new_n243_), .C1(new_n247_), .C2(new_n249_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n252_), .A2(new_n273_), .A3(new_n275_), .A4(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(KEYINPUT71), .A2(KEYINPUT7), .ZN(new_n278_));
  INV_X1    g077(.A(G99gat), .ZN(new_n279_));
  INV_X1    g078(.A(G106gat), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n278_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(KEYINPUT71), .A2(KEYINPUT7), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT72), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n282_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n285_));
  NOR2_X1   g084(.A1(G99gat), .A2(G106gat), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n278_), .A4(new_n286_), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n283_), .A2(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n259_), .A2(new_n261_), .A3(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n245_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT8), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n292_), .A2(KEYINPUT73), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n293_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n283_), .A2(new_n287_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n296_), .A2(new_n261_), .A3(new_n259_), .A4(new_n289_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n295_), .B1(new_n297_), .B2(new_n245_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n277_), .B1(new_n294_), .B2(new_n298_), .ZN(new_n299_));
  OR2_X1    g098(.A1(KEYINPUT74), .A2(G71gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(KEYINPUT74), .A2(G71gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(G78gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n300_), .A2(G78gat), .A3(new_n301_), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(G57gat), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n307_), .A2(G64gat), .ZN(new_n308_));
  INV_X1    g107(.A(G64gat), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n309_), .A2(G57gat), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT75), .B1(new_n308_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT11), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(G57gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n307_), .A2(G64gat), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT75), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n311_), .A2(new_n312_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n306_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT76), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n311_), .A2(new_n316_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n319_), .B1(new_n320_), .B2(KEYINPUT11), .ZN(new_n321_));
  AOI211_X1 g120(.A(KEYINPUT76), .B(new_n312_), .C1(new_n311_), .C2(new_n316_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n318_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  AND3_X1   g122(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n315_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT11), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT76), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n320_), .A2(new_n319_), .A3(KEYINPUT11), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n327_), .A2(new_n328_), .A3(new_n317_), .A4(new_n306_), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n323_), .A2(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n299_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G230gat), .A2(G233gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT64), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n299_), .A2(new_n330_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT78), .ZN(new_n336_));
  AOI21_X1  g135(.A(KEYINPUT12), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT12), .ZN(new_n338_));
  AOI211_X1 g137(.A(KEYINPUT78), .B(new_n338_), .C1(new_n299_), .C2(new_n330_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n334_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT77), .B1(new_n299_), .B2(new_n330_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n291_), .A2(new_n293_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n297_), .A2(new_n295_), .A3(new_n245_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n323_), .A2(new_n329_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .A4(new_n277_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n341_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n335_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n333_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n340_), .A2(new_n350_), .ZN(new_n351_));
  XOR2_X1   g150(.A(G120gat), .B(G148gat), .Z(new_n352_));
  XNOR2_X1  g151(.A(G176gat), .B(G204gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n351_), .A2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n351_), .A2(new_n357_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n241_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n351_), .A2(new_n357_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n351_), .A2(new_n357_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n361_), .A2(KEYINPUT13), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n360_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT80), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n360_), .A2(new_n363_), .A3(KEYINPUT80), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n240_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G231gat), .A2(G233gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n213_), .B(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(new_n345_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT17), .ZN(new_n372_));
  XOR2_X1   g171(.A(G127gat), .B(G155gat), .Z(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT16), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G183gat), .B(G211gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  OR3_X1    g175(.A1(new_n371_), .A2(new_n372_), .A3(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(KEYINPUT17), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n371_), .A2(new_n378_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n368_), .A2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(G176gat), .B1(KEYINPUT91), .B2(KEYINPUT22), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(G169gat), .ZN(new_n383_));
  INV_X1    g182(.A(G183gat), .ZN(new_n384_));
  INV_X1    g183(.A(G190gat), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n384_), .A2(new_n385_), .A3(KEYINPUT23), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT23), .B1(new_n384_), .B2(new_n385_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(G183gat), .A2(G190gat), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n383_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n388_), .B(KEYINPUT90), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n392_), .A2(new_n386_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT26), .B(G190gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT25), .B(G183gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(G169gat), .A2(G176gat), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT24), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  AND2_X1   g198(.A1(G169gat), .A2(G176gat), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n400_), .A2(new_n397_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n396_), .B(new_n399_), .C1(new_n398_), .C2(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n391_), .B1(new_n393_), .B2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G71gat), .B(G99gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(G43gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n403_), .B(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(G113gat), .B(G120gat), .Z(new_n407_));
  XNOR2_X1  g206(.A(G127gat), .B(G134gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n406_), .B(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G227gat), .A2(G233gat), .ZN(new_n411_));
  INV_X1    g210(.A(G15gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT30), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT31), .ZN(new_n415_));
  XOR2_X1   g214(.A(new_n410_), .B(new_n415_), .Z(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT97), .B(G204gat), .ZN(new_n417_));
  MUX2_X1   g216(.A(G204gat), .B(new_n417_), .S(G197gat), .Z(new_n418_));
  XNOR2_X1  g217(.A(G211gat), .B(G218gat), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT21), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n418_), .A2(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n418_), .A2(KEYINPUT21), .ZN(new_n423_));
  INV_X1    g222(.A(G197gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n417_), .A2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n420_), .B1(G197gat), .B2(G204gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n419_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n422_), .B1(new_n423_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT102), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n431_), .B1(new_n393_), .B2(new_n390_), .ZN(new_n432_));
  OAI221_X1 g231(.A(KEYINPUT102), .B1(G183gat), .B2(G190gat), .C1(new_n392_), .C2(new_n386_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT22), .B(G169gat), .ZN(new_n434_));
  INV_X1    g233(.A(G176gat), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n400_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n432_), .A2(new_n433_), .A3(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT101), .B(KEYINPUT24), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n387_), .A2(new_n388_), .B1(new_n438_), .B2(new_n397_), .ZN(new_n439_));
  XOR2_X1   g238(.A(new_n395_), .B(KEYINPUT100), .Z(new_n440_));
  INV_X1    g239(.A(new_n394_), .ZN(new_n441_));
  OAI221_X1 g240(.A(new_n439_), .B1(new_n401_), .B2(new_n438_), .C1(new_n440_), .C2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n430_), .B1(new_n437_), .B2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT20), .B1(new_n403_), .B2(new_n429_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G226gat), .A2(G233gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT19), .ZN(new_n447_));
  XOR2_X1   g246(.A(new_n447_), .B(KEYINPUT99), .Z(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n437_), .A2(new_n430_), .A3(new_n442_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT20), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n451_), .B1(new_n403_), .B2(new_n429_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n445_), .A2(new_n449_), .B1(new_n453_), .B2(new_n447_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n448_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n447_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n450_), .A2(new_n456_), .A3(new_n452_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G8gat), .B(G36gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT18), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G64gat), .B(G92gat), .ZN(new_n461_));
  XOR2_X1   g260(.A(new_n460_), .B(new_n461_), .Z(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT32), .ZN(new_n463_));
  MUX2_X1   g262(.A(new_n454_), .B(new_n458_), .S(new_n463_), .Z(new_n464_));
  XNOR2_X1  g263(.A(G1gat), .B(G29gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(G85gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT0), .B(G57gat), .ZN(new_n467_));
  XOR2_X1   g266(.A(new_n466_), .B(new_n467_), .Z(new_n468_));
  NOR2_X1   g267(.A1(G141gat), .A2(G148gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT3), .ZN(new_n470_));
  INV_X1    g269(.A(G141gat), .ZN(new_n471_));
  INV_X1    g270(.A(G148gat), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT93), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT2), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT2), .ZN(new_n476_));
  OAI211_X1 g275(.A(KEYINPUT93), .B(new_n476_), .C1(new_n471_), .C2(new_n472_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n470_), .A2(new_n475_), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT94), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G155gat), .A2(G162gat), .ZN(new_n481_));
  NOR2_X1   g280(.A1(G155gat), .A2(G162gat), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n480_), .A2(new_n481_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n409_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n481_), .B1(new_n482_), .B2(KEYINPUT1), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT92), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n488_), .B1(KEYINPUT1), .B2(new_n481_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n486_), .A2(new_n487_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  OR3_X1    g290(.A1(new_n491_), .A2(new_n469_), .A3(new_n473_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n484_), .A2(new_n485_), .A3(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n483_), .A2(new_n481_), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n478_), .A2(new_n479_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n478_), .A2(new_n479_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n494_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NOR3_X1   g296(.A1(new_n491_), .A2(new_n469_), .A3(new_n473_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n409_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n493_), .A2(KEYINPUT4), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G225gat), .A2(G233gat), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT4), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n503_), .B(new_n409_), .C1(new_n497_), .C2(new_n498_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n500_), .A2(new_n502_), .A3(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n493_), .A2(new_n501_), .A3(new_n499_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n468_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n507_), .A2(KEYINPUT103), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n505_), .A2(new_n468_), .A3(new_n506_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n509_), .B1(new_n507_), .B2(KEYINPUT103), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n464_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n462_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n458_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n455_), .A2(new_n457_), .A3(new_n462_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n505_), .A2(new_n506_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(KEYINPUT33), .A3(new_n468_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT33), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n509_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n500_), .A2(new_n501_), .A3(new_n504_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n468_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n493_), .A2(new_n502_), .A3(new_n499_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n516_), .A2(new_n518_), .A3(new_n520_), .A4(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n511_), .A2(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(KEYINPUT29), .B1(new_n497_), .B2(new_n498_), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n527_), .A2(new_n303_), .A3(new_n429_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n303_), .B1(new_n527_), .B2(new_n429_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n280_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n429_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(G78gat), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n527_), .A2(new_n303_), .A3(new_n429_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(G106gat), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(G233gat), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n535_), .A2(KEYINPUT96), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(KEYINPUT96), .ZN(new_n537_));
  OAI21_X1  g336(.A(G228gat), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT98), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n538_), .B1(new_n429_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n530_), .A2(new_n534_), .A3(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n541_), .B1(new_n530_), .B2(new_n534_), .ZN(new_n543_));
  XOR2_X1   g342(.A(G22gat), .B(G50gat), .Z(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  XOR2_X1   g344(.A(KEYINPUT95), .B(KEYINPUT28), .Z(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n497_), .A2(new_n498_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT29), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n547_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n548_), .A2(new_n549_), .A3(new_n547_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n545_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  AND3_X1   g352(.A1(new_n551_), .A2(new_n545_), .A3(new_n552_), .ZN(new_n554_));
  OAI22_X1  g353(.A1(new_n542_), .A2(new_n543_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n530_), .A2(new_n534_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(new_n540_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n554_), .A2(new_n553_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n530_), .A2(new_n534_), .A3(new_n541_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n557_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n555_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n526_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n555_), .A2(new_n560_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT104), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n564_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n507_), .A2(KEYINPUT103), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n507_), .A2(KEYINPUT103), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n566_), .A2(KEYINPUT104), .A3(new_n509_), .A4(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT27), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n514_), .A2(KEYINPUT27), .ZN(new_n570_));
  NOR3_X1   g369(.A1(new_n443_), .A2(new_n448_), .A3(new_n444_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n456_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n512_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n569_), .A2(new_n515_), .B1(new_n570_), .B2(new_n573_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n563_), .A2(new_n565_), .A3(new_n568_), .A4(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n416_), .B1(new_n562_), .B2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n565_), .A2(new_n568_), .A3(new_n416_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n574_), .A2(new_n555_), .A3(new_n560_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT105), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT105), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n574_), .A2(new_n555_), .A3(new_n560_), .A4(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n577_), .B1(new_n579_), .B2(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n576_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT34), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n585_), .A2(KEYINPUT35), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(KEYINPUT35), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n277_), .B(new_n215_), .C1(new_n294_), .C2(new_n298_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n207_), .B1(new_n344_), .B2(new_n277_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n588_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT83), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n207_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n299_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n596_), .A2(new_n589_), .A3(new_n586_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n589_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n598_), .A2(KEYINPUT83), .A3(new_n588_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G190gat), .B(G218gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT81), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G134gat), .B(G162gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT36), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n605_), .B(KEYINPUT82), .Z(new_n606_));
  NAND4_X1  g405(.A1(new_n594_), .A2(new_n597_), .A3(new_n599_), .A4(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT84), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n603_), .B(KEYINPUT36), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n597_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n610_));
  AOI21_X1  g409(.A(KEYINPUT83), .B1(new_n598_), .B2(new_n588_), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n608_), .B(new_n609_), .C1(new_n610_), .C2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n594_), .A2(new_n597_), .A3(new_n599_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n608_), .B1(new_n614_), .B2(new_n609_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n607_), .B1(new_n613_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(KEYINPUT107), .B1(new_n583_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT107), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n619_), .B(new_n616_), .C1(new_n576_), .C2(new_n582_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n381_), .B1(new_n618_), .B2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n565_), .A2(new_n568_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n202_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n562_), .A2(new_n575_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n416_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n579_), .A2(new_n581_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n622_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(new_n628_), .A3(new_n416_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n626_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n614_), .A2(new_n609_), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n631_), .A2(KEYINPUT37), .A3(new_n607_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT37), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n632_), .B1(new_n616_), .B2(new_n633_), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n380_), .B(KEYINPUT85), .Z(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n630_), .A2(new_n637_), .A3(new_n368_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT106), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT106), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n630_), .A2(new_n368_), .A3(new_n640_), .A4(new_n637_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n639_), .A2(new_n202_), .A3(new_n622_), .A4(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n623_), .B1(new_n643_), .B2(KEYINPUT38), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n643_), .A2(KEYINPUT108), .A3(KEYINPUT38), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT108), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT38), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n646_), .B1(new_n642_), .B2(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n644_), .B1(new_n645_), .B2(new_n648_), .ZN(G1324gat));
  INV_X1    g448(.A(KEYINPUT40), .ZN(new_n650_));
  INV_X1    g449(.A(new_n574_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n639_), .A2(new_n209_), .A3(new_n651_), .A4(new_n641_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT109), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  AOI211_X1 g453(.A(new_n574_), .B(new_n381_), .C1(new_n618_), .C2(new_n620_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n654_), .B1(new_n655_), .B2(new_n209_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n621_), .A2(new_n651_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(KEYINPUT39), .A3(G8gat), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n650_), .B1(new_n653_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT109), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n652_), .B(new_n661_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n662_), .A2(KEYINPUT40), .A3(new_n658_), .A4(new_n656_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n660_), .A2(new_n663_), .ZN(G1325gat));
  NAND2_X1  g463(.A1(new_n621_), .A2(new_n416_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(G15gat), .ZN(new_n666_));
  XOR2_X1   g465(.A(KEYINPUT110), .B(KEYINPUT41), .Z(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n638_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n670_), .A2(new_n412_), .A3(new_n416_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n665_), .A2(G15gat), .A3(new_n667_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n669_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT111), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n669_), .A2(KEYINPUT111), .A3(new_n671_), .A4(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1326gat));
  INV_X1    g476(.A(G22gat), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n670_), .A2(new_n678_), .A3(new_n563_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT42), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n621_), .A2(new_n563_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n681_), .B2(G22gat), .ZN(new_n682_));
  AOI211_X1 g481(.A(KEYINPUT42), .B(new_n678_), .C1(new_n621_), .C2(new_n563_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n679_), .B1(new_n682_), .B2(new_n683_), .ZN(G1327gat));
  NOR2_X1   g483(.A1(new_n635_), .A2(new_n616_), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n630_), .A2(new_n368_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(G29gat), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n686_), .A2(new_n687_), .A3(new_n622_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n634_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n689_), .B1(new_n576_), .B2(new_n582_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n691_), .B1(new_n689_), .B2(KEYINPUT112), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n635_), .B1(new_n690_), .B2(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n630_), .A2(new_n689_), .A3(new_n692_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n694_), .A2(new_n368_), .A3(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n694_), .A2(new_n695_), .A3(KEYINPUT44), .A4(new_n368_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n698_), .A2(new_n622_), .A3(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT113), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G29gat), .B1(new_n700_), .B2(new_n701_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n688_), .B1(new_n702_), .B2(new_n703_), .ZN(G1328gat));
  NAND3_X1  g503(.A1(new_n698_), .A2(new_n651_), .A3(new_n699_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(G36gat), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n574_), .A2(G36gat), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n686_), .A2(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT45), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n706_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT46), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n706_), .A2(KEYINPUT46), .A3(new_n709_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1329gat));
  NAND3_X1  g513(.A1(new_n698_), .A2(new_n416_), .A3(new_n699_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(G43gat), .ZN(new_n716_));
  INV_X1    g515(.A(G43gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n686_), .A2(new_n717_), .A3(new_n416_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(KEYINPUT114), .B(KEYINPUT47), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n716_), .A2(new_n718_), .A3(new_n720_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1330gat));
  INV_X1    g523(.A(G50gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n686_), .A2(new_n725_), .A3(new_n563_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n698_), .A2(new_n563_), .A3(new_n699_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT115), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n727_), .A2(new_n728_), .A3(G50gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n727_), .B2(G50gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n726_), .B1(new_n729_), .B2(new_n730_), .ZN(G1331gat));
  NAND2_X1  g530(.A1(new_n366_), .A2(new_n367_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n240_), .ZN(new_n733_));
  NOR4_X1   g532(.A1(new_n583_), .A2(new_n636_), .A3(new_n732_), .A4(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(new_n307_), .A3(new_n622_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n732_), .A2(new_n733_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(new_n635_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n620_), .B2(new_n618_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(new_n622_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n739_), .B2(new_n307_), .ZN(G1332gat));
  NAND3_X1  g539(.A1(new_n734_), .A2(new_n309_), .A3(new_n651_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT48), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n738_), .A2(new_n651_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n743_), .B2(G64gat), .ZN(new_n744_));
  AOI211_X1 g543(.A(KEYINPUT48), .B(new_n309_), .C1(new_n738_), .C2(new_n651_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n741_), .B1(new_n744_), .B2(new_n745_), .ZN(G1333gat));
  INV_X1    g545(.A(G71gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n734_), .A2(new_n747_), .A3(new_n416_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n738_), .A2(new_n416_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(KEYINPUT116), .B(KEYINPUT49), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n749_), .A2(G71gat), .A3(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n749_), .B2(G71gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(G1334gat));
  NAND3_X1  g552(.A1(new_n734_), .A2(new_n303_), .A3(new_n563_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n738_), .A2(new_n563_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(G78gat), .ZN(new_n757_));
  AOI211_X1 g556(.A(KEYINPUT50), .B(new_n303_), .C1(new_n738_), .C2(new_n563_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(G1335gat));
  NAND3_X1  g558(.A1(new_n694_), .A2(new_n695_), .A3(new_n736_), .ZN(new_n760_));
  OAI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n628_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n583_), .A2(new_n733_), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n732_), .A2(new_n635_), .A3(new_n616_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(G85gat), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n764_), .A2(new_n765_), .A3(new_n622_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n761_), .A2(new_n766_), .ZN(G1336gat));
  OAI21_X1  g566(.A(G92gat), .B1(new_n760_), .B2(new_n574_), .ZN(new_n768_));
  INV_X1    g567(.A(G92gat), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n764_), .A2(new_n769_), .A3(new_n651_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(G1337gat));
  OAI21_X1  g570(.A(G99gat), .B1(new_n760_), .B2(new_n625_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n764_), .B(new_n416_), .C1(new_n269_), .C2(new_n271_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g574(.A1(new_n694_), .A2(new_n695_), .A3(new_n563_), .A4(new_n736_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(G106gat), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n561_), .A2(new_n263_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n762_), .A2(new_n763_), .A3(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n781_), .B(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n776_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n779_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g585(.A1(new_n360_), .A2(new_n363_), .A3(new_n240_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n637_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n789_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(new_n636_), .B2(new_n787_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n238_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n233_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n231_), .A2(new_n221_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n214_), .A2(new_n220_), .A3(new_n232_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n238_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n795_), .A2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n799_), .B1(new_n351_), .B2(new_n357_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n337_), .A2(new_n339_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n333_), .B1(new_n801_), .B2(new_n348_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n340_), .A2(new_n803_), .ZN(new_n804_));
  OAI211_X1 g603(.A(KEYINPUT55), .B(new_n334_), .C1(new_n337_), .C2(new_n339_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n802_), .A2(new_n804_), .A3(new_n805_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n806_), .A2(KEYINPUT56), .A3(new_n356_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT56), .B1(new_n806_), .B2(new_n356_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n800_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT58), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n634_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n806_), .A2(new_n356_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT56), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n806_), .A2(KEYINPUT56), .A3(new_n356_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n816_), .A2(KEYINPUT119), .A3(KEYINPUT58), .A4(new_n800_), .ZN(new_n817_));
  OAI211_X1 g616(.A(KEYINPUT58), .B(new_n800_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT119), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n811_), .A2(new_n817_), .A3(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n358_), .A2(new_n240_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n824_));
  OAI22_X1  g623(.A1(new_n358_), .A2(new_n359_), .B1(new_n798_), .B2(new_n795_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n822_), .B1(new_n826_), .B2(new_n616_), .ZN(new_n827_));
  AOI211_X1 g626(.A(KEYINPUT57), .B(new_n617_), .C1(new_n824_), .C2(new_n825_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n821_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n635_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n793_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n627_), .A2(new_n622_), .A3(new_n416_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n833_), .A2(KEYINPUT59), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n380_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n793_), .B1(new_n829_), .B2(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n837_), .A2(new_n833_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT59), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n835_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(G113gat), .B1(new_n840_), .B2(new_n240_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n838_), .ZN(new_n842_));
  OR2_X1    g641(.A1(new_n240_), .A2(G113gat), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n841_), .B1(new_n842_), .B2(new_n843_), .ZN(G1340gat));
  OAI21_X1  g643(.A(G120gat), .B1(new_n840_), .B2(new_n732_), .ZN(new_n845_));
  INV_X1    g644(.A(G120gat), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(new_n732_), .B2(KEYINPUT60), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(KEYINPUT60), .B2(new_n846_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n845_), .B1(new_n842_), .B2(new_n848_), .ZN(G1341gat));
  OAI21_X1  g648(.A(G127gat), .B1(new_n840_), .B2(new_n836_), .ZN(new_n850_));
  OR2_X1    g649(.A1(new_n830_), .A2(G127gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n842_), .B2(new_n851_), .ZN(G1342gat));
  INV_X1    g651(.A(G134gat), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(new_n842_), .B2(new_n616_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(KEYINPUT120), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n856_), .B(new_n853_), .C1(new_n842_), .C2(new_n616_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n840_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n634_), .A2(new_n853_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(KEYINPUT121), .ZN(new_n860_));
  AOI22_X1  g659(.A1(new_n855_), .A2(new_n857_), .B1(new_n858_), .B2(new_n860_), .ZN(G1343gat));
  INV_X1    g660(.A(new_n837_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n622_), .A2(new_n563_), .A3(new_n574_), .A4(new_n625_), .ZN(new_n863_));
  XOR2_X1   g662(.A(new_n863_), .B(KEYINPUT122), .Z(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n865_), .A2(new_n240_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(new_n471_), .ZN(G1344gat));
  NOR2_X1   g666(.A1(new_n865_), .A2(new_n732_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(new_n472_), .ZN(G1345gat));
  NOR2_X1   g668(.A1(new_n865_), .A2(new_n830_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(KEYINPUT61), .B(G155gat), .ZN(new_n871_));
  XOR2_X1   g670(.A(new_n870_), .B(new_n871_), .Z(G1346gat));
  OAI21_X1  g671(.A(G162gat), .B1(new_n865_), .B2(new_n634_), .ZN(new_n873_));
  OR2_X1    g672(.A1(new_n616_), .A2(G162gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n865_), .B2(new_n874_), .ZN(G1347gat));
  INV_X1    g674(.A(KEYINPUT62), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n577_), .A2(new_n574_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n561_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n733_), .A2(new_n362_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n880_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n825_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n616_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(KEYINPUT57), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n826_), .A2(new_n822_), .A3(new_n616_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n635_), .B1(new_n886_), .B2(new_n821_), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n733_), .B(new_n879_), .C1(new_n887_), .C2(new_n793_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT123), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n888_), .A2(new_n889_), .A3(G169gat), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n889_), .B1(new_n888_), .B2(G169gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n876_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n892_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n894_), .A2(KEYINPUT62), .A3(new_n890_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT124), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n896_), .B1(new_n831_), .B2(new_n878_), .ZN(new_n897_));
  OAI211_X1 g696(.A(KEYINPUT124), .B(new_n879_), .C1(new_n887_), .C2(new_n793_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n733_), .A2(new_n434_), .ZN(new_n900_));
  XOR2_X1   g699(.A(new_n900_), .B(KEYINPUT125), .Z(new_n901_));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n901_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n893_), .A2(new_n895_), .A3(new_n902_), .ZN(G1348gat));
  INV_X1    g702(.A(new_n732_), .ZN(new_n904_));
  AOI21_X1  g703(.A(G176gat), .B1(new_n899_), .B2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n862_), .A2(new_n561_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n904_), .A2(G176gat), .A3(new_n877_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(KEYINPUT126), .B1(new_n905_), .B2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT126), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n732_), .B1(new_n897_), .B2(new_n898_), .ZN(new_n911_));
  OAI221_X1 g710(.A(new_n910_), .B1(new_n906_), .B2(new_n907_), .C1(new_n911_), .C2(G176gat), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n909_), .A2(new_n912_), .ZN(G1349gat));
  AND2_X1   g712(.A1(new_n380_), .A2(new_n440_), .ZN(new_n914_));
  NAND4_X1  g713(.A1(new_n862_), .A2(new_n635_), .A3(new_n561_), .A4(new_n877_), .ZN(new_n915_));
  AOI22_X1  g714(.A1(new_n899_), .A2(new_n914_), .B1(new_n915_), .B2(new_n384_), .ZN(G1350gat));
  NAND3_X1  g715(.A1(new_n899_), .A2(new_n617_), .A3(new_n394_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n634_), .B1(new_n897_), .B2(new_n898_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n918_), .B2(new_n385_), .ZN(G1351gat));
  NAND4_X1  g718(.A1(new_n628_), .A2(new_n563_), .A3(new_n651_), .A4(new_n625_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n837_), .A2(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n733_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n904_), .ZN(new_n924_));
  MUX2_X1   g723(.A(new_n417_), .B(G204gat), .S(new_n924_), .Z(G1353gat));
  NOR3_X1   g724(.A1(new_n837_), .A2(new_n836_), .A3(new_n920_), .ZN(new_n926_));
  NOR3_X1   g725(.A1(new_n926_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n927_));
  XOR2_X1   g726(.A(KEYINPUT63), .B(G211gat), .Z(new_n928_));
  AOI21_X1  g727(.A(new_n927_), .B1(new_n926_), .B2(new_n928_), .ZN(G1354gat));
  INV_X1    g728(.A(G218gat), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n921_), .A2(new_n930_), .A3(new_n617_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n837_), .A2(new_n634_), .A3(new_n920_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n930_), .B2(new_n932_), .ZN(G1355gat));
endmodule


