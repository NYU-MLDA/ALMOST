//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 0 1 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n606_, new_n607_, new_n608_, new_n609_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n802_, new_n803_, new_n804_, new_n805_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n817_, new_n818_, new_n819_, new_n821_, new_n822_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n861_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_;
  OR3_X1    g000(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n202_));
  OAI21_X1  g001(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G183gat), .A2(G190gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  OR2_X1    g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n204_), .B1(new_n210_), .B2(KEYINPUT75), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n210_), .A2(KEYINPUT75), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT24), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT74), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT74), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n216_), .A2(new_n219_), .A3(new_n207_), .A4(new_n209_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n214_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(KEYINPUT24), .A3(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT25), .B(G183gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT26), .B(G190gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n218_), .A2(new_n220_), .A3(new_n223_), .A4(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n213_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G71gat), .B(G99gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(G43gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n228_), .B(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(G127gat), .B(G134gat), .Z(new_n232_));
  XOR2_X1   g031(.A(G113gat), .B(G120gat), .Z(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n231_), .B(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G227gat), .A2(G233gat), .ZN(new_n237_));
  INV_X1    g036(.A(G15gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT30), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT31), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n236_), .B(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT77), .ZN(new_n243_));
  INV_X1    g042(.A(G155gat), .ZN(new_n244_));
  INV_X1    g043(.A(G162gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G155gat), .A2(G162gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT1), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT1), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(G155gat), .A3(G162gat), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT77), .B1(G155gat), .B2(G162gat), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n246_), .A2(new_n248_), .A3(new_n250_), .A4(new_n251_), .ZN(new_n252_));
  AND2_X1   g051(.A1(G141gat), .A2(G148gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT76), .ZN(new_n254_));
  INV_X1    g053(.A(G141gat), .ZN(new_n255_));
  INV_X1    g054(.A(G148gat), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n254_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT76), .B1(G141gat), .B2(G148gat), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n253_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n252_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT78), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT78), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n252_), .A2(new_n259_), .A3(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT79), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT79), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n266_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT2), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n269_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n253_), .A2(KEYINPUT2), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT3), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n272_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n268_), .A2(new_n270_), .A3(new_n271_), .A4(new_n273_), .ZN(new_n274_));
  AND3_X1   g073(.A1(new_n246_), .A2(new_n251_), .A3(new_n247_), .ZN(new_n275_));
  AOI22_X1  g074(.A1(new_n261_), .A2(new_n263_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT28), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT29), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n276_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n265_), .A2(new_n267_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n271_), .A2(new_n270_), .A3(new_n273_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n275_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n252_), .A2(new_n259_), .A3(new_n262_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n262_), .B1(new_n252_), .B2(new_n259_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n282_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT28), .B1(new_n285_), .B2(KEYINPUT29), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G22gat), .B(G50gat), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n279_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n287_), .B1(new_n279_), .B2(new_n286_), .ZN(new_n290_));
  OR3_X1    g089(.A1(new_n289_), .A2(KEYINPUT80), .A3(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(G211gat), .B(G218gat), .Z(new_n292_));
  INV_X1    g091(.A(G197gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(G204gat), .ZN(new_n294_));
  INV_X1    g093(.A(G204gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G197gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT21), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n292_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT81), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(new_n293_), .A3(G204gat), .ZN(new_n302_));
  OAI211_X1 g101(.A(KEYINPUT21), .B(new_n302_), .C1(new_n297_), .C2(new_n301_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n300_), .A2(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n298_), .A2(new_n299_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n292_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n307_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n308_));
  INV_X1    g107(.A(G228gat), .ZN(new_n309_));
  INV_X1    g108(.A(G233gat), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  OAI221_X1 g111(.A(new_n307_), .B1(new_n309_), .B2(new_n310_), .C1(new_n276_), .C2(new_n278_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G78gat), .B(G106gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n315_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n312_), .A2(new_n313_), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT80), .B1(new_n289_), .B2(new_n290_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n291_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT82), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n318_), .A2(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n289_), .A2(new_n290_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n312_), .A2(new_n313_), .A3(KEYINPUT82), .A4(new_n317_), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n323_), .A2(new_n324_), .A3(new_n316_), .A4(new_n325_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n321_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT98), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n285_), .A2(new_n235_), .ZN(new_n330_));
  OAI211_X1 g129(.A(new_n234_), .B(new_n282_), .C1(new_n284_), .C2(new_n283_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G225gat), .A2(G233gat), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n330_), .A2(KEYINPUT4), .A3(new_n331_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT4), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n285_), .A2(new_n336_), .A3(new_n235_), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n332_), .B(KEYINPUT90), .Z(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT91), .B1(new_n335_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n338_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n261_), .A2(new_n263_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n234_), .B1(new_n342_), .B2(new_n282_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n341_), .B1(new_n343_), .B2(new_n336_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT91), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n330_), .A2(KEYINPUT4), .A3(new_n331_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n334_), .B1(new_n340_), .B2(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G57gat), .B(G85gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT93), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(G1gat), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n349_), .A2(KEYINPUT93), .ZN(new_n352_));
  INV_X1    g151(.A(G1gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n349_), .A2(KEYINPUT93), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n351_), .A2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT92), .B(KEYINPUT0), .ZN(new_n357_));
  INV_X1    g156(.A(G29gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n356_), .B(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n329_), .B1(new_n348_), .B2(new_n360_), .ZN(new_n361_));
  NOR3_X1   g160(.A1(new_n335_), .A2(KEYINPUT91), .A3(new_n339_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n345_), .B1(new_n344_), .B2(new_n346_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n333_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n360_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n364_), .A2(KEYINPUT98), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n340_), .A2(new_n347_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n360_), .A2(new_n333_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT97), .B1(new_n367_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT97), .ZN(new_n371_));
  AOI211_X1 g170(.A(new_n371_), .B(new_n368_), .C1(new_n340_), .C2(new_n347_), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n361_), .B(new_n366_), .C1(new_n370_), .C2(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT20), .B1(new_n228_), .B2(new_n307_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT84), .B(KEYINPUT24), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(new_n222_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT85), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n375_), .A2(KEYINPUT85), .A3(new_n222_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n378_), .A2(new_n221_), .A3(new_n379_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n207_), .A2(new_n209_), .ZN(new_n381_));
  OR2_X1    g180(.A1(KEYINPUT84), .A2(KEYINPUT24), .ZN(new_n382_));
  NAND2_X1  g181(.A1(KEYINPUT84), .A2(KEYINPUT24), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(new_n214_), .A3(new_n383_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n226_), .A2(new_n381_), .A3(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n381_), .A2(KEYINPUT86), .A3(new_n208_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT86), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n204_), .B1(new_n210_), .B2(new_n387_), .ZN(new_n388_));
  AOI22_X1  g187(.A1(new_n380_), .A2(new_n385_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n300_), .A2(new_n303_), .B1(new_n305_), .B2(new_n292_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n392_));
  AND2_X1   g191(.A1(G226gat), .A2(G233gat), .ZN(new_n393_));
  XOR2_X1   g192(.A(new_n392_), .B(new_n393_), .Z(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NOR3_X1   g194(.A1(new_n374_), .A2(new_n391_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT20), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n397_), .B1(new_n228_), .B2(new_n307_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n389_), .A2(KEYINPUT96), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n390_), .B1(new_n389_), .B2(KEYINPUT96), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n398_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n396_), .B1(new_n402_), .B2(new_n395_), .ZN(new_n403_));
  AOI211_X1 g202(.A(new_n397_), .B(new_n395_), .C1(new_n228_), .C2(new_n307_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT87), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n389_), .A2(new_n405_), .A3(new_n390_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n405_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n404_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n395_), .B1(new_n374_), .B2(new_n391_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(KEYINPUT89), .ZN(new_n413_));
  XOR2_X1   g212(.A(G8gat), .B(G36gat), .Z(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G64gat), .B(G92gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT32), .ZN(new_n418_));
  MUX2_X1   g217(.A(new_n403_), .B(new_n411_), .S(new_n418_), .Z(new_n419_));
  NAND2_X1  g218(.A1(new_n373_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n417_), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n226_), .A2(new_n220_), .A3(new_n223_), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n422_), .A2(new_n218_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n423_));
  OAI211_X1 g222(.A(KEYINPUT20), .B(new_n394_), .C1(new_n423_), .C2(new_n390_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n380_), .A2(new_n385_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n388_), .A2(new_n386_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT87), .B1(new_n427_), .B2(new_n307_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n424_), .B1(new_n428_), .B2(new_n406_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n307_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n397_), .B1(new_n423_), .B2(new_n390_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n394_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n421_), .B1(new_n429_), .B2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n409_), .A2(new_n410_), .A3(new_n417_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n346_), .A2(new_n337_), .A3(new_n332_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n330_), .A2(new_n331_), .A3(new_n338_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n365_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT95), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT95), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n365_), .A2(new_n436_), .A3(new_n440_), .A4(new_n437_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n435_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n369_), .B(KEYINPUT33), .C1(new_n362_), .C2(new_n363_), .ZN(new_n443_));
  OR2_X1    g242(.A1(new_n443_), .A2(KEYINPUT94), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(KEYINPUT94), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n369_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT33), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n442_), .A2(new_n444_), .A3(new_n445_), .A4(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n328_), .B1(new_n420_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT27), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n435_), .A2(new_n451_), .ZN(new_n452_));
  OAI211_X1 g251(.A(KEYINPUT27), .B(new_n434_), .C1(new_n403_), .C2(new_n417_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NOR3_X1   g253(.A1(new_n373_), .A2(new_n327_), .A3(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n242_), .B1(new_n450_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT99), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n452_), .A2(new_n453_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n327_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT100), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n458_), .A2(KEYINPUT100), .A3(new_n327_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n373_), .A2(new_n242_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT99), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n466_), .B(new_n242_), .C1(new_n450_), .C2(new_n455_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n457_), .A2(new_n465_), .A3(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(G29gat), .B(G36gat), .Z(new_n469_));
  XOR2_X1   g268(.A(G43gat), .B(G50gat), .Z(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G29gat), .B(G36gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G43gat), .B(G50gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n471_), .A2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT15), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G15gat), .B(G22gat), .ZN(new_n477_));
  INV_X1    g276(.A(G8gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT14), .B1(new_n353_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G1gat), .B(G8gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n476_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n475_), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G229gat), .A2(G233gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n482_), .B(new_n484_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n489_), .A2(G229gat), .A3(G233gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G113gat), .B(G141gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G169gat), .B(G197gat), .ZN(new_n493_));
  XOR2_X1   g292(.A(new_n492_), .B(new_n493_), .Z(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT70), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n491_), .A2(new_n495_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n496_), .A2(KEYINPUT71), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n488_), .A2(new_n490_), .A3(new_n494_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n498_), .B1(new_n496_), .B2(KEYINPUT71), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n500_), .A2(KEYINPUT72), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(KEYINPUT72), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT73), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n468_), .A2(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(G85gat), .B(G92gat), .Z(new_n506_));
  NOR2_X1   g305(.A1(G99gat), .A2(G106gat), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT7), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G99gat), .A2(G106gat), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT6), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n506_), .B1(new_n509_), .B2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT8), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT64), .B(G85gat), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(G92gat), .ZN(new_n517_));
  OR3_X1    g316(.A1(new_n516_), .A2(KEYINPUT9), .A3(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n512_), .B1(KEYINPUT9), .B2(new_n506_), .ZN(new_n519_));
  XOR2_X1   g318(.A(KEYINPUT10), .B(G99gat), .Z(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n518_), .B(new_n519_), .C1(G106gat), .C2(new_n521_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n514_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G57gat), .B(G64gat), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n524_), .A2(KEYINPUT11), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G71gat), .B(G78gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n525_), .A2(new_n526_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n524_), .A2(KEYINPUT11), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n527_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n523_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(G230gat), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n531_), .B1(new_n532_), .B2(new_n310_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT65), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n534_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n523_), .A2(new_n530_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT12), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n535_), .A2(new_n536_), .A3(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n531_), .ZN(new_n541_));
  OAI211_X1 g340(.A(G230gat), .B(G233gat), .C1(new_n541_), .C2(new_n537_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(KEYINPUT66), .B(KEYINPUT5), .Z(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT67), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G120gat), .B(G148gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G176gat), .B(G204gat), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n547_), .B(new_n548_), .Z(new_n549_));
  OR2_X1    g348(.A1(new_n543_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n543_), .A2(new_n549_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT13), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n550_), .A2(KEYINPUT13), .A3(new_n551_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n523_), .A2(new_n475_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G232gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT34), .ZN(new_n559_));
  INV_X1    g358(.A(new_n476_), .ZN(new_n560_));
  OAI221_X1 g359(.A(new_n557_), .B1(KEYINPUT35), .B2(new_n559_), .C1(new_n560_), .C2(new_n523_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(KEYINPUT35), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G190gat), .B(G218gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G134gat), .B(G162gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n566_), .A2(KEYINPUT36), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n563_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n566_), .B(KEYINPUT36), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n563_), .A2(new_n569_), .ZN(new_n570_));
  OR3_X1    g369(.A1(new_n568_), .A2(new_n570_), .A3(KEYINPUT37), .ZN(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT37), .B1(new_n568_), .B2(new_n570_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G231gat), .A2(G233gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n482_), .B(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n576_), .B(new_n530_), .Z(new_n577_));
  XNOR2_X1  g376(.A(G127gat), .B(G155gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G183gat), .B(G211gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT69), .B(KEYINPUT16), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT68), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT17), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n582_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n582_), .A2(new_n584_), .ZN(new_n586_));
  OR3_X1    g385(.A1(new_n577_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n577_), .A2(new_n585_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n574_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n505_), .A2(new_n556_), .A3(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n591_), .B(KEYINPUT101), .Z(new_n592_));
  NAND3_X1  g391(.A1(new_n592_), .A2(new_n353_), .A3(new_n373_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT38), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n556_), .A2(new_n503_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n596_), .A2(new_n589_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n568_), .A2(new_n570_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT102), .Z(new_n599_));
  AND2_X1   g398(.A1(new_n468_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n597_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n373_), .ZN(new_n602_));
  OAI21_X1  g401(.A(G1gat), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n593_), .A2(new_n594_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n595_), .A2(new_n603_), .A3(new_n604_), .ZN(G1324gat));
  NAND3_X1  g404(.A1(new_n592_), .A2(new_n478_), .A3(new_n454_), .ZN(new_n606_));
  OAI21_X1  g405(.A(G8gat), .B1(new_n601_), .B2(new_n458_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT39), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n609_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g409(.A(G15gat), .B1(new_n601_), .B2(new_n242_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT41), .Z(new_n612_));
  INV_X1    g411(.A(new_n242_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n592_), .A2(new_n238_), .A3(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(G1326gat));
  INV_X1    g414(.A(G22gat), .ZN(new_n616_));
  INV_X1    g415(.A(new_n601_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n327_), .B(KEYINPUT103), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n616_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n619_), .B(KEYINPUT42), .Z(new_n620_));
  NAND3_X1  g419(.A1(new_n592_), .A2(new_n616_), .A3(new_n618_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(G1327gat));
  NAND3_X1  g421(.A1(new_n556_), .A2(new_n503_), .A3(new_n589_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT104), .ZN(new_n625_));
  OAI21_X1  g424(.A(KEYINPUT43), .B1(new_n573_), .B2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n467_), .A2(new_n465_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n602_), .A2(new_n328_), .A3(new_n458_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n433_), .A2(new_n434_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n439_), .A2(new_n441_), .ZN(new_n630_));
  AND4_X1   g429(.A1(new_n445_), .A2(new_n629_), .A3(new_n448_), .A4(new_n630_), .ZN(new_n631_));
  AOI22_X1  g430(.A1(new_n631_), .A2(new_n444_), .B1(new_n373_), .B2(new_n419_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n628_), .B1(new_n632_), .B2(new_n328_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n466_), .B1(new_n633_), .B2(new_n242_), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n626_), .B(new_n574_), .C1(new_n627_), .C2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n626_), .B1(new_n468_), .B2(new_n574_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n624_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT106), .ZN(new_n639_));
  XNOR2_X1  g438(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n638_), .A2(new_n639_), .A3(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n574_), .B1(new_n627_), .B2(new_n634_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n626_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n623_), .B1(new_n645_), .B2(new_n635_), .ZN(new_n646_));
  OAI21_X1  g445(.A(KEYINPUT106), .B1(new_n646_), .B2(new_n640_), .ZN(new_n647_));
  AOI22_X1  g446(.A1(new_n642_), .A2(new_n647_), .B1(KEYINPUT44), .B2(new_n646_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n648_), .A2(new_n373_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n598_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n589_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n556_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n505_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n373_), .A2(new_n358_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT107), .ZN(new_n656_));
  OAI22_X1  g455(.A1(new_n649_), .A2(new_n358_), .B1(new_n654_), .B2(new_n656_), .ZN(G1328gat));
  INV_X1    g456(.A(new_n654_), .ZN(new_n658_));
  INV_X1    g457(.A(G36gat), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n658_), .A2(new_n659_), .A3(new_n454_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT45), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n642_), .A2(new_n647_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n458_), .B1(new_n646_), .B2(KEYINPUT44), .ZN(new_n663_));
  AOI211_X1 g462(.A(KEYINPUT108), .B(new_n659_), .C1(new_n662_), .C2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT108), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n639_), .B1(new_n638_), .B2(new_n641_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n646_), .A2(KEYINPUT106), .A3(new_n640_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n663_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n665_), .B1(new_n668_), .B2(G36gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n661_), .B1(new_n664_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT46), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OAI211_X1 g471(.A(KEYINPUT46), .B(new_n661_), .C1(new_n664_), .C2(new_n669_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1329gat));
  NAND3_X1  g473(.A1(new_n648_), .A2(G43gat), .A3(new_n613_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n654_), .A2(new_n242_), .ZN(new_n676_));
  XOR2_X1   g475(.A(KEYINPUT109), .B(G43gat), .Z(new_n677_));
  OAI21_X1  g476(.A(new_n675_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g478(.A(G50gat), .B1(new_n658_), .B2(new_n618_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n328_), .A2(G50gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n648_), .B2(new_n681_), .ZN(G1331gat));
  INV_X1    g481(.A(G57gat), .ZN(new_n683_));
  INV_X1    g482(.A(new_n503_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n556_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n468_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(new_n590_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n683_), .B1(new_n688_), .B2(new_n602_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n556_), .A2(new_n504_), .A3(new_n589_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n600_), .A2(new_n690_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n691_), .A2(new_n683_), .A3(new_n602_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n689_), .B1(new_n692_), .B2(KEYINPUT110), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n693_), .B1(KEYINPUT110), .B2(new_n692_), .ZN(G1332gat));
  OAI21_X1  g493(.A(G64gat), .B1(new_n691_), .B2(new_n458_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT48), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n458_), .A2(G64gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n696_), .B1(new_n688_), .B2(new_n697_), .ZN(G1333gat));
  OAI21_X1  g497(.A(G71gat), .B1(new_n691_), .B2(new_n242_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT49), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n242_), .A2(G71gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n700_), .B1(new_n688_), .B2(new_n701_), .ZN(G1334gat));
  INV_X1    g501(.A(G78gat), .ZN(new_n703_));
  INV_X1    g502(.A(new_n691_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n704_), .B2(new_n618_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT50), .Z(new_n706_));
  NAND2_X1  g505(.A1(new_n618_), .A2(new_n703_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT111), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n706_), .B1(new_n688_), .B2(new_n708_), .ZN(G1335gat));
  NAND2_X1  g508(.A1(new_n687_), .A2(new_n652_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(G85gat), .B1(new_n711_), .B2(new_n373_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT112), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n684_), .A2(new_n589_), .ZN(new_n714_));
  AOI211_X1 g513(.A(new_n556_), .B(new_n714_), .C1(new_n645_), .C2(new_n635_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n602_), .A2(new_n516_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n713_), .B1(new_n715_), .B2(new_n716_), .ZN(G1336gat));
  NAND3_X1  g516(.A1(new_n711_), .A2(new_n517_), .A3(new_n454_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n715_), .A2(new_n454_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n719_), .B2(new_n517_), .ZN(G1337gat));
  NOR2_X1   g519(.A1(new_n242_), .A2(new_n521_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT113), .B1(new_n711_), .B2(new_n721_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n715_), .A2(new_n613_), .ZN(new_n723_));
  INV_X1    g522(.A(G99gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n722_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g525(.A(G106gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n711_), .A2(new_n727_), .A3(new_n328_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT52), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n715_), .A2(new_n328_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n730_), .B2(G106gat), .ZN(new_n731_));
  AOI211_X1 g530(.A(KEYINPUT52), .B(new_n727_), .C1(new_n715_), .C2(new_n328_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI22_X1  g533(.A1(new_n501_), .A2(new_n502_), .B1(new_n543_), .B2(new_n549_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT55), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n540_), .A2(new_n736_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n535_), .A2(new_n539_), .A3(KEYINPUT55), .A4(new_n536_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n539_), .A2(new_n531_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n739_), .A2(G230gat), .A3(G233gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n737_), .A2(new_n738_), .A3(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n549_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT114), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(KEYINPUT56), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT56), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n741_), .A2(KEYINPUT114), .A3(new_n747_), .A4(new_n742_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n735_), .A2(new_n745_), .A3(new_n746_), .A4(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n498_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n486_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n487_), .B1(new_n751_), .B2(KEYINPUT115), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n752_), .B1(KEYINPUT115), .B2(new_n751_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n494_), .B1(new_n489_), .B2(new_n487_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n750_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n552_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n749_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n650_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT57), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n598_), .B1(new_n749_), .B2(new_n756_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT57), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n551_), .A2(new_n755_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n741_), .A2(new_n747_), .A3(new_n742_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n746_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT116), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT58), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n765_), .A2(new_n766_), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n767_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n746_), .A2(new_n763_), .A3(new_n764_), .A4(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n768_), .A2(new_n574_), .A3(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n760_), .A2(new_n762_), .A3(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n590_), .A2(new_n556_), .ZN(new_n773_));
  OAI21_X1  g572(.A(KEYINPUT54), .B1(new_n773_), .B2(new_n504_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n504_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT54), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n775_), .A2(new_n556_), .A3(new_n776_), .A4(new_n590_), .ZN(new_n777_));
  AOI22_X1  g576(.A1(new_n772_), .A2(new_n589_), .B1(new_n774_), .B2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n463_), .A2(new_n613_), .A3(new_n373_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(G113gat), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(new_n781_), .A3(new_n503_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT59), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT117), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(KEYINPUT117), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n784_), .B(new_n786_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n762_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n771_), .B1(new_n761_), .B2(KEYINPUT57), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n589_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n774_), .A2(new_n777_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT117), .ZN(new_n793_));
  INV_X1    g592(.A(new_n779_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n792_), .A2(new_n793_), .A3(KEYINPUT59), .A4(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n775_), .B1(new_n787_), .B2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n782_), .B1(new_n796_), .B2(new_n781_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT118), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT118), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n799_), .B(new_n782_), .C1(new_n796_), .C2(new_n781_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(G1340gat));
  INV_X1    g600(.A(G120gat), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n802_), .B1(new_n556_), .B2(KEYINPUT60), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n780_), .B(new_n803_), .C1(KEYINPUT60), .C2(new_n802_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n556_), .B1(new_n787_), .B2(new_n795_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(new_n802_), .ZN(G1341gat));
  AOI21_X1  g605(.A(G127gat), .B1(new_n780_), .B2(new_n651_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n787_), .A2(new_n795_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n651_), .A2(G127gat), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT119), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n807_), .B1(new_n808_), .B2(new_n810_), .ZN(G1342gat));
  INV_X1    g610(.A(G134gat), .ZN(new_n812_));
  INV_X1    g611(.A(new_n599_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n780_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n573_), .B1(new_n787_), .B2(new_n795_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n814_), .B1(new_n815_), .B2(new_n812_), .ZN(G1343gat));
  NOR3_X1   g615(.A1(new_n602_), .A2(new_n327_), .A3(new_n454_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n792_), .A2(new_n242_), .A3(new_n817_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n818_), .A2(new_n684_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(new_n255_), .ZN(G1344gat));
  NOR2_X1   g619(.A1(new_n818_), .A2(new_n556_), .ZN(new_n821_));
  XOR2_X1   g620(.A(KEYINPUT120), .B(G148gat), .Z(new_n822_));
  XNOR2_X1  g621(.A(new_n821_), .B(new_n822_), .ZN(G1345gat));
  INV_X1    g622(.A(new_n818_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n824_), .A2(KEYINPUT121), .A3(new_n651_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT121), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n818_), .B2(new_n589_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(KEYINPUT61), .B(G155gat), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n828_), .B(new_n829_), .ZN(G1346gat));
  OAI21_X1  g629(.A(G162gat), .B1(new_n818_), .B2(new_n573_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n813_), .A2(new_n245_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n818_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT122), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n833_), .B(new_n834_), .ZN(G1347gat));
  INV_X1    g634(.A(KEYINPUT124), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n602_), .A2(new_n454_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n837_), .A2(new_n242_), .ZN(new_n838_));
  XOR2_X1   g637(.A(new_n838_), .B(KEYINPUT123), .Z(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(new_n618_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n792_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n503_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT62), .ZN(new_n844_));
  AND4_X1   g643(.A1(new_n836_), .A2(new_n843_), .A3(new_n844_), .A4(G169gat), .ZN(new_n845_));
  INV_X1    g644(.A(G169gat), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n846_), .B1(KEYINPUT124), .B2(KEYINPUT62), .ZN(new_n847_));
  AOI22_X1  g646(.A1(new_n843_), .A2(new_n847_), .B1(new_n836_), .B2(new_n844_), .ZN(new_n848_));
  XOR2_X1   g647(.A(KEYINPUT22), .B(G169gat), .Z(new_n849_));
  OAI22_X1  g648(.A1(new_n845_), .A2(new_n848_), .B1(new_n843_), .B2(new_n849_), .ZN(G1348gat));
  AOI21_X1  g649(.A(G176gat), .B1(new_n842_), .B2(new_n685_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n778_), .A2(new_n328_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n839_), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n853_), .A2(G176gat), .A3(new_n685_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n851_), .B1(new_n852_), .B2(new_n854_), .ZN(G1349gat));
  NOR3_X1   g654(.A1(new_n841_), .A2(new_n224_), .A3(new_n589_), .ZN(new_n856_));
  INV_X1    g655(.A(G183gat), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n852_), .A2(new_n651_), .A3(new_n853_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n856_), .B1(new_n857_), .B2(new_n858_), .ZN(G1350gat));
  OAI21_X1  g658(.A(G190gat), .B1(new_n841_), .B2(new_n573_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n813_), .A2(new_n225_), .ZN(new_n861_));
  XOR2_X1   g660(.A(new_n861_), .B(KEYINPUT125), .Z(new_n862_));
  OAI21_X1  g661(.A(new_n860_), .B1(new_n841_), .B2(new_n862_), .ZN(G1351gat));
  NOR2_X1   g662(.A1(new_n837_), .A2(new_n327_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n792_), .A2(new_n242_), .A3(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT126), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n792_), .A2(KEYINPUT126), .A3(new_n242_), .A4(new_n864_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n503_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G197gat), .ZN(G1352gat));
  AOI21_X1  g670(.A(new_n556_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(KEYINPUT127), .B2(new_n295_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT127), .B(G204gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n872_), .B2(new_n874_), .ZN(G1353gat));
  XNOR2_X1  g674(.A(KEYINPUT63), .B(G211gat), .ZN(new_n876_));
  AOI211_X1 g675(.A(new_n589_), .B(new_n876_), .C1(new_n867_), .C2(new_n868_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n869_), .A2(new_n651_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n877_), .B1(new_n878_), .B2(new_n879_), .ZN(G1354gat));
  INV_X1    g679(.A(G218gat), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n869_), .A2(new_n881_), .A3(new_n813_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n573_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n881_), .B2(new_n883_), .ZN(G1355gat));
endmodule


