//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 1 0 1 0 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 1 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n887_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n919_, new_n920_, new_n922_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n936_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT21), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G218gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G211gat), .ZN(new_n208_));
  INV_X1    g007(.A(G211gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G218gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT91), .ZN(new_n211_));
  AND3_X1   g010(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n211_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  AND2_X1   g013(.A1(G197gat), .A2(G204gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G197gat), .A2(G204gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n205_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT90), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n206_), .B1(new_n214_), .B2(new_n219_), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n204_), .A2(new_n205_), .ZN(new_n221_));
  AOI21_X1  g020(.A(KEYINPUT90), .B1(new_n204_), .B2(new_n205_), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n221_), .B(new_n222_), .C1(new_n212_), .C2(new_n213_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n220_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT22), .B(G169gat), .ZN(new_n225_));
  INV_X1    g024(.A(G176gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT80), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n227_), .B(new_n230_), .C1(new_n233_), .C2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT79), .ZN(new_n236_));
  INV_X1    g035(.A(G169gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n236_), .A2(new_n237_), .A3(new_n226_), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT79), .B1(G169gat), .B2(G176gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT24), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT26), .B(G190gat), .ZN(new_n243_));
  INV_X1    g042(.A(G183gat), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT25), .B1(new_n244_), .B2(KEYINPUT78), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT78), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT25), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n246_), .A2(new_n247_), .A3(G183gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n243_), .A2(new_n245_), .A3(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n231_), .B(KEYINPUT23), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n242_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n228_), .B(KEYINPUT80), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n238_), .A2(KEYINPUT24), .A3(new_n239_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n235_), .B1(new_n251_), .B2(new_n254_), .ZN(new_n255_));
  OAI211_X1 g054(.A(KEYINPUT94), .B(KEYINPUT20), .C1(new_n224_), .C2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n250_), .B1(G183gat), .B2(G190gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT95), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n225_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT22), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n260_), .A2(G169gat), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n237_), .A2(KEYINPUT22), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT95), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n259_), .A2(new_n263_), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n257_), .B(new_n230_), .C1(new_n264_), .C2(G176gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT25), .B(G183gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n243_), .A2(new_n266_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n238_), .A2(KEYINPUT24), .A3(new_n228_), .A4(new_n239_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n242_), .A2(new_n250_), .A3(new_n267_), .A4(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n265_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(new_n224_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n256_), .A2(new_n271_), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n252_), .A2(new_n253_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n273_), .A2(new_n250_), .A3(new_n249_), .A4(new_n242_), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n274_), .A2(new_n220_), .A3(new_n223_), .A4(new_n235_), .ZN(new_n275_));
  AOI21_X1  g074(.A(KEYINPUT94), .B1(new_n275_), .B2(KEYINPUT20), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n203_), .B1(new_n272_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n224_), .A2(new_n255_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n265_), .A2(new_n220_), .A3(new_n223_), .A4(new_n269_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n203_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n278_), .A2(new_n279_), .A3(KEYINPUT20), .A4(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n277_), .A2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G8gat), .B(G36gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT18), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G64gat), .B(G92gat), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n284_), .B(new_n285_), .Z(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n282_), .A2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n277_), .A2(new_n286_), .A3(new_n281_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT27), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(KEYINPUT98), .B(KEYINPUT20), .Z(new_n293_));
  NAND3_X1  g092(.A1(new_n278_), .A2(new_n279_), .A3(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(new_n203_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT99), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n294_), .A2(KEYINPUT99), .A3(new_n203_), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT20), .B1(new_n224_), .B2(new_n255_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT94), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(new_n271_), .A3(new_n256_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n297_), .B(new_n298_), .C1(new_n203_), .C2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n287_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n304_), .A2(KEYINPUT27), .A3(new_n289_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n292_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(KEYINPUT87), .A2(G155gat), .A3(G162gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(KEYINPUT87), .B1(G155gat), .B2(G162gat), .ZN(new_n309_));
  OAI22_X1  g108(.A1(new_n308_), .A2(new_n309_), .B1(G155gat), .B2(G162gat), .ZN(new_n310_));
  NOR2_X1   g109(.A1(G141gat), .A2(G148gat), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT3), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n311_), .A2(KEYINPUT88), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT88), .ZN(new_n314_));
  OAI22_X1  g113(.A1(new_n314_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G141gat), .A2(G148gat), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n316_), .A2(KEYINPUT2), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(KEYINPUT2), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n313_), .B(new_n315_), .C1(new_n317_), .C2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n310_), .B1(new_n319_), .B2(KEYINPUT89), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n316_), .B(KEYINPUT2), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT89), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n321_), .A2(new_n322_), .A3(new_n315_), .A4(new_n313_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n309_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT1), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(new_n325_), .A3(new_n307_), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT1), .B1(new_n308_), .B2(new_n309_), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n326_), .B(new_n327_), .C1(G155gat), .C2(G162gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n316_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n329_), .A2(new_n311_), .ZN(new_n330_));
  AOI22_X1  g129(.A1(new_n320_), .A2(new_n323_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT29), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n224_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT92), .ZN(new_n334_));
  INV_X1    g133(.A(G228gat), .ZN(new_n335_));
  INV_X1    g134(.A(G233gat), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n334_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G78gat), .B(G106gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT93), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n333_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n339_), .B1(new_n333_), .B2(new_n337_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G22gat), .B(G50gat), .ZN(new_n343_));
  OR3_X1    g142(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n319_), .A2(KEYINPUT89), .ZN(new_n345_));
  INV_X1    g144(.A(new_n310_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(new_n323_), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n328_), .A2(new_n330_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  OR3_X1    g148(.A1(new_n349_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT28), .B1(new_n349_), .B2(KEYINPUT29), .ZN(new_n351_));
  NAND3_X1  g150(.A1(KEYINPUT92), .A2(G228gat), .A3(G233gat), .ZN(new_n352_));
  AND3_X1   g151(.A1(new_n350_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n352_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n343_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n344_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n355_), .B1(new_n344_), .B2(new_n356_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n306_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G127gat), .B(G134gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G113gat), .B(G120gat), .ZN(new_n363_));
  AND3_X1   g162(.A1(new_n362_), .A2(new_n363_), .A3(KEYINPUT84), .ZN(new_n364_));
  AOI21_X1  g163(.A(KEYINPUT84), .B1(new_n362_), .B2(new_n363_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT85), .B1(new_n362_), .B2(new_n363_), .ZN(new_n367_));
  INV_X1    g166(.A(G134gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(G127gat), .ZN(new_n369_));
  INV_X1    g168(.A(G127gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(G134gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(G120gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(G113gat), .ZN(new_n374_));
  INV_X1    g173(.A(G113gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(G120gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT85), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n372_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n367_), .A2(new_n379_), .ZN(new_n380_));
  NOR3_X1   g179(.A1(new_n366_), .A2(new_n380_), .A3(KEYINPUT86), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT86), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n372_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n378_), .B1(new_n372_), .B2(new_n377_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT84), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n386_), .B1(new_n372_), .B2(new_n377_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n362_), .A2(new_n363_), .A3(KEYINPUT84), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n382_), .B1(new_n385_), .B2(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n381_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT31), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT83), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT81), .B(KEYINPUT30), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n255_), .B(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n396_), .A2(KEYINPUT82), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n394_), .B(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(KEYINPUT82), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G71gat), .B(G99gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(G43gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G227gat), .A2(G233gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(G15gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n401_), .B(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n399_), .A2(new_n404_), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n398_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n398_), .A2(new_n405_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G1gat), .B(G29gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(G85gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT0), .B(G57gat), .ZN(new_n412_));
  XOR2_X1   g211(.A(new_n411_), .B(new_n412_), .Z(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT86), .B1(new_n366_), .B2(new_n380_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n385_), .A2(new_n382_), .A3(new_n389_), .ZN(new_n416_));
  AOI22_X1  g215(.A1(new_n415_), .A2(new_n416_), .B1(new_n348_), .B2(new_n347_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT4), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G225gat), .A2(G233gat), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT97), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT96), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n362_), .B(new_n363_), .ZN(new_n425_));
  AND4_X1   g224(.A1(new_n424_), .A2(new_n347_), .A3(new_n348_), .A4(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n349_), .B1(new_n381_), .B2(new_n390_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n424_), .B1(new_n331_), .B2(new_n425_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n426_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n423_), .B1(new_n429_), .B2(new_n418_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n331_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n347_), .A2(new_n348_), .A3(new_n425_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT96), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n431_), .B1(new_n417_), .B2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n434_), .A2(KEYINPUT97), .A3(KEYINPUT4), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n422_), .B1(new_n430_), .B2(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n429_), .A2(new_n421_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n414_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n422_), .ZN(new_n439_));
  NOR3_X1   g238(.A1(new_n429_), .A2(new_n423_), .A3(new_n418_), .ZN(new_n440_));
  AOI21_X1  g239(.A(KEYINPUT97), .B1(new_n434_), .B2(KEYINPUT4), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n439_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n437_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n443_), .A3(new_n413_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n438_), .A2(new_n444_), .ZN(new_n445_));
  NOR3_X1   g244(.A1(new_n361_), .A2(new_n409_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n286_), .A2(KEYINPUT32), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n303_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n277_), .A2(new_n447_), .A3(new_n281_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n451_), .B1(new_n444_), .B2(new_n438_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n419_), .A2(new_n420_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n453_), .B1(new_n430_), .B2(new_n435_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n414_), .B1(new_n429_), .B2(new_n420_), .ZN(new_n455_));
  OAI211_X1 g254(.A(new_n289_), .B(new_n288_), .C1(new_n454_), .C2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT33), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n456_), .B1(new_n457_), .B2(new_n444_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n430_), .A2(new_n435_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n437_), .B1(new_n459_), .B2(new_n439_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(KEYINPUT33), .A3(new_n413_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n452_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT100), .B1(new_n462_), .B2(new_n359_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n444_), .A2(new_n457_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n453_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n455_), .B1(new_n459_), .B2(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n466_), .A2(new_n290_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n464_), .A2(new_n467_), .A3(new_n461_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n451_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n445_), .A2(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n359_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT100), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n306_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n438_), .A2(new_n444_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(new_n359_), .A3(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n463_), .A2(new_n473_), .A3(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n446_), .B1(new_n477_), .B2(new_n409_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G15gat), .B(G22gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT71), .B(G8gat), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n480_), .A2(G1gat), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT14), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n479_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G1gat), .B(G8gat), .ZN(new_n484_));
  XOR2_X1   g283(.A(new_n483_), .B(new_n484_), .Z(new_n485_));
  XNOR2_X1  g284(.A(G29gat), .B(G36gat), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT69), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G43gat), .B(G50gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n485_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT77), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n485_), .A2(new_n490_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G229gat), .A2(G233gat), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n485_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n490_), .B(KEYINPUT15), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n493_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n498_), .B1(new_n497_), .B2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G113gat), .B(G141gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G169gat), .B(G197gat), .ZN(new_n504_));
  XOR2_X1   g303(.A(new_n503_), .B(new_n504_), .Z(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n502_), .B(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n478_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(G230gat), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n509_), .A2(new_n336_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G57gat), .B(G64gat), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n512_), .A2(KEYINPUT11), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(KEYINPUT11), .ZN(new_n514_));
  XOR2_X1   g313(.A(G71gat), .B(G78gat), .Z(new_n515_));
  NAND3_X1  g314(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n514_), .A2(new_n515_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT7), .ZN(new_n520_));
  INV_X1    g319(.A(G99gat), .ZN(new_n521_));
  INV_X1    g320(.A(G106gat), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n520_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT65), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n523_), .A2(KEYINPUT65), .A3(new_n524_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G99gat), .A2(G106gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT6), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n527_), .A2(new_n528_), .A3(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(G85gat), .B(G92gat), .Z(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT8), .B1(new_n533_), .B2(KEYINPUT66), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT66), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n535_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n525_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(new_n530_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT64), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n537_), .A2(new_n530_), .A3(KEYINPUT64), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT8), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n532_), .A2(new_n543_), .ZN(new_n544_));
  OAI22_X1  g343(.A1(new_n534_), .A2(new_n536_), .B1(new_n542_), .B2(new_n544_), .ZN(new_n545_));
  XOR2_X1   g344(.A(KEYINPUT10), .B(G99gat), .Z(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n522_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n532_), .A2(KEYINPUT9), .ZN(new_n548_));
  INV_X1    g347(.A(G85gat), .ZN(new_n549_));
  INV_X1    g348(.A(G92gat), .ZN(new_n550_));
  OR3_X1    g349(.A1(new_n549_), .A2(new_n550_), .A3(KEYINPUT9), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n547_), .A2(new_n548_), .A3(new_n530_), .A4(new_n551_), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n545_), .A2(KEYINPUT67), .A3(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(KEYINPUT67), .B1(new_n545_), .B2(new_n552_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n519_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT67), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n544_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n531_), .A2(new_n532_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n543_), .B1(new_n558_), .B2(new_n535_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n536_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n557_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n552_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n556_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n545_), .A2(KEYINPUT67), .A3(new_n552_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n563_), .A2(new_n518_), .A3(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n511_), .B1(new_n555_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n545_), .A2(new_n552_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n567_), .A2(KEYINPUT12), .A3(new_n519_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT12), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n569_), .B1(new_n555_), .B2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n553_), .A2(new_n554_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n510_), .B1(new_n572_), .B2(new_n518_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n566_), .B1(new_n571_), .B2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G120gat), .B(G148gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT5), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G176gat), .B(G204gat), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n576_), .B(new_n577_), .Z(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n574_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n574_), .A2(new_n579_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT13), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n580_), .B(new_n581_), .C1(KEYINPUT68), .C2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n567_), .A2(new_n500_), .A3(KEYINPUT70), .ZN(new_n588_));
  AOI21_X1  g387(.A(KEYINPUT70), .B1(new_n567_), .B2(new_n500_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n572_), .A2(new_n490_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT34), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT35), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n592_), .A2(new_n596_), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n563_), .A2(new_n490_), .A3(new_n564_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n567_), .A2(new_n500_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n594_), .A2(KEYINPUT35), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n596_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  OR3_X1    g401(.A1(new_n598_), .A2(new_n599_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT36), .ZN(new_n604_));
  XOR2_X1   g403(.A(G134gat), .B(G162gat), .Z(new_n605_));
  XNOR2_X1  g404(.A(G190gat), .B(G218gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n597_), .A2(new_n603_), .A3(new_n604_), .A4(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n604_), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n607_), .A2(new_n604_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n595_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n598_), .A2(new_n599_), .A3(new_n602_), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n609_), .B(new_n610_), .C1(new_n611_), .C2(new_n612_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n608_), .A2(new_n613_), .A3(KEYINPUT37), .ZN(new_n614_));
  AOI21_X1  g413(.A(KEYINPUT37), .B1(new_n608_), .B2(new_n613_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n518_), .B(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n499_), .B(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(KEYINPUT73), .B(KEYINPUT16), .Z(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT74), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G127gat), .B(G155gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G183gat), .B(G211gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n625_), .A2(KEYINPUT72), .A3(KEYINPUT17), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n619_), .B(new_n626_), .C1(KEYINPUT17), .C2(new_n625_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n627_), .B1(new_n619_), .B2(new_n626_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT75), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n616_), .A2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT76), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n508_), .A2(new_n587_), .A3(new_n631_), .ZN(new_n632_));
  OR3_X1    g431(.A1(new_n632_), .A2(G1gat), .A3(new_n475_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n634_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n608_), .A2(new_n613_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n478_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n587_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n640_), .A2(new_n507_), .A3(new_n628_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G1gat), .B1(new_n642_), .B2(new_n475_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n635_), .A2(new_n636_), .A3(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT102), .ZN(G1324gat));
  OAI21_X1  g444(.A(G8gat), .B1(new_n642_), .B2(new_n474_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT39), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n474_), .A2(new_n480_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n647_), .B1(new_n632_), .B2(new_n648_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g449(.A(G15gat), .B1(new_n642_), .B2(new_n409_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n652_), .ZN(new_n654_));
  OR3_X1    g453(.A1(new_n632_), .A2(G15gat), .A3(new_n409_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n653_), .A2(new_n654_), .A3(new_n655_), .ZN(G1326gat));
  INV_X1    g455(.A(new_n359_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G22gat), .B1(new_n642_), .B2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT42), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n657_), .A2(G22gat), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT104), .Z(new_n661_));
  OAI21_X1  g460(.A(new_n659_), .B1(new_n632_), .B2(new_n661_), .ZN(G1327gat));
  NOR3_X1   g461(.A1(new_n640_), .A2(new_n629_), .A3(new_n637_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n508_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  OR3_X1    g464(.A1(new_n665_), .A2(G29gat), .A3(new_n475_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n476_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n667_));
  AOI211_X1 g466(.A(KEYINPUT100), .B(new_n359_), .C1(new_n468_), .C2(new_n470_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n409_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n446_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n616_), .A2(KEYINPUT43), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n674_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT37), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n637_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n608_), .A2(new_n613_), .A3(KEYINPUT37), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n677_), .A2(KEYINPUT105), .A3(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n675_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n475_), .A2(new_n359_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n682_), .A2(new_n306_), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT33), .B1(new_n460_), .B2(new_n413_), .ZN(new_n684_));
  NOR4_X1   g483(.A1(new_n436_), .A2(new_n457_), .A3(new_n437_), .A4(new_n414_), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n684_), .A2(new_n685_), .A3(new_n456_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n657_), .B1(new_n686_), .B2(new_n452_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n683_), .B1(new_n687_), .B2(KEYINPUT100), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n408_), .B1(new_n688_), .B2(new_n473_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n681_), .B1(new_n689_), .B2(new_n446_), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT106), .B1(new_n690_), .B2(KEYINPUT43), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n680_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n692_), .A2(new_n693_), .A3(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n673_), .B1(new_n691_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n507_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n629_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n587_), .A2(new_n697_), .A3(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n696_), .A2(KEYINPUT44), .A3(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702_));
  INV_X1    g501(.A(new_n673_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n693_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n704_));
  OAI211_X1 g503(.A(KEYINPUT106), .B(KEYINPUT43), .C1(new_n478_), .C2(new_n680_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n703_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n702_), .B1(new_n706_), .B2(new_n699_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n701_), .A2(new_n707_), .A3(new_n445_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n708_), .A2(new_n709_), .A3(G29gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n708_), .B2(G29gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n666_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT108), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n714_), .B(new_n666_), .C1(new_n710_), .C2(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1328gat));
  NAND3_X1  g515(.A1(new_n701_), .A2(new_n707_), .A3(new_n306_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(G36gat), .ZN(new_n718_));
  INV_X1    g517(.A(G36gat), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n664_), .A2(new_n719_), .A3(new_n306_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT45), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n718_), .A2(new_n721_), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT46), .Z(G1329gat));
  AND2_X1   g522(.A1(new_n701_), .A2(new_n707_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n724_), .A2(G43gat), .A3(new_n408_), .ZN(new_n725_));
  INV_X1    g524(.A(G43gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n726_), .B1(new_n665_), .B2(new_n409_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g528(.A(G50gat), .B1(new_n664_), .B2(new_n359_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n359_), .A2(G50gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n724_), .B2(new_n731_), .ZN(G1331gat));
  NOR2_X1   g531(.A1(new_n697_), .A2(new_n698_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n639_), .A2(new_n640_), .A3(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G57gat), .B1(new_n734_), .B2(new_n475_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n631_), .A2(new_n640_), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n736_), .A2(KEYINPUT109), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n478_), .A2(new_n697_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(KEYINPUT109), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n737_), .A2(new_n738_), .A3(new_n739_), .ZN(new_n740_));
  OR2_X1    g539(.A1(new_n475_), .A2(G57gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n735_), .B1(new_n740_), .B2(new_n741_), .ZN(G1332gat));
  OAI21_X1  g541(.A(G64gat), .B1(new_n734_), .B2(new_n474_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT48), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n474_), .A2(G64gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n744_), .B1(new_n740_), .B2(new_n745_), .ZN(G1333gat));
  OAI21_X1  g545(.A(G71gat), .B1(new_n734_), .B2(new_n409_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT49), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n409_), .A2(G71gat), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT110), .Z(new_n750_));
  OAI21_X1  g549(.A(new_n748_), .B1(new_n740_), .B2(new_n750_), .ZN(G1334gat));
  OAI21_X1  g550(.A(G78gat), .B1(new_n734_), .B2(new_n657_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT50), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n657_), .A2(G78gat), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n753_), .B1(new_n740_), .B2(new_n754_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT111), .Z(G1335gat));
  NOR3_X1   g555(.A1(new_n587_), .A2(new_n629_), .A3(new_n637_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n738_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(new_n549_), .A3(new_n445_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n640_), .A2(new_n507_), .A3(new_n698_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n706_), .A2(new_n475_), .A3(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n759_), .B1(new_n761_), .B2(new_n549_), .ZN(G1336gat));
  NAND3_X1  g561(.A1(new_n758_), .A2(new_n550_), .A3(new_n306_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n706_), .A2(new_n474_), .A3(new_n760_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(new_n550_), .ZN(G1337gat));
  NAND3_X1  g564(.A1(new_n758_), .A2(new_n408_), .A3(new_n546_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT112), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT51), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n706_), .A2(new_n409_), .A3(new_n760_), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n767_), .B(new_n769_), .C1(new_n521_), .C2(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n768_), .A2(KEYINPUT51), .ZN(new_n772_));
  XOR2_X1   g571(.A(new_n771_), .B(new_n772_), .Z(G1338gat));
  NAND3_X1  g572(.A1(new_n758_), .A2(new_n522_), .A3(new_n359_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n706_), .A2(new_n760_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n359_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n775_), .B1(new_n777_), .B2(G106gat), .ZN(new_n778_));
  AOI211_X1 g577(.A(KEYINPUT52), .B(new_n522_), .C1(new_n776_), .C2(new_n359_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n774_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n780_), .B(new_n782_), .ZN(G1339gat));
  NAND3_X1  g582(.A1(new_n587_), .A2(new_n733_), .A3(new_n616_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n784_), .A2(KEYINPUT54), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(KEYINPUT54), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT119), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n788_), .A2(KEYINPUT57), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n506_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT118), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n791_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n501_), .A2(new_n497_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n792_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n502_), .A2(new_n505_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n797_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n581_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n507_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n518_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n568_), .B1(new_n803_), .B2(KEYINPUT12), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n565_), .A2(new_n511_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n802_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n571_), .A2(new_n573_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n809_), .A2(new_n802_), .A3(KEYINPUT55), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n511_), .B1(new_n571_), .B2(new_n565_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT116), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n815_));
  AOI211_X1 g614(.A(new_n815_), .B(new_n812_), .C1(new_n808_), .C2(new_n810_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n578_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT56), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT117), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n801_), .B1(new_n817_), .B2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT55), .B1(new_n809_), .B2(new_n802_), .ZN(new_n821_));
  AOI211_X1 g620(.A(KEYINPUT115), .B(new_n807_), .C1(new_n571_), .C2(new_n573_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n813_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n815_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n811_), .A2(KEYINPUT116), .A3(new_n813_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n579_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n819_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n798_), .B1(new_n820_), .B2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n789_), .B1(new_n829_), .B2(new_n638_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n798_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n800_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n817_), .A2(new_n819_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n831_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n789_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n834_), .A2(new_n637_), .A3(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT58), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n797_), .A2(new_n799_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n826_), .B2(new_n818_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n817_), .A2(KEYINPUT56), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n837_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n616_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n817_), .A2(KEYINPUT56), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n826_), .A2(new_n818_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n843_), .A2(new_n844_), .A3(KEYINPUT58), .A4(new_n838_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n841_), .A2(new_n842_), .A3(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n830_), .A2(new_n836_), .A3(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n787_), .B1(new_n847_), .B2(new_n628_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n361_), .A2(new_n409_), .A3(new_n475_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  OAI211_X1 g650(.A(KEYINPUT120), .B(new_n375_), .C1(new_n851_), .C2(new_n507_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n853_));
  INV_X1    g652(.A(new_n850_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n848_), .A2(new_n507_), .A3(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n853_), .B1(new_n855_), .B2(G113gat), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n852_), .A2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n787_), .B1(new_n847_), .B2(new_n698_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n858_), .A2(KEYINPUT59), .A3(new_n854_), .ZN(new_n859_));
  OAI21_X1  g658(.A(KEYINPUT59), .B1(new_n848_), .B2(new_n854_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  OAI211_X1 g661(.A(KEYINPUT121), .B(KEYINPUT59), .C1(new_n848_), .C2(new_n854_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n859_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n507_), .A2(new_n375_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n857_), .B1(new_n864_), .B2(new_n865_), .ZN(G1340gat));
  OAI21_X1  g665(.A(new_n373_), .B1(new_n587_), .B2(KEYINPUT60), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n867_), .B1(KEYINPUT60), .B2(new_n373_), .ZN(new_n868_));
  OR2_X1    g667(.A1(new_n851_), .A2(new_n868_), .ZN(new_n869_));
  AOI211_X1 g668(.A(new_n587_), .B(new_n859_), .C1(new_n862_), .C2(new_n863_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n870_), .B2(new_n373_), .ZN(G1341gat));
  OAI211_X1 g670(.A(KEYINPUT122), .B(new_n370_), .C1(new_n851_), .C2(new_n698_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n848_), .A2(new_n698_), .A3(new_n854_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n874_), .B2(G127gat), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n872_), .A2(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n628_), .A2(new_n370_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n876_), .B1(new_n864_), .B2(new_n877_), .ZN(G1342gat));
  NAND4_X1  g677(.A1(new_n849_), .A2(new_n368_), .A3(new_n638_), .A4(new_n850_), .ZN(new_n879_));
  AOI211_X1 g678(.A(new_n616_), .B(new_n859_), .C1(new_n862_), .C2(new_n863_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(new_n368_), .ZN(G1343gat));
  NOR4_X1   g680(.A1(new_n408_), .A2(new_n657_), .A3(new_n475_), .A4(new_n306_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n848_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n697_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n640_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g687(.A1(new_n884_), .A2(new_n629_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(KEYINPUT123), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT123), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n884_), .A2(new_n891_), .A3(new_n629_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(KEYINPUT61), .B(G155gat), .ZN(new_n893_));
  AND3_X1   g692(.A1(new_n890_), .A2(new_n892_), .A3(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n893_), .B1(new_n890_), .B2(new_n892_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1346gat));
  AOI21_X1  g695(.A(G162gat), .B1(new_n884_), .B2(new_n638_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n681_), .A2(G162gat), .ZN(new_n898_));
  XOR2_X1   g697(.A(new_n898_), .B(KEYINPUT124), .Z(new_n899_));
  AOI21_X1  g698(.A(new_n897_), .B1(new_n884_), .B2(new_n899_), .ZN(G1347gat));
  NOR2_X1   g699(.A1(new_n409_), .A2(new_n445_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n901_), .A2(new_n657_), .A3(new_n306_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n858_), .A2(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n237_), .B1(new_n903_), .B2(new_n697_), .ZN(new_n904_));
  OR2_X1    g703(.A1(new_n904_), .A2(KEYINPUT62), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(KEYINPUT62), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n903_), .A2(new_n697_), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n905_), .B(new_n906_), .C1(new_n264_), .C2(new_n907_), .ZN(G1348gat));
  INV_X1    g707(.A(KEYINPUT125), .ZN(new_n909_));
  INV_X1    g708(.A(new_n902_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n849_), .A2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n640_), .A2(G176gat), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n858_), .A2(new_n587_), .A3(new_n902_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n914_), .A2(G176gat), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n909_), .B1(new_n913_), .B2(new_n915_), .ZN(new_n916_));
  OAI221_X1 g715(.A(KEYINPUT125), .B1(new_n914_), .B2(G176gat), .C1(new_n911_), .C2(new_n912_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1349gat));
  NAND3_X1  g717(.A1(new_n849_), .A2(new_n629_), .A3(new_n910_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n628_), .A2(new_n266_), .ZN(new_n920_));
  AOI22_X1  g719(.A1(new_n919_), .A2(new_n244_), .B1(new_n903_), .B2(new_n920_), .ZN(G1350gat));
  NAND3_X1  g720(.A1(new_n903_), .A2(new_n243_), .A3(new_n638_), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n858_), .A2(new_n616_), .A3(new_n902_), .ZN(new_n923_));
  INV_X1    g722(.A(G190gat), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n922_), .B1(new_n923_), .B2(new_n924_), .ZN(G1351gat));
  XNOR2_X1  g724(.A(KEYINPUT127), .B(G197gat), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT127), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n927_), .A2(G197gat), .ZN(new_n928_));
  OR2_X1    g727(.A1(new_n408_), .A2(new_n682_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT126), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n306_), .B1(new_n929_), .B2(new_n930_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n931_), .B1(new_n930_), .B2(new_n929_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n849_), .A2(new_n932_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n933_), .A2(new_n507_), .ZN(new_n934_));
  MUX2_X1   g733(.A(new_n926_), .B(new_n928_), .S(new_n934_), .Z(G1352gat));
  INV_X1    g734(.A(new_n933_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(new_n640_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g737(.A1(new_n933_), .A2(new_n628_), .ZN(new_n939_));
  OR2_X1    g738(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  XOR2_X1   g740(.A(KEYINPUT63), .B(G211gat), .Z(new_n942_));
  AOI21_X1  g741(.A(new_n941_), .B1(new_n939_), .B2(new_n942_), .ZN(G1354gat));
  OAI21_X1  g742(.A(G218gat), .B1(new_n933_), .B2(new_n616_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n638_), .A2(new_n207_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n944_), .B1(new_n933_), .B2(new_n945_), .ZN(G1355gat));
endmodule


