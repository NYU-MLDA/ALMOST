//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n659_, new_n660_, new_n661_,
    new_n663_, new_n664_, new_n665_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n786_, new_n787_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n794_, new_n796_, new_n797_, new_n799_, new_n800_,
    new_n801_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n822_, new_n823_, new_n824_, new_n826_, new_n827_, new_n828_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_;
  XNOR2_X1  g000(.A(G85gat), .B(G92gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT6), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT6), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n206_), .A2(G99gat), .A3(G106gat), .ZN(new_n207_));
  AND2_X1   g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT7), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n203_), .B1(new_n208_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT8), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(KEYINPUT66), .A3(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT9), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n202_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT10), .B(G99gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT64), .B(G106gat), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n205_), .A2(new_n207_), .ZN(new_n225_));
  INV_X1    g024(.A(G92gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT65), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(G92gat), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n227_), .A2(new_n229_), .A3(new_n217_), .A4(G85gat), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n219_), .A2(new_n224_), .A3(new_n225_), .A4(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n232_), .B(new_n203_), .C1(new_n208_), .C2(new_n213_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT8), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n225_), .A2(new_n212_), .A3(new_n211_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n232_), .B1(new_n235_), .B2(new_n203_), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n216_), .B(new_n231_), .C1(new_n234_), .C2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G57gat), .B(G64gat), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n238_), .A2(KEYINPUT11), .ZN(new_n239_));
  XOR2_X1   g038(.A(G71gat), .B(G78gat), .Z(new_n240_));
  OR2_X1    g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n238_), .A2(KEYINPUT11), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n239_), .A2(new_n240_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n237_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT68), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT67), .B1(new_n237_), .B2(new_n244_), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n230_), .B(new_n225_), .C1(new_n220_), .C2(new_n222_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n248_), .A2(new_n218_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n212_), .ZN(new_n250_));
  NOR3_X1   g049(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n202_), .B1(new_n252_), .B2(new_n225_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n215_), .B1(new_n253_), .B2(new_n232_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n214_), .A2(KEYINPUT66), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n249_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n256_), .A2(new_n257_), .A3(new_n258_), .A4(new_n216_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n237_), .A2(new_n260_), .A3(new_n244_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n246_), .A2(new_n247_), .A3(new_n259_), .A4(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G230gat), .A2(G233gat), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n245_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n256_), .A2(new_n257_), .A3(new_n216_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n237_), .A2(KEYINPUT12), .A3(new_n244_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n268_), .A2(new_n263_), .A3(new_n269_), .A4(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G120gat), .B(G148gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT5), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(G176gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(G204gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n265_), .A2(new_n271_), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n265_), .A2(KEYINPUT70), .A3(new_n271_), .A4(new_n275_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n265_), .A2(new_n271_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n275_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n280_), .A2(KEYINPUT71), .A3(new_n283_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT72), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n288_), .B1(new_n289_), .B2(KEYINPUT13), .ZN(new_n290_));
  XOR2_X1   g089(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n291_));
  NAND3_X1  g090(.A1(new_n286_), .A2(new_n287_), .A3(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT75), .B(G15gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(G22gat), .ZN(new_n296_));
  INV_X1    g095(.A(G1gat), .ZN(new_n297_));
  INV_X1    g096(.A(G8gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT14), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(G1gat), .B(G8gat), .Z(new_n301_));
  XOR2_X1   g100(.A(new_n300_), .B(new_n301_), .Z(new_n302_));
  XNOR2_X1  g101(.A(G29gat), .B(G36gat), .ZN(new_n303_));
  INV_X1    g102(.A(G43gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(G50gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n307_), .A2(KEYINPUT15), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(KEYINPUT15), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n302_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT78), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n307_), .B(KEYINPUT15), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT78), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n312_), .A2(new_n313_), .A3(new_n302_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G229gat), .A2(G233gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n307_), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n302_), .A2(new_n316_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n311_), .A2(new_n314_), .A3(new_n315_), .A4(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n302_), .B(new_n316_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n315_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G113gat), .B(G141gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT79), .ZN(new_n324_));
  INV_X1    g123(.A(G169gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n326_), .B(G197gat), .Z(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n322_), .A2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n318_), .A2(new_n321_), .A3(new_n327_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n294_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G127gat), .B(G134gat), .ZN(new_n334_));
  INV_X1    g133(.A(G113gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(G120gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G183gat), .A2(G190gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT23), .ZN(new_n339_));
  OR3_X1    g138(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n340_));
  INV_X1    g139(.A(G176gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n325_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G169gat), .A2(G176gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n342_), .A2(KEYINPUT24), .A3(new_n343_), .ZN(new_n344_));
  AND3_X1   g143(.A1(new_n339_), .A2(new_n340_), .A3(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT25), .B(G183gat), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n346_), .A2(KEYINPUT80), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT26), .B(G190gat), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT80), .ZN(new_n349_));
  INV_X1    g148(.A(G183gat), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n350_), .A2(KEYINPUT25), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n348_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n345_), .B1(new_n347_), .B2(new_n352_), .ZN(new_n353_));
  OR2_X1    g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354_));
  AOI22_X1  g153(.A1(new_n339_), .A2(new_n354_), .B1(G169gat), .B2(G176gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT22), .B(G169gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT81), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n357_), .B1(new_n325_), .B2(KEYINPUT22), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n341_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n355_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n353_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n337_), .B(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(KEYINPUT30), .B(G71gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT82), .B(G99gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT31), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G15gat), .B(G43gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n367_), .B(new_n368_), .Z(new_n369_));
  NAND2_X1  g168(.A1(G227gat), .A2(G233gat), .ZN(new_n370_));
  XOR2_X1   g169(.A(new_n369_), .B(new_n370_), .Z(new_n371_));
  XNOR2_X1  g170(.A(new_n365_), .B(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT91), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G211gat), .B(G218gat), .ZN(new_n375_));
  XOR2_X1   g174(.A(G197gat), .B(G204gat), .Z(new_n376_));
  OAI21_X1  g175(.A(new_n375_), .B1(new_n376_), .B2(KEYINPUT21), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(KEYINPUT21), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(new_n361_), .A3(new_n353_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n356_), .B(KEYINPUT89), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n341_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n348_), .A2(new_n346_), .ZN(new_n383_));
  AOI22_X1  g182(.A1(new_n382_), .A2(new_n355_), .B1(new_n383_), .B2(new_n345_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n380_), .B(KEYINPUT20), .C1(new_n384_), .C2(new_n379_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G226gat), .A2(G233gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT19), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n385_), .A2(KEYINPUT90), .A3(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT90), .B1(new_n385_), .B2(new_n387_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT20), .ZN(new_n390_));
  XOR2_X1   g189(.A(new_n377_), .B(new_n378_), .Z(new_n391_));
  AOI21_X1  g190(.A(new_n390_), .B1(new_n391_), .B2(new_n362_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n387_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n384_), .A2(new_n379_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n392_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n388_), .A2(new_n389_), .A3(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G8gat), .B(G36gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT18), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(G64gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(new_n226_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n374_), .B1(new_n397_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n397_), .A2(new_n401_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n385_), .A2(new_n387_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT90), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n385_), .A2(KEYINPUT90), .A3(new_n387_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(new_n395_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n401_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(KEYINPUT91), .A3(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n402_), .A2(new_n403_), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT27), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G228gat), .A2(G233gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT86), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(G155gat), .A2(G162gat), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT83), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G155gat), .A2(G162gat), .ZN(new_n420_));
  NOR2_X1   g219(.A1(G141gat), .A2(G148gat), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT3), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(KEYINPUT84), .A2(KEYINPUT2), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G141gat), .A2(G148gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  AOI22_X1  g225(.A1(KEYINPUT84), .A2(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n426_), .B1(new_n427_), .B2(new_n424_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n419_), .B(new_n420_), .C1(new_n423_), .C2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n421_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n417_), .B(KEYINPUT83), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n420_), .B(KEYINPUT1), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n430_), .B(new_n425_), .C1(new_n431_), .C2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n429_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT29), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n416_), .B1(new_n391_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  XOR2_X1   g236(.A(G78gat), .B(G106gat), .Z(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n391_), .A2(new_n435_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n414_), .A2(KEYINPUT86), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n416_), .A2(new_n441_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n437_), .B(new_n439_), .C1(new_n440_), .C2(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n440_), .A2(new_n442_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n438_), .B1(new_n444_), .B2(new_n436_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT88), .B1(new_n446_), .B2(KEYINPUT87), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT87), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT88), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n443_), .A2(new_n445_), .A3(new_n448_), .A4(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n447_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n446_), .A2(KEYINPUT87), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n434_), .A2(KEYINPUT29), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT28), .ZN(new_n454_));
  XOR2_X1   g253(.A(G22gat), .B(G50gat), .Z(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT85), .ZN(new_n456_));
  XOR2_X1   g255(.A(new_n454_), .B(new_n456_), .Z(new_n457_));
  NAND2_X1  g256(.A1(new_n452_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n451_), .A2(new_n458_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n447_), .A2(new_n452_), .A3(new_n457_), .A4(new_n450_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(G120gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n336_), .B(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(new_n433_), .A3(new_n429_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n337_), .A2(new_n434_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(new_n465_), .A3(KEYINPUT4), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT92), .B1(new_n465_), .B2(KEYINPUT4), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G225gat), .A2(G233gat), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT92), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT4), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n337_), .A2(new_n470_), .A3(new_n471_), .A4(new_n434_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n466_), .A2(new_n467_), .A3(new_n469_), .A4(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n464_), .A2(new_n468_), .A3(new_n465_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  XOR2_X1   g274(.A(KEYINPUT93), .B(KEYINPUT0), .Z(new_n476_));
  XNOR2_X1  g275(.A(G1gat), .B(G29gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G57gat), .B(G85gat), .ZN(new_n479_));
  XOR2_X1   g278(.A(new_n478_), .B(new_n479_), .Z(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n475_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n473_), .A2(new_n480_), .A3(new_n474_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n385_), .A2(new_n387_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n393_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n403_), .B(KEYINPUT27), .C1(new_n401_), .C2(new_n488_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n413_), .A2(new_n461_), .A3(new_n485_), .A4(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n408_), .A2(KEYINPUT91), .A3(new_n409_), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT91), .B1(new_n408_), .B2(new_n409_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .A4(new_n472_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n464_), .A2(new_n469_), .A3(new_n465_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(new_n481_), .A3(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n483_), .B(KEYINPUT33), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n494_), .A2(new_n403_), .A3(new_n497_), .A4(new_n498_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n406_), .A2(new_n395_), .A3(KEYINPUT94), .A4(new_n407_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n401_), .A2(KEYINPUT32), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n500_), .A2(new_n501_), .A3(new_n488_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT94), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n501_), .B1(new_n397_), .B2(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n484_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n461_), .B1(new_n499_), .B2(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n373_), .B1(new_n491_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n413_), .A2(new_n489_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n485_), .A2(new_n372_), .ZN(new_n509_));
  NOR3_X1   g308(.A1(new_n508_), .A2(new_n461_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n507_), .A2(new_n511_), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n333_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(KEYINPUT74), .A2(KEYINPUT37), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT74), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT37), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n312_), .A2(new_n237_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n256_), .A2(new_n307_), .A3(new_n216_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G232gat), .A2(G233gat), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n520_), .B(KEYINPUT73), .Z(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT34), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n518_), .B(new_n519_), .C1(KEYINPUT35), .C2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(KEYINPUT35), .ZN(new_n524_));
  XOR2_X1   g323(.A(new_n523_), .B(new_n524_), .Z(new_n525_));
  XNOR2_X1  g324(.A(G190gat), .B(G218gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(G134gat), .ZN(new_n527_));
  INV_X1    g326(.A(G162gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT36), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n525_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n523_), .B(new_n524_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n529_), .A2(new_n530_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n514_), .B(new_n517_), .C1(new_n532_), .C2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n525_), .A2(new_n531_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n538_), .A2(new_n515_), .A3(new_n516_), .A4(new_n535_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G231gat), .A2(G233gat), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n541_), .B(KEYINPUT76), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n302_), .B(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(new_n244_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G127gat), .B(G155gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT16), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(new_n350_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(G211gat), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n544_), .A2(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n548_), .B1(new_n544_), .B2(KEYINPUT77), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT17), .ZN(new_n551_));
  OR3_X1    g350(.A1(new_n549_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n551_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n540_), .A2(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n513_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n556_), .A2(new_n297_), .A3(new_n484_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT38), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n532_), .A2(new_n536_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n560_), .A2(new_n554_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n513_), .A2(new_n561_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n562_), .A2(new_n484_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n558_), .B1(new_n297_), .B2(new_n563_), .ZN(G1324gat));
  NAND3_X1  g363(.A1(new_n556_), .A2(new_n298_), .A3(new_n508_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT39), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n562_), .A2(new_n508_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n566_), .B1(new_n567_), .B2(G8gat), .ZN(new_n568_));
  AOI211_X1 g367(.A(KEYINPUT39), .B(new_n298_), .C1(new_n562_), .C2(new_n508_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n565_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n570_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g370(.A(G15gat), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n572_), .B1(new_n562_), .B2(new_n372_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT41), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n556_), .A2(new_n572_), .A3(new_n372_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(G1326gat));
  INV_X1    g375(.A(G22gat), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n461_), .A2(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n578_), .B(KEYINPUT95), .Z(new_n579_));
  NAND2_X1  g378(.A1(new_n556_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT42), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n562_), .A2(new_n461_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n581_), .B1(new_n582_), .B2(G22gat), .ZN(new_n583_));
  AOI211_X1 g382(.A(KEYINPUT42), .B(new_n577_), .C1(new_n562_), .C2(new_n461_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n580_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT96), .ZN(G1327gat));
  INV_X1    g385(.A(KEYINPUT43), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n512_), .A2(new_n587_), .A3(new_n540_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT97), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n507_), .A2(new_n589_), .A3(new_n511_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n402_), .A2(new_n403_), .A3(new_n410_), .A4(new_n497_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n498_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n505_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n461_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n372_), .B1(new_n595_), .B2(new_n490_), .ZN(new_n596_));
  OAI21_X1  g395(.A(KEYINPUT97), .B1(new_n596_), .B2(new_n510_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n590_), .A2(new_n597_), .A3(new_n540_), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n598_), .A2(KEYINPUT98), .A3(KEYINPUT43), .ZN(new_n599_));
  AOI21_X1  g398(.A(KEYINPUT98), .B1(new_n598_), .B2(KEYINPUT43), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n588_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n601_), .A2(new_n554_), .A3(new_n333_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT44), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n601_), .A2(KEYINPUT44), .A3(new_n554_), .A4(new_n333_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n604_), .A2(new_n484_), .A3(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(G29gat), .ZN(new_n607_));
  INV_X1    g406(.A(new_n554_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n608_), .A2(new_n559_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n513_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT99), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT99), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n513_), .A2(new_n612_), .A3(new_n609_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n485_), .A2(G29gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT100), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n607_), .B1(new_n614_), .B2(new_n616_), .ZN(G1328gat));
  INV_X1    g416(.A(KEYINPUT46), .ZN(new_n618_));
  INV_X1    g417(.A(G36gat), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n605_), .A2(new_n508_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n619_), .B1(new_n620_), .B2(new_n604_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n611_), .A2(new_n619_), .A3(new_n508_), .A4(new_n613_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT45), .Z(new_n623_));
  OAI21_X1  g422(.A(new_n618_), .B1(new_n621_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n604_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n605_), .A2(new_n508_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G36gat), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n622_), .B(KEYINPUT45), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(KEYINPUT46), .A3(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n624_), .A2(new_n629_), .ZN(G1329gat));
  OAI21_X1  g429(.A(new_n304_), .B1(new_n614_), .B2(new_n373_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n605_), .A2(G43gat), .A3(new_n372_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n631_), .B1(new_n625_), .B2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g433(.A(new_n614_), .ZN(new_n635_));
  AOI21_X1  g434(.A(G50gat), .B1(new_n635_), .B2(new_n461_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n605_), .A2(G50gat), .A3(new_n461_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n636_), .B1(new_n637_), .B2(new_n604_), .ZN(G1331gat));
  AOI21_X1  g437(.A(new_n331_), .B1(new_n507_), .B2(new_n511_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n639_), .A2(new_n561_), .A3(new_n294_), .ZN(new_n640_));
  INV_X1    g439(.A(G57gat), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n640_), .A2(new_n641_), .A3(new_n485_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n512_), .A2(new_n332_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT101), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n639_), .A2(KEYINPUT101), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n293_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(new_n555_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n649_), .A2(KEYINPUT102), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(KEYINPUT102), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(new_n484_), .A3(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n642_), .B1(new_n652_), .B2(new_n641_), .ZN(G1332gat));
  INV_X1    g452(.A(new_n508_), .ZN(new_n654_));
  OAI21_X1  g453(.A(G64gat), .B1(new_n640_), .B2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT48), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n654_), .A2(G64gat), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n656_), .B1(new_n648_), .B2(new_n657_), .ZN(G1333gat));
  OAI21_X1  g457(.A(G71gat), .B1(new_n640_), .B2(new_n373_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT49), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n373_), .A2(G71gat), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n660_), .B1(new_n648_), .B2(new_n661_), .ZN(G1334gat));
  OAI21_X1  g461(.A(G78gat), .B1(new_n640_), .B2(new_n594_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT50), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n594_), .A2(G78gat), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n664_), .B1(new_n648_), .B2(new_n665_), .ZN(G1335gat));
  NAND2_X1  g465(.A1(new_n647_), .A2(new_n609_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(G85gat), .B1(new_n668_), .B2(new_n484_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n293_), .A2(new_n608_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n601_), .A2(new_n332_), .A3(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n484_), .A2(G85gat), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT103), .Z(new_n674_));
  AOI21_X1  g473(.A(new_n669_), .B1(new_n672_), .B2(new_n674_), .ZN(G1336gat));
  OAI21_X1  g474(.A(new_n226_), .B1(new_n667_), .B2(new_n654_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n676_), .B(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n508_), .A2(new_n227_), .A3(new_n229_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT105), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n672_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n678_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT106), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n678_), .A2(KEYINPUT106), .A3(new_n681_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1337gat));
  OAI21_X1  g485(.A(G99gat), .B1(new_n671_), .B2(new_n373_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n668_), .A2(new_n221_), .A3(new_n372_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g489(.A1(new_n668_), .A2(new_n223_), .A3(new_n461_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(KEYINPUT107), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n668_), .A2(new_n693_), .A3(new_n223_), .A4(new_n461_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n601_), .A2(new_n332_), .A3(new_n461_), .A4(new_n670_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(G106gat), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT52), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n696_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n695_), .A2(new_n699_), .A3(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT53), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT53), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n695_), .A2(new_n699_), .A3(new_n703_), .A4(new_n700_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(G1339gat));
  AOI21_X1  g504(.A(new_n331_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT54), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n555_), .A2(new_n706_), .A3(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n555_), .B2(new_n706_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n331_), .A2(new_n280_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n257_), .B1(new_n256_), .B2(new_n216_), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n269_), .B(new_n270_), .C1(new_n712_), .C2(new_n266_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n713_), .A2(new_n714_), .A3(new_n264_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n713_), .B2(new_n264_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT55), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n271_), .B(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(KEYINPUT109), .B1(new_n717_), .B2(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n266_), .B1(new_n237_), .B2(new_n244_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n721_), .B1(KEYINPUT12), .B2(new_n712_), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n722_), .A2(new_n718_), .A3(new_n263_), .A4(new_n269_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n271_), .A2(KEYINPUT55), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n725_), .B(new_n726_), .C1(new_n716_), .C2(new_n715_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n720_), .A2(new_n282_), .A3(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT56), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n720_), .A2(KEYINPUT56), .A3(new_n282_), .A4(new_n727_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n711_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n302_), .B(new_n307_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n328_), .B1(new_n733_), .B2(new_n320_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT110), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT110), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n736_), .B(new_n328_), .C1(new_n733_), .C2(new_n320_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n311_), .A2(new_n314_), .A3(new_n320_), .A4(new_n317_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n735_), .A2(new_n737_), .A3(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n330_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n559_), .B1(new_n732_), .B2(new_n741_), .ZN(new_n742_));
  XOR2_X1   g541(.A(KEYINPUT111), .B(KEYINPUT57), .Z(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT112), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n742_), .A2(new_n746_), .A3(new_n743_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(new_n748_));
  OAI211_X1 g547(.A(KEYINPUT57), .B(new_n559_), .C1(new_n732_), .C2(new_n741_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT116), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT114), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n751_), .A2(KEYINPUT58), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT113), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n730_), .A2(new_n753_), .A3(new_n731_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n740_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n755_), .B(new_n280_), .C1(new_n731_), .C2(new_n753_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n752_), .B1(new_n754_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n756_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n752_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n730_), .A2(new_n753_), .A3(new_n731_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n758_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n757_), .A2(new_n540_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT115), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT115), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n757_), .A2(new_n761_), .A3(new_n764_), .A4(new_n540_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n748_), .A2(new_n750_), .A3(new_n763_), .A4(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n710_), .B1(new_n766_), .B2(new_n554_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n654_), .A2(new_n484_), .A3(new_n594_), .A4(new_n372_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(G113gat), .B1(new_n769_), .B2(new_n331_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n750_), .A2(new_n762_), .A3(new_n744_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n710_), .B1(new_n771_), .B2(new_n554_), .ZN(new_n772_));
  XOR2_X1   g571(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n773_));
  NOR3_X1   g572(.A1(new_n772_), .A2(new_n768_), .A3(new_n773_), .ZN(new_n774_));
  OR2_X1    g573(.A1(new_n767_), .A2(new_n768_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(KEYINPUT59), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n332_), .A2(new_n335_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n770_), .B1(new_n776_), .B2(new_n777_), .ZN(G1340gat));
  OAI21_X1  g577(.A(new_n462_), .B1(new_n293_), .B2(KEYINPUT60), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n769_), .B(new_n779_), .C1(KEYINPUT60), .C2(new_n462_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n776_), .A2(new_n294_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(new_n462_), .ZN(G1341gat));
  AOI21_X1  g581(.A(G127gat), .B1(new_n769_), .B2(new_n608_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n608_), .A2(G127gat), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n776_), .B2(new_n784_), .ZN(G1342gat));
  AOI21_X1  g584(.A(G134gat), .B1(new_n769_), .B2(new_n560_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n540_), .A2(G134gat), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n776_), .B2(new_n787_), .ZN(G1343gat));
  NAND3_X1  g587(.A1(new_n654_), .A2(new_n484_), .A3(new_n461_), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n767_), .A2(new_n372_), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n331_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(KEYINPUT118), .B(G141gat), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n791_), .B(new_n792_), .ZN(G1344gat));
  NAND2_X1  g592(.A1(new_n790_), .A2(new_n294_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g594(.A1(new_n790_), .A2(new_n608_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(KEYINPUT61), .B(G155gat), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n796_), .B(new_n797_), .ZN(G1346gat));
  AOI21_X1  g597(.A(G162gat), .B1(new_n790_), .B2(new_n560_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n540_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n800_), .A2(new_n528_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n799_), .B1(new_n790_), .B2(new_n801_), .ZN(G1347gat));
  INV_X1    g601(.A(KEYINPUT119), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n654_), .A2(new_n509_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n594_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n772_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n331_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n803_), .B1(new_n808_), .B2(new_n325_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n807_), .A2(KEYINPUT119), .A3(G169gat), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(KEYINPUT62), .A3(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n808_), .A2(new_n381_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT62), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n803_), .B(new_n813_), .C1(new_n808_), .C2(new_n325_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n811_), .A2(new_n812_), .A3(new_n814_), .ZN(G1348gat));
  AOI21_X1  g614(.A(G176gat), .B1(new_n806_), .B2(new_n294_), .ZN(new_n816_));
  XOR2_X1   g615(.A(new_n816_), .B(KEYINPUT120), .Z(new_n817_));
  NOR2_X1   g616(.A1(new_n767_), .A2(new_n461_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(KEYINPUT121), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n819_), .A2(G176gat), .A3(new_n294_), .A4(new_n804_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n817_), .A2(new_n820_), .ZN(G1349gat));
  INV_X1    g620(.A(new_n806_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n822_), .A2(new_n554_), .A3(new_n346_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n819_), .A2(new_n608_), .A3(new_n804_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n823_), .B1(new_n824_), .B2(new_n350_), .ZN(G1350gat));
  OAI21_X1  g624(.A(G190gat), .B1(new_n822_), .B2(new_n800_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n560_), .A2(new_n348_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT122), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n826_), .B1(new_n822_), .B2(new_n828_), .ZN(G1351gat));
  NOR4_X1   g628(.A1(new_n654_), .A2(new_n484_), .A3(new_n594_), .A4(new_n372_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n749_), .A2(KEYINPUT116), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n749_), .A2(KEYINPUT116), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n742_), .A2(new_n746_), .A3(new_n743_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n746_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n836_));
  OAI22_X1  g635(.A1(new_n833_), .A2(new_n834_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n763_), .A2(new_n765_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n554_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n710_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n831_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n331_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n294_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(G204gat), .ZN(G1353gat));
  NOR3_X1   g644(.A1(new_n767_), .A2(new_n554_), .A3(new_n831_), .ZN(new_n846_));
  XOR2_X1   g645(.A(KEYINPUT63), .B(G211gat), .Z(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT123), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  AND4_X1   g647(.A1(KEYINPUT123), .A2(new_n841_), .A3(new_n608_), .A4(new_n847_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  AOI211_X1 g650(.A(KEYINPUT124), .B(new_n851_), .C1(new_n841_), .C2(new_n608_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT124), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n763_), .A2(new_n765_), .ZN(new_n854_));
  OR2_X1    g653(.A1(new_n749_), .A2(KEYINPUT116), .ZN(new_n855_));
  AOI22_X1  g654(.A1(new_n745_), .A2(new_n747_), .B1(new_n855_), .B2(new_n832_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n608_), .B1(new_n854_), .B2(new_n856_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n608_), .B(new_n830_), .C1(new_n857_), .C2(new_n710_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n853_), .B1(new_n858_), .B2(new_n850_), .ZN(new_n859_));
  OAI22_X1  g658(.A1(new_n848_), .A2(new_n849_), .B1(new_n852_), .B2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT125), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT124), .B1(new_n846_), .B2(new_n851_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n858_), .A2(new_n853_), .A3(new_n850_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT125), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n864_), .B(new_n865_), .C1(new_n848_), .C2(new_n849_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n861_), .A2(new_n866_), .ZN(G1354gat));
  NAND2_X1  g666(.A1(new_n841_), .A2(new_n560_), .ZN(new_n868_));
  XOR2_X1   g667(.A(new_n868_), .B(KEYINPUT126), .Z(new_n869_));
  INV_X1    g668(.A(G218gat), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n800_), .A2(new_n870_), .ZN(new_n871_));
  AOI22_X1  g670(.A1(new_n869_), .A2(new_n870_), .B1(new_n841_), .B2(new_n871_), .ZN(G1355gat));
endmodule


