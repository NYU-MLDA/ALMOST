//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n791_, new_n792_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n809_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n820_, new_n821_, new_n822_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n845_, new_n846_,
    new_n847_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT6), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(KEYINPUT10), .B(G99gat), .Z(new_n206_));
  AOI21_X1  g005(.A(new_n204_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT9), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G92gat), .ZN(new_n209_));
  INV_X1    g008(.A(G85gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n208_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214_));
  AND2_X1   g013(.A1(G85gat), .A2(G92gat), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n214_), .B1(new_n215_), .B2(KEYINPUT9), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT66), .B1(new_n213_), .B2(new_n216_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n207_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT70), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT70), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n223_), .B(new_n207_), .C1(new_n219_), .C2(new_n220_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n215_), .A2(new_n214_), .ZN(new_n225_));
  OR2_X1    g024(.A1(G99gat), .A2(G106gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT7), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n225_), .B1(new_n227_), .B2(new_n204_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT8), .B1(new_n228_), .B2(KEYINPUT68), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT68), .B1(new_n228_), .B2(KEYINPUT67), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n222_), .A2(new_n224_), .A3(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(G43gat), .B(G50gat), .Z(new_n233_));
  XNOR2_X1  g032(.A(G29gat), .B(G36gat), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n234_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n237_), .B(KEYINPUT15), .Z(new_n238_));
  NAND2_X1  g037(.A1(new_n232_), .A2(new_n238_), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n221_), .A2(new_n231_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n237_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT72), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n239_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G232gat), .A2(G233gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT34), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  AOI22_X1  g046(.A1(new_n232_), .A2(new_n238_), .B1(new_n241_), .B2(new_n240_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n246_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(new_n243_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n247_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT35), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n248_), .A2(new_n252_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n247_), .A2(new_n250_), .A3(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(G190gat), .B(G218gat), .Z(new_n256_));
  XNOR2_X1  g055(.A(G134gat), .B(G162gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT36), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n253_), .A2(new_n255_), .A3(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(KEYINPUT73), .B1(new_n253_), .B2(new_n255_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n258_), .A2(new_n259_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n261_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT73), .ZN(new_n265_));
  INV_X1    g064(.A(new_n255_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT35), .B1(new_n247_), .B2(new_n250_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n265_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n263_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT37), .B1(new_n264_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n268_), .A2(new_n269_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n262_), .A2(new_n263_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT37), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .A4(new_n261_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n271_), .A2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G15gat), .B(G22gat), .ZN(new_n277_));
  INV_X1    g076(.A(G1gat), .ZN(new_n278_));
  INV_X1    g077(.A(G8gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT14), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n277_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G1gat), .B(G8gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G231gat), .A2(G233gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G57gat), .B(G64gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT11), .ZN(new_n287_));
  XOR2_X1   g086(.A(G71gat), .B(G78gat), .Z(new_n288_));
  OR2_X1    g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n286_), .A2(KEYINPUT11), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n288_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n289_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(new_n285_), .B(new_n292_), .Z(new_n293_));
  XNOR2_X1  g092(.A(G127gat), .B(G155gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT16), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G183gat), .B(G211gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT17), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n298_), .B(KEYINPUT74), .Z(new_n299_));
  NAND2_X1  g098(.A1(new_n293_), .A2(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n300_), .B(KEYINPUT75), .Z(new_n301_));
  XNOR2_X1  g100(.A(new_n297_), .B(KEYINPUT17), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n293_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n276_), .A2(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(new_n305_), .B(KEYINPUT76), .Z(new_n306_));
  NAND2_X1  g105(.A1(new_n240_), .A2(new_n292_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT12), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n240_), .A2(new_n292_), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n289_), .B(KEYINPUT12), .C1(new_n290_), .C2(new_n291_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  AOI22_X1  g110(.A1(new_n308_), .A2(new_n309_), .B1(new_n232_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G230gat), .A2(G233gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n309_), .A2(KEYINPUT69), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n240_), .A2(new_n292_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT69), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n307_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n315_), .A2(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n314_), .B1(new_n313_), .B2(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(G120gat), .B(G148gat), .Z(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT5), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G176gat), .B(G204gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n320_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT13), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT71), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n325_), .A2(KEYINPUT13), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n325_), .A2(KEYINPUT13), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n329_), .A2(KEYINPUT71), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n283_), .A2(new_n237_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n333_), .B1(new_n238_), .B2(new_n283_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G229gat), .A2(G233gat), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n283_), .B(new_n237_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n338_), .A2(new_n335_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G113gat), .B(G141gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G169gat), .B(G197gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NOR3_X1   g142(.A1(new_n337_), .A2(new_n339_), .A3(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n344_), .B(KEYINPUT78), .Z(new_n345_));
  OAI21_X1  g144(.A(new_n343_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT77), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n345_), .B(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n332_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT98), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT20), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G226gat), .A2(G233gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT19), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT23), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n355_), .A2(G183gat), .A3(G190gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT79), .ZN(new_n357_));
  INV_X1    g156(.A(G183gat), .ZN(new_n358_));
  INV_X1    g157(.A(G190gat), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT23), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT79), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n361_), .A2(new_n355_), .A3(G183gat), .A4(G190gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n357_), .A2(new_n360_), .A3(new_n362_), .ZN(new_n363_));
  OR2_X1    g162(.A1(G169gat), .A2(G176gat), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n364_), .A2(KEYINPUT24), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT80), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n363_), .A2(KEYINPUT80), .A3(new_n365_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT25), .B(G183gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT26), .B(G190gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G169gat), .A2(G176gat), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n372_), .A2(KEYINPUT24), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n370_), .A2(new_n371_), .B1(new_n373_), .B2(new_n364_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n368_), .A2(new_n369_), .A3(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT22), .B(G169gat), .ZN(new_n376_));
  INV_X1    g175(.A(G176gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n378_), .A2(KEYINPUT81), .ZN(new_n379_));
  INV_X1    g178(.A(new_n372_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n360_), .A2(new_n356_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n358_), .A2(new_n359_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n380_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n378_), .A2(KEYINPUT81), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n379_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n375_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(G204gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(G197gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(KEYINPUT89), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT89), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(G204gat), .ZN(new_n391_));
  AOI21_X1  g190(.A(G197gat), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n388_), .B1(new_n392_), .B2(KEYINPUT90), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT89), .B(G204gat), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT90), .ZN(new_n395_));
  NOR3_X1   g194(.A1(new_n394_), .A2(new_n395_), .A3(G197gat), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT21), .B1(new_n393_), .B2(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(G197gat), .A2(G204gat), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(G197gat), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n399_), .B1(new_n394_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT21), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G211gat), .B(G218gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT91), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT91), .ZN(new_n405_));
  INV_X1    g204(.A(G211gat), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n406_), .A2(G218gat), .ZN(new_n407_));
  INV_X1    g206(.A(G218gat), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n408_), .A2(G211gat), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n405_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n401_), .A2(new_n402_), .B1(new_n404_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n397_), .A2(new_n411_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n404_), .A2(new_n410_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n401_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(KEYINPUT21), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n412_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n386_), .A2(new_n416_), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n380_), .A2(KEYINPUT94), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n380_), .A2(KEYINPUT94), .ZN(new_n419_));
  AOI22_X1  g218(.A1(new_n418_), .A2(new_n419_), .B1(new_n377_), .B2(new_n376_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n363_), .A2(KEYINPUT95), .A3(new_n382_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(KEYINPUT95), .B1(new_n363_), .B2(new_n382_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n420_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n365_), .A2(new_n381_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(new_n374_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n413_), .A2(KEYINPUT21), .ZN(new_n428_));
  AOI22_X1  g227(.A1(new_n428_), .A2(new_n414_), .B1(new_n397_), .B2(new_n411_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  AOI211_X1 g229(.A(new_n352_), .B(new_n354_), .C1(new_n417_), .C2(new_n430_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n375_), .A2(new_n412_), .A3(new_n385_), .A4(new_n415_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n363_), .A2(new_n382_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT95), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n421_), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n436_), .A2(new_n420_), .B1(new_n374_), .B2(new_n425_), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n432_), .B(KEYINPUT20), .C1(new_n437_), .C2(new_n429_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n354_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT96), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n438_), .A2(KEYINPUT96), .A3(new_n354_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n431_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G8gat), .B(G36gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT18), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G64gat), .B(G92gat), .ZN(new_n446_));
  XOR2_X1   g245(.A(new_n445_), .B(new_n446_), .Z(new_n447_));
  OAI21_X1  g246(.A(new_n351_), .B1(new_n443_), .B2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n352_), .B1(new_n417_), .B2(new_n430_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n354_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n438_), .A2(KEYINPUT96), .A3(new_n354_), .ZN(new_n452_));
  AOI21_X1  g251(.A(KEYINPUT96), .B1(new_n438_), .B2(new_n354_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n451_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n447_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(KEYINPUT98), .A3(new_n455_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n451_), .B(new_n447_), .C1(new_n452_), .C2(new_n453_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT97), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n441_), .A2(new_n442_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT97), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n459_), .A2(new_n460_), .A3(new_n451_), .A4(new_n447_), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n448_), .A2(new_n456_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n462_), .A2(KEYINPUT27), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n438_), .A2(new_n450_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n464_), .B1(new_n449_), .B2(new_n354_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(new_n455_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(KEYINPUT27), .A3(new_n457_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n463_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G155gat), .A2(G162gat), .ZN(new_n469_));
  OR2_X1    g268(.A1(G155gat), .A2(G162gat), .ZN(new_n470_));
  NOR2_X1   g269(.A1(G141gat), .A2(G148gat), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT3), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G141gat), .A2(G148gat), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT2), .ZN(new_n474_));
  AOI22_X1  g273(.A1(new_n471_), .A2(new_n472_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n475_), .B1(new_n472_), .B2(new_n471_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT87), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n469_), .B(new_n470_), .C1(new_n476_), .C2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT88), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n469_), .A2(KEYINPUT85), .A3(KEYINPUT1), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n470_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT86), .ZN(new_n484_));
  AOI21_X1  g283(.A(KEYINPUT85), .B1(new_n469_), .B2(KEYINPUT1), .ZN(new_n485_));
  OR3_X1    g284(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n484_), .B1(new_n483_), .B2(new_n485_), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n486_), .B(new_n487_), .C1(KEYINPUT1), .C2(new_n469_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n471_), .B(KEYINPUT84), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(new_n473_), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n481_), .A2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n429_), .B1(new_n491_), .B2(KEYINPUT29), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G228gat), .A2(G233gat), .ZN(new_n493_));
  XOR2_X1   g292(.A(new_n492_), .B(new_n493_), .Z(new_n494_));
  XOR2_X1   g293(.A(G78gat), .B(G106gat), .Z(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT92), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT93), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n491_), .A2(KEYINPUT29), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT28), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G22gat), .B(G50gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n498_), .A2(new_n502_), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n494_), .A2(new_n496_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n503_), .A2(new_n497_), .A3(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n497_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n506_), .A2(new_n502_), .A3(new_n498_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n468_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n386_), .B(KEYINPUT30), .ZN(new_n511_));
  XOR2_X1   g310(.A(G71gat), .B(G99gat), .Z(new_n512_));
  NAND2_X1  g311(.A1(G227gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G15gat), .B(G43gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT82), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n514_), .B(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n511_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT31), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G127gat), .B(G134gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT83), .ZN(new_n521_));
  XOR2_X1   g320(.A(G113gat), .B(G120gat), .Z(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n519_), .A2(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n519_), .A2(new_n523_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n523_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n491_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n481_), .A2(new_n490_), .A3(new_n523_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G225gat), .A2(G233gat), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n528_), .A2(KEYINPUT4), .A3(new_n529_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n530_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n533_), .B1(new_n528_), .B2(KEYINPUT4), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n531_), .B1(new_n532_), .B2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G1gat), .B(G29gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT0), .ZN(new_n537_));
  INV_X1    g336(.A(G57gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(G85gat), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n535_), .A2(new_n541_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n531_), .B(new_n540_), .C1(new_n532_), .C2(new_n534_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n526_), .A2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n510_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n468_), .A2(new_n545_), .A3(new_n508_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n447_), .A2(KEYINPUT32), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n542_), .A2(new_n543_), .B1(new_n550_), .B2(new_n465_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n459_), .A2(new_n451_), .A3(new_n549_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n552_), .A2(KEYINPUT101), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(KEYINPUT101), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n551_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT102), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n551_), .B(KEYINPUT102), .C1(new_n553_), .C2(new_n554_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT100), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT33), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n543_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n528_), .A2(KEYINPUT4), .A3(new_n529_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n563_), .B(new_n533_), .C1(KEYINPUT4), .C2(new_n528_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n564_), .A2(KEYINPUT33), .A3(new_n531_), .A4(new_n540_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n528_), .A2(new_n529_), .A3(new_n533_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n530_), .B1(new_n528_), .B2(KEYINPUT4), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n541_), .B(new_n566_), .C1(new_n532_), .C2(new_n567_), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n562_), .A2(new_n565_), .A3(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n569_), .B1(new_n462_), .B2(KEYINPUT99), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n448_), .A2(new_n456_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n458_), .A2(new_n461_), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n571_), .A2(KEYINPUT99), .A3(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n560_), .B1(new_n570_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n571_), .A2(new_n572_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT99), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n462_), .A2(KEYINPUT99), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n577_), .A2(KEYINPUT100), .A3(new_n578_), .A4(new_n569_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n559_), .B1(new_n574_), .B2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n548_), .B1(new_n580_), .B2(new_n508_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n526_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n547_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n350_), .A2(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n306_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n586_), .A2(new_n278_), .A3(new_n544_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT38), .ZN(new_n588_));
  INV_X1    g387(.A(new_n304_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n350_), .A2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n264_), .A2(new_n270_), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n591_), .B(KEYINPUT103), .Z(new_n592_));
  NAND2_X1  g391(.A1(new_n584_), .A2(new_n592_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n590_), .A2(new_n545_), .A3(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n588_), .B1(new_n278_), .B2(new_n594_), .ZN(G1324gat));
  INV_X1    g394(.A(new_n468_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n586_), .A2(new_n279_), .A3(new_n596_), .ZN(new_n597_));
  NOR3_X1   g396(.A1(new_n590_), .A2(new_n468_), .A3(new_n593_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT104), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT39), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n279_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n600_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n601_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n597_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT40), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  OAI211_X1 g406(.A(KEYINPUT40), .B(new_n597_), .C1(new_n603_), .C2(new_n604_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(G1325gat));
  NOR2_X1   g408(.A1(new_n590_), .A2(new_n593_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(new_n526_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(G15gat), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n612_), .A2(KEYINPUT41), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(KEYINPUT41), .ZN(new_n614_));
  INV_X1    g413(.A(G15gat), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n586_), .A2(new_n615_), .A3(new_n526_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n613_), .A2(new_n614_), .A3(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT105), .ZN(G1326gat));
  INV_X1    g417(.A(G22gat), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n619_), .B1(new_n610_), .B2(new_n508_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT42), .Z(new_n621_));
  NAND2_X1  g420(.A1(new_n508_), .A2(new_n619_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT106), .Z(new_n623_));
  NAND2_X1  g422(.A1(new_n586_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n621_), .A2(new_n624_), .ZN(G1327gat));
  NOR2_X1   g424(.A1(new_n591_), .A2(new_n589_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n585_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(G29gat), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(new_n629_), .A3(new_n544_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT44), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n271_), .A2(new_n275_), .ZN(new_n632_));
  NOR4_X1   g431(.A1(new_n583_), .A2(new_n632_), .A3(KEYINPUT107), .A4(KEYINPUT43), .ZN(new_n633_));
  OAI21_X1  g432(.A(KEYINPUT43), .B1(new_n583_), .B2(new_n632_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT107), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  OR3_X1    g435(.A1(new_n583_), .A2(KEYINPUT43), .A3(new_n632_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n633_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n350_), .A2(new_n304_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n631_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n639_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n583_), .A2(KEYINPUT43), .A3(new_n632_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n642_), .B1(new_n635_), .B2(new_n634_), .ZN(new_n643_));
  OAI211_X1 g442(.A(KEYINPUT44), .B(new_n641_), .C1(new_n643_), .C2(new_n633_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n640_), .A2(KEYINPUT108), .A3(new_n644_), .A4(new_n544_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n645_), .A2(G29gat), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n640_), .A2(new_n544_), .A3(new_n644_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT108), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT109), .B1(new_n646_), .B2(new_n649_), .ZN(new_n650_));
  AND4_X1   g449(.A1(KEYINPUT109), .A2(new_n649_), .A3(G29gat), .A4(new_n645_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n630_), .B1(new_n650_), .B2(new_n651_), .ZN(G1328gat));
  XOR2_X1   g451(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n468_), .A2(G36gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n654_), .B1(new_n628_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n655_), .ZN(new_n657_));
  NOR4_X1   g456(.A1(new_n585_), .A2(new_n627_), .A3(new_n657_), .A4(new_n653_), .ZN(new_n658_));
  OAI22_X1  g457(.A1(new_n656_), .A2(new_n658_), .B1(KEYINPUT111), .B2(KEYINPUT46), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n640_), .A2(new_n596_), .A3(new_n644_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(G36gat), .B2(new_n660_), .ZN(new_n661_));
  AND2_X1   g460(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(G1329gat));
  INV_X1    g462(.A(G43gat), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n628_), .A2(new_n664_), .A3(new_n526_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n640_), .A2(new_n526_), .A3(new_n644_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n666_), .B2(new_n664_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT47), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(G1330gat));
  INV_X1    g468(.A(G50gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n628_), .A2(new_n670_), .A3(new_n508_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n640_), .A2(new_n508_), .A3(new_n644_), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n672_), .A2(KEYINPUT112), .A3(G50gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(KEYINPUT112), .B1(new_n672_), .B2(G50gat), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n671_), .B1(new_n673_), .B2(new_n674_), .ZN(G1331gat));
  NAND2_X1  g474(.A1(new_n332_), .A2(new_n349_), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n306_), .A2(new_n583_), .A3(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n677_), .A2(new_n538_), .A3(new_n544_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n593_), .A2(new_n676_), .A3(new_n304_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G57gat), .B1(new_n680_), .B2(new_n545_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n678_), .A2(new_n681_), .ZN(G1332gat));
  INV_X1    g481(.A(G64gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n683_), .B1(new_n679_), .B2(new_n596_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  XOR2_X1   g484(.A(KEYINPUT113), .B(KEYINPUT48), .Z(new_n686_));
  OR2_X1    g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n686_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n677_), .A2(new_n683_), .A3(new_n596_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n687_), .A2(new_n688_), .A3(new_n689_), .ZN(G1333gat));
  INV_X1    g489(.A(G71gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n691_), .B1(new_n679_), .B2(new_n526_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT49), .Z(new_n693_));
  NAND3_X1  g492(.A1(new_n677_), .A2(new_n691_), .A3(new_n526_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1334gat));
  INV_X1    g494(.A(G78gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n696_), .B1(new_n679_), .B2(new_n508_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT50), .Z(new_n698_));
  NAND3_X1  g497(.A1(new_n677_), .A2(new_n696_), .A3(new_n508_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1335gat));
  NOR3_X1   g499(.A1(new_n676_), .A2(new_n583_), .A3(new_n627_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n701_), .A2(new_n210_), .A3(new_n544_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n676_), .A2(new_n589_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n638_), .A2(new_n545_), .A3(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n702_), .B1(new_n705_), .B2(new_n210_), .ZN(G1336gat));
  AOI21_X1  g505(.A(G92gat), .B1(new_n701_), .B2(new_n596_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n638_), .A2(new_n704_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n468_), .A2(new_n209_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n707_), .B1(new_n708_), .B2(new_n709_), .ZN(G1337gat));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n526_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n526_), .A2(new_n206_), .ZN(new_n712_));
  AOI22_X1  g511(.A1(new_n711_), .A2(G99gat), .B1(new_n701_), .B2(new_n712_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT51), .Z(G1338gat));
  XNOR2_X1  g513(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n508_), .B(new_n703_), .C1(new_n643_), .C2(new_n633_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(G106gat), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT52), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n701_), .A2(new_n205_), .A3(new_n508_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n715_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n717_), .A2(KEYINPUT52), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT52), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(new_n716_), .B2(G106gat), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n719_), .B(new_n715_), .C1(new_n721_), .C2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n720_), .A2(new_n725_), .ZN(G1339gat));
  NAND3_X1  g525(.A1(new_n305_), .A2(new_n349_), .A3(new_n326_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT54), .Z(new_n728_));
  OR2_X1    g527(.A1(new_n320_), .A2(new_n324_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(new_n348_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT115), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT55), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n314_), .A2(new_n731_), .A3(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n733_), .B1(new_n313_), .B2(new_n312_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n732_), .B1(new_n314_), .B2(new_n731_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n324_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT56), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  OAI211_X1 g537(.A(KEYINPUT56), .B(new_n324_), .C1(new_n734_), .C2(new_n735_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n730_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n343_), .B1(new_n338_), .B2(new_n335_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT116), .ZN(new_n742_));
  AOI22_X1  g541(.A1(new_n334_), .A2(new_n336_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n743_), .B1(new_n742_), .B2(new_n741_), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n325_), .A2(new_n346_), .A3(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n591_), .B1(new_n740_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT57), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT57), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n748_), .B(new_n591_), .C1(new_n740_), .C2(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n735_), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n751_), .B(new_n733_), .C1(new_n313_), .C2(new_n312_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n752_), .A2(KEYINPUT117), .A3(KEYINPUT56), .A4(new_n324_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT117), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n739_), .A2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n753_), .A2(new_n755_), .A3(new_n738_), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n729_), .A2(new_n346_), .A3(new_n744_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT58), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n756_), .A2(KEYINPUT58), .A3(new_n757_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(new_n276_), .A3(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n589_), .B1(new_n750_), .B2(new_n762_), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n728_), .A2(new_n763_), .ZN(new_n764_));
  NOR3_X1   g563(.A1(new_n510_), .A2(new_n545_), .A3(new_n582_), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT119), .Z(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT120), .Z(new_n767_));
  NOR2_X1   g566(.A1(new_n767_), .A2(KEYINPUT59), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n764_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n766_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n750_), .A2(new_n762_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT118), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n750_), .A2(new_n762_), .A3(KEYINPUT118), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n304_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n728_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n770_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT59), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n769_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(G113gat), .B1(new_n780_), .B2(new_n349_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n778_), .ZN(new_n782_));
  OR3_X1    g581(.A1(new_n782_), .A2(G113gat), .A3(new_n349_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(G1340gat));
  INV_X1    g583(.A(new_n332_), .ZN(new_n785_));
  OAI21_X1  g584(.A(G120gat), .B1(new_n780_), .B2(new_n785_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n785_), .A2(KEYINPUT60), .A3(G120gat), .ZN(new_n787_));
  AND2_X1   g586(.A1(KEYINPUT60), .A2(G120gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n778_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n786_), .A2(new_n789_), .ZN(G1341gat));
  OAI21_X1  g589(.A(G127gat), .B1(new_n780_), .B2(new_n304_), .ZN(new_n791_));
  OR3_X1    g590(.A1(new_n782_), .A2(G127gat), .A3(new_n304_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(G1342gat));
  INV_X1    g592(.A(new_n592_), .ZN(new_n794_));
  AOI21_X1  g593(.A(G134gat), .B1(new_n778_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n780_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(KEYINPUT121), .B(G134gat), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n632_), .A2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n795_), .B1(new_n796_), .B2(new_n798_), .ZN(G1343gat));
  AOI21_X1  g598(.A(new_n589_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n800_), .A2(new_n728_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n596_), .A2(new_n509_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n803_), .A2(new_n545_), .A3(new_n526_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n801_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n348_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n332_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g609(.A1(new_n776_), .A2(new_n777_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT122), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n589_), .A4(new_n804_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n589_), .B(new_n804_), .C1(new_n800_), .C2(new_n728_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT122), .ZN(new_n815_));
  XOR2_X1   g614(.A(KEYINPUT61), .B(G155gat), .Z(new_n816_));
  AND3_X1   g615(.A1(new_n813_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n816_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(G1346gat));
  INV_X1    g618(.A(G162gat), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n806_), .A2(new_n820_), .A3(new_n794_), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n801_), .A2(new_n632_), .A3(new_n805_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n820_), .B2(new_n822_), .ZN(G1347gat));
  NOR2_X1   g622(.A1(new_n468_), .A2(new_n546_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n509_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n764_), .A2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n827_), .A2(new_n376_), .A3(new_n348_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n824_), .A2(new_n348_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT123), .ZN(new_n830_));
  OR2_X1    g629(.A1(new_n829_), .A2(KEYINPUT123), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n764_), .A2(new_n509_), .A3(new_n830_), .A4(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT62), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n832_), .A2(new_n833_), .A3(G169gat), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n832_), .B2(G169gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n828_), .B1(new_n834_), .B2(new_n835_), .ZN(G1348gat));
  OAI211_X1 g635(.A(new_n332_), .B(new_n826_), .C1(new_n728_), .C2(new_n763_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n377_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n332_), .A2(G176gat), .A3(new_n509_), .A4(new_n824_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n801_), .B2(new_n839_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(KEYINPUT124), .ZN(G1349gat));
  NAND2_X1  g640(.A1(new_n827_), .A2(new_n589_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n842_), .A2(new_n370_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n843_), .B1(new_n358_), .B2(new_n842_), .ZN(G1350gat));
  NAND3_X1  g643(.A1(new_n827_), .A2(new_n371_), .A3(new_n794_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n827_), .A2(new_n276_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n845_), .B1(new_n847_), .B2(new_n359_), .ZN(G1351gat));
  NOR4_X1   g647(.A1(new_n468_), .A2(new_n509_), .A3(new_n544_), .A4(new_n526_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n811_), .A2(new_n849_), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n850_), .A2(G197gat), .A3(new_n348_), .ZN(new_n851_));
  AOI21_X1  g650(.A(G197gat), .B1(new_n850_), .B2(new_n348_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1352gat));
  INV_X1    g652(.A(KEYINPUT125), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n850_), .A2(new_n854_), .A3(new_n394_), .A4(new_n332_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n811_), .A2(new_n332_), .A3(new_n849_), .ZN(new_n856_));
  AOI21_X1  g655(.A(KEYINPUT125), .B1(new_n856_), .B2(G204gat), .ZN(new_n857_));
  INV_X1    g656(.A(new_n394_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n856_), .A2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n855_), .B1(new_n857_), .B2(new_n859_), .ZN(G1353gat));
  OR2_X1    g659(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n304_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT126), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n850_), .A2(new_n861_), .A3(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n861_), .B1(new_n850_), .B2(new_n863_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n864_), .A2(new_n865_), .ZN(G1354gat));
  NAND2_X1  g665(.A1(new_n850_), .A2(new_n794_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n276_), .A2(G218gat), .ZN(new_n868_));
  XOR2_X1   g667(.A(new_n868_), .B(KEYINPUT127), .Z(new_n869_));
  AOI22_X1  g668(.A1(new_n867_), .A2(new_n408_), .B1(new_n850_), .B2(new_n869_), .ZN(G1355gat));
endmodule


