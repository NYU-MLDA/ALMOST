//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n786_, new_n787_, new_n788_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n800_, new_n801_, new_n802_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n907_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n949_, new_n950_, new_n951_, new_n953_, new_n954_,
    new_n956_, new_n957_, new_n958_, new_n960_, new_n962_, new_n963_,
    new_n964_, new_n966_, new_n967_, new_n968_;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  INV_X1    g001(.A(G176gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT88), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT88), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G176gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT22), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n207_), .A2(G169gat), .ZN(new_n208_));
  OAI211_X1 g007(.A(new_n204_), .B(new_n206_), .C1(new_n208_), .C2(KEYINPUT87), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT87), .ZN(new_n210_));
  INV_X1    g009(.A(G169gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT22), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n207_), .A2(G169gat), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n210_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n202_), .B1(new_n209_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT89), .ZN(new_n216_));
  INV_X1    g015(.A(G183gat), .ZN(new_n217_));
  INV_X1    g016(.A(G190gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT23), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT23), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(G183gat), .A3(G190gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n217_), .A2(new_n218_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n216_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n215_), .A2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n222_), .A2(new_n216_), .A3(new_n223_), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n221_), .A2(KEYINPUT86), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n221_), .A2(KEYINPUT86), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n219_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n211_), .A2(new_n203_), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n230_), .A2(KEYINPUT24), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n217_), .A2(KEYINPUT25), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT25), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(G183gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n218_), .A2(KEYINPUT26), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT26), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(G190gat), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n232_), .A2(new_n234_), .A3(new_n235_), .A4(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n230_), .A2(KEYINPUT24), .A3(new_n202_), .ZN(new_n239_));
  AND3_X1   g038(.A1(new_n231_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  AOI22_X1  g039(.A1(new_n225_), .A2(new_n226_), .B1(new_n229_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G227gat), .A2(G233gat), .ZN(new_n242_));
  XOR2_X1   g041(.A(new_n242_), .B(G15gat), .Z(new_n243_));
  XNOR2_X1  g042(.A(new_n241_), .B(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT31), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n245_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G71gat), .B(G99gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(G43gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT90), .B(KEYINPUT30), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G127gat), .B(G134gat), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(G113gat), .B(G120gat), .Z(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT91), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G113gat), .B(G120gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT92), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n253_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n258_), .B1(new_n253_), .B2(new_n257_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n256_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n253_), .A2(new_n257_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT92), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n253_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT91), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n265_), .B1(new_n253_), .B2(new_n257_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n263_), .A2(new_n264_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n261_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n252_), .B(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n248_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n246_), .A2(new_n247_), .A3(new_n269_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G1gat), .B(G29gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(G85gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT0), .B(G57gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT2), .ZN(new_n279_));
  INV_X1    g078(.A(G141gat), .ZN(new_n280_));
  INV_X1    g079(.A(G148gat), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n279_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT3), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n283_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n282_), .A2(new_n284_), .A3(new_n285_), .A4(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G155gat), .A2(G162gat), .ZN(new_n288_));
  OR2_X1    g087(.A1(G155gat), .A2(G162gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(G141gat), .B(G148gat), .Z(new_n291_));
  NAND2_X1  g090(.A1(new_n288_), .A2(KEYINPUT1), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(new_n289_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n288_), .A2(KEYINPUT1), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n291_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n290_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n261_), .A2(new_n296_), .A3(new_n267_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT4), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n262_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n253_), .A2(new_n257_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n290_), .B(new_n295_), .C1(new_n301_), .C2(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n298_), .B1(new_n297_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G225gat), .A2(G233gat), .ZN(new_n305_));
  NOR3_X1   g104(.A1(new_n300_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n297_), .A2(new_n303_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n305_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n278_), .B1(new_n306_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT103), .ZN(new_n311_));
  INV_X1    g110(.A(new_n304_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n305_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n312_), .A2(new_n313_), .A3(new_n299_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(new_n277_), .A3(new_n308_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n310_), .A2(new_n311_), .A3(new_n315_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n314_), .A2(KEYINPUT103), .A3(new_n277_), .A4(new_n308_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n273_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G78gat), .B(G106gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  AND2_X1   g120(.A1(G228gat), .A2(G233gat), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(G211gat), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n324_), .A2(G218gat), .ZN(new_n325_));
  INV_X1    g124(.A(G218gat), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n326_), .A2(G211gat), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT95), .B1(new_n325_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(G211gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n324_), .A2(G218gat), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT95), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n329_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n328_), .A2(new_n332_), .ZN(new_n333_));
  XOR2_X1   g132(.A(G197gat), .B(G204gat), .Z(new_n334_));
  NAND3_X1  g133(.A1(new_n334_), .A2(KEYINPUT94), .A3(KEYINPUT21), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT94), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G197gat), .B(G204gat), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT21), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n337_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n338_), .A2(new_n339_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n336_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT96), .ZN(new_n344_));
  AND3_X1   g143(.A1(new_n329_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n331_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n344_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n328_), .A2(KEYINPUT96), .A3(new_n332_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n347_), .A2(new_n348_), .A3(new_n341_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT97), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n347_), .A2(new_n348_), .A3(KEYINPUT97), .A4(new_n341_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n343_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT93), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n323_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n290_), .A2(new_n295_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT29), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n353_), .A2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n355_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n351_), .A2(new_n352_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n343_), .ZN(new_n362_));
  AOI221_X4 g161(.A(new_n358_), .B1(new_n354_), .B2(new_n323_), .C1(new_n361_), .C2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n321_), .B1(new_n360_), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n334_), .A2(KEYINPUT21), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n365_), .B1(new_n333_), .B2(new_n344_), .ZN(new_n366_));
  AOI21_X1  g165(.A(KEYINPUT97), .B1(new_n366_), .B2(new_n348_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n352_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n362_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n358_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(KEYINPUT93), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(new_n372_), .A3(new_n323_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n355_), .A2(new_n359_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(new_n374_), .A3(new_n320_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n364_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n356_), .A2(new_n357_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT28), .ZN(new_n378_));
  XOR2_X1   g177(.A(G22gat), .B(G50gat), .Z(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n376_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n375_), .A2(KEYINPUT98), .ZN(new_n382_));
  OAI211_X1 g181(.A(KEYINPUT99), .B(new_n321_), .C1(new_n360_), .C2(new_n363_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT98), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n373_), .A2(new_n374_), .A3(new_n384_), .A4(new_n320_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n382_), .A2(new_n383_), .A3(new_n385_), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n378_), .B(new_n379_), .Z(new_n387_));
  AOI21_X1  g186(.A(new_n320_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n387_), .B1(new_n388_), .B2(KEYINPUT99), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n381_), .B1(new_n386_), .B2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G8gat), .B(G36gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT18), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G64gat), .B(G92gat), .ZN(new_n393_));
  XOR2_X1   g192(.A(new_n392_), .B(new_n393_), .Z(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT20), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n396_), .B1(new_n353_), .B2(new_n241_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G226gat), .A2(G233gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT19), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n229_), .A2(new_n223_), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n204_), .A2(new_n206_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n212_), .A2(new_n213_), .ZN(new_n403_));
  AOI22_X1  g202(.A1(new_n402_), .A2(new_n403_), .B1(G169gat), .B2(G176gat), .ZN(new_n404_));
  AOI22_X1  g203(.A1(new_n401_), .A2(new_n404_), .B1(new_n240_), .B2(new_n222_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n369_), .A2(new_n406_), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n397_), .A2(new_n400_), .A3(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n396_), .B1(new_n353_), .B2(new_n405_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n225_), .A2(new_n226_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n240_), .A2(new_n229_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n369_), .A2(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n400_), .B1(new_n409_), .B2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n395_), .B1(new_n408_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT104), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n362_), .B(new_n405_), .C1(new_n367_), .C2(new_n368_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT20), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n353_), .A2(new_n241_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n399_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n397_), .A2(new_n400_), .A3(new_n407_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT104), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(new_n423_), .A3(new_n395_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n416_), .A2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT20), .B1(new_n369_), .B2(new_n412_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n353_), .A2(new_n405_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n399_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n409_), .A2(new_n400_), .A3(new_n413_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(KEYINPUT100), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT100), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n409_), .A2(new_n413_), .A3(new_n431_), .A4(new_n400_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n395_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT27), .B1(new_n425_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n429_), .A2(KEYINPUT100), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n400_), .B1(new_n397_), .B2(new_n407_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n432_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(new_n394_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT27), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n430_), .A2(new_n395_), .A3(new_n432_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  AOI211_X1 g240(.A(new_n319_), .B(new_n390_), .C1(new_n434_), .C2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n387_), .B1(new_n364_), .B2(new_n375_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n382_), .A2(new_n383_), .A3(new_n385_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT99), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n380_), .B1(new_n364_), .B2(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n443_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n437_), .A2(new_n394_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT101), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n449_), .A2(KEYINPUT33), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n310_), .A2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n305_), .B1(new_n300_), .B2(new_n304_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT102), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  OAI211_X1 g253(.A(KEYINPUT102), .B(new_n305_), .C1(new_n300_), .C2(new_n304_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n297_), .A2(new_n303_), .A3(new_n313_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n454_), .A2(new_n277_), .A3(new_n455_), .A4(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n450_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n278_), .B(new_n458_), .C1(new_n306_), .C2(new_n309_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n451_), .A2(new_n457_), .A3(new_n459_), .ZN(new_n460_));
  NOR3_X1   g259(.A1(new_n448_), .A2(new_n433_), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n394_), .A2(KEYINPUT32), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n422_), .A2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n464_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n463_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n447_), .B1(new_n461_), .B2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n423_), .B1(new_n422_), .B2(new_n395_), .ZN(new_n469_));
  AOI211_X1 g268(.A(KEYINPUT104), .B(new_n394_), .C1(new_n420_), .C2(new_n421_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n439_), .B1(new_n471_), .B2(new_n438_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n438_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n390_), .A2(new_n318_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n468_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n273_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n442_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G230gat), .A2(G233gat), .ZN(new_n479_));
  XOR2_X1   g278(.A(new_n479_), .B(KEYINPUT64), .Z(new_n480_));
  INV_X1    g279(.A(G85gat), .ZN(new_n481_));
  INV_X1    g280(.A(G92gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT9), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G85gat), .A2(G92gat), .ZN(new_n485_));
  AND3_X1   g284(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  AOI22_X1  g286(.A1(new_n483_), .A2(new_n485_), .B1(new_n484_), .B2(G92gat), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n489_), .A3(KEYINPUT65), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G99gat), .A2(G106gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT6), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT6), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n493_), .A2(G99gat), .A3(G106gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT66), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n492_), .A2(new_n494_), .A3(KEYINPUT66), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  XOR2_X1   g298(.A(KEYINPUT10), .B(G99gat), .Z(new_n500_));
  INV_X1    g299(.A(G106gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT65), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n503_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n490_), .A2(new_n499_), .A3(new_n502_), .A4(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G57gat), .B(G64gat), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n506_), .A2(KEYINPUT11), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(KEYINPUT11), .ZN(new_n508_));
  XOR2_X1   g307(.A(G71gat), .B(G78gat), .Z(new_n509_));
  NAND3_X1  g308(.A1(new_n507_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n508_), .A2(new_n509_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT7), .ZN(new_n513_));
  INV_X1    g312(.A(G99gat), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(new_n514_), .A3(new_n501_), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n497_), .A2(new_n498_), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT8), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n483_), .A2(new_n485_), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n515_), .A2(new_n516_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT67), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT67), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n515_), .A2(new_n524_), .A3(new_n516_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(new_n495_), .A3(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n519_), .B1(new_n526_), .B2(new_n520_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n505_), .B(new_n512_), .C1(new_n521_), .C2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT12), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n520_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT8), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n512_), .B1(new_n533_), .B2(new_n505_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n529_), .A2(new_n534_), .ZN(new_n535_));
  AOI211_X1 g334(.A(KEYINPUT12), .B(new_n512_), .C1(new_n533_), .C2(new_n505_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n480_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT69), .ZN(new_n538_));
  INV_X1    g337(.A(new_n480_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n512_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n521_), .A2(new_n527_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n505_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n540_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n543_), .A2(KEYINPUT12), .A3(new_n528_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n533_), .A2(new_n505_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT12), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n545_), .A2(new_n546_), .A3(new_n540_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n539_), .B1(new_n544_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT69), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  OR3_X1    g349(.A1(new_n545_), .A2(KEYINPUT68), .A3(new_n540_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n543_), .A2(KEYINPUT68), .A3(new_n528_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(new_n539_), .A3(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n538_), .A2(new_n550_), .A3(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(G120gat), .B(G148gat), .Z(new_n555_));
  XNOR2_X1  g354(.A(G176gat), .B(G204gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n560_), .A2(KEYINPUT70), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT72), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n554_), .B(new_n562_), .Z(new_n563_));
  INV_X1    g362(.A(KEYINPUT13), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n554_), .B(new_n562_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(KEYINPUT13), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G29gat), .B(G36gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G43gat), .B(G50gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT73), .B(KEYINPUT15), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G15gat), .B(G22gat), .ZN(new_n574_));
  INV_X1    g373(.A(G1gat), .ZN(new_n575_));
  INV_X1    g374(.A(G8gat), .ZN(new_n576_));
  OAI21_X1  g375(.A(KEYINPUT14), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n574_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G1gat), .B(G8gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n573_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT84), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G229gat), .A2(G233gat), .ZN(new_n583_));
  INV_X1    g382(.A(new_n580_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(new_n571_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT84), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n573_), .A2(new_n586_), .A3(new_n580_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n582_), .A2(new_n583_), .A3(new_n585_), .A4(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT83), .ZN(new_n589_));
  INV_X1    g388(.A(new_n585_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n584_), .A2(new_n571_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n589_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n584_), .A2(new_n571_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n593_), .A2(KEYINPUT83), .A3(new_n585_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n588_), .B1(new_n595_), .B2(new_n583_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G113gat), .B(G141gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G169gat), .B(G197gat), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n597_), .B(new_n598_), .Z(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n596_), .A2(new_n600_), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n588_), .B(new_n599_), .C1(new_n595_), .C2(new_n583_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT85), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n478_), .A2(new_n568_), .A3(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT37), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G190gat), .B(G218gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G134gat), .B(G162gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n609_), .B(KEYINPUT36), .Z(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT76), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G232gat), .A2(G233gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT34), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n614_), .A2(KEYINPUT35), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n545_), .A2(new_n573_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT74), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n541_), .A2(new_n542_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n571_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n616_), .A2(new_n617_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n615_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n614_), .A2(KEYINPUT35), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n615_), .A2(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n620_), .A2(new_n616_), .A3(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT75), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n620_), .A2(new_n616_), .A3(KEYINPUT75), .A4(new_n625_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n612_), .B1(new_n623_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n609_), .A2(KEYINPUT36), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n623_), .A2(new_n630_), .A3(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n606_), .B1(new_n632_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n634_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n610_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n637_), .B1(new_n623_), .B2(new_n630_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n636_), .A2(new_n638_), .A3(KEYINPUT37), .ZN(new_n639_));
  OAI21_X1  g438(.A(KEYINPUT77), .B1(new_n635_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n638_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n641_), .A2(new_n606_), .A3(new_n634_), .ZN(new_n642_));
  OAI21_X1  g441(.A(KEYINPUT37), .B1(new_n636_), .B2(new_n631_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT77), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n642_), .A2(new_n643_), .A3(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n640_), .A2(new_n645_), .ZN(new_n646_));
  XOR2_X1   g445(.A(G127gat), .B(G155gat), .Z(new_n647_));
  XNOR2_X1  g446(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(G183gat), .B(G211gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT17), .Z(new_n652_));
  NAND2_X1  g451(.A1(G231gat), .A2(G233gat), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n580_), .B(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(new_n512_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n652_), .A2(new_n655_), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n656_), .A2(KEYINPUT81), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n655_), .A2(KEYINPUT78), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n655_), .A2(KEYINPUT78), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT80), .B(KEYINPUT17), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n658_), .A2(new_n659_), .A3(new_n651_), .A4(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n656_), .A2(KEYINPUT81), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n657_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT82), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n663_), .B(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n646_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n605_), .A2(new_n666_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT105), .Z(new_n668_));
  INV_X1    g467(.A(new_n318_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(new_n575_), .A3(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT38), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n671_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n565_), .A2(new_n567_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(new_n603_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n675_), .A2(new_n663_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n636_), .A2(new_n638_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n478_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(G1gat), .B1(new_n679_), .B2(new_n318_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n672_), .A2(new_n673_), .A3(new_n680_), .ZN(G1324gat));
  NAND3_X1  g480(.A1(new_n668_), .A2(new_n576_), .A3(new_n474_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n676_), .A2(new_n474_), .A3(new_n678_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(G8gat), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n684_), .A2(KEYINPUT39), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n684_), .A2(KEYINPUT39), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n682_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT40), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OAI211_X1 g488(.A(new_n682_), .B(KEYINPUT40), .C1(new_n686_), .C2(new_n685_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1325gat));
  OAI21_X1  g490(.A(G15gat), .B1(new_n679_), .B2(new_n477_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT41), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n667_), .A2(G15gat), .A3(new_n477_), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1326gat));
  OAI21_X1  g494(.A(G22gat), .B1(new_n679_), .B2(new_n447_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT42), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n447_), .A2(G22gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n697_), .B1(new_n667_), .B2(new_n698_), .ZN(G1327gat));
  INV_X1    g498(.A(new_n665_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n677_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n605_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(G29gat), .B1(new_n704_), .B2(new_n669_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n674_), .A2(new_n665_), .A3(new_n603_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n446_), .A2(new_n383_), .A3(new_n382_), .A4(new_n385_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n669_), .B1(new_n709_), .B2(new_n381_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n710_), .B1(new_n473_), .B2(new_n472_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n273_), .B1(new_n711_), .B2(new_n468_), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n646_), .B(new_n708_), .C1(new_n712_), .C2(new_n442_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n434_), .A2(new_n441_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n319_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n715_), .A2(new_n447_), .A3(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n438_), .A2(new_n440_), .ZN(new_n718_));
  OAI22_X1  g517(.A1(new_n718_), .A2(new_n460_), .B1(new_n466_), .B2(new_n465_), .ZN(new_n719_));
  AOI22_X1  g518(.A1(new_n715_), .A2(new_n710_), .B1(new_n719_), .B2(new_n447_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n717_), .B1(new_n720_), .B2(new_n273_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n708_), .B1(new_n721_), .B2(new_n646_), .ZN(new_n722_));
  OAI211_X1 g521(.A(KEYINPUT44), .B(new_n707_), .C1(new_n714_), .C2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT106), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n640_), .A2(new_n645_), .ZN(new_n725_));
  OAI21_X1  g524(.A(KEYINPUT43), .B1(new_n478_), .B2(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n706_), .B1(new_n726_), .B2(new_n713_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n727_), .A2(new_n728_), .A3(KEYINPUT44), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n730_));
  INV_X1    g529(.A(new_n727_), .ZN(new_n731_));
  AOI22_X1  g530(.A1(new_n724_), .A2(new_n729_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n669_), .A2(G29gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n705_), .B1(new_n732_), .B2(new_n733_), .ZN(G1328gat));
  XNOR2_X1  g533(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(G36gat), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n605_), .A2(new_n737_), .A3(new_n474_), .A4(new_n702_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n738_), .B(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n731_), .A2(new_n730_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n723_), .A2(KEYINPUT106), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n728_), .B1(new_n727_), .B2(KEYINPUT44), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n474_), .B(new_n741_), .C1(new_n742_), .C2(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n740_), .B1(new_n744_), .B2(G36gat), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n736_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n737_), .B1(new_n732_), .B2(new_n474_), .ZN(new_n748_));
  OAI211_X1 g547(.A(KEYINPUT107), .B(new_n735_), .C1(new_n748_), .C2(new_n740_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1329gat));
  AOI21_X1  g549(.A(G43gat), .B1(new_n704_), .B2(new_n273_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n273_), .A2(G43gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n732_), .B2(new_n752_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n753_), .B(new_n755_), .ZN(G1330gat));
  INV_X1    g555(.A(G50gat), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n757_), .B1(new_n732_), .B2(new_n390_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n703_), .A2(G50gat), .A3(new_n447_), .ZN(new_n759_));
  OAI21_X1  g558(.A(KEYINPUT110), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n741_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n761_));
  OAI21_X1  g560(.A(G50gat), .B1(new_n761_), .B2(new_n447_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT110), .ZN(new_n763_));
  INV_X1    g562(.A(new_n759_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n762_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n760_), .A2(new_n765_), .ZN(G1331gat));
  INV_X1    g565(.A(G57gat), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n674_), .A2(new_n603_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n768_), .A2(new_n666_), .A3(new_n721_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n767_), .B1(new_n769_), .B2(new_n318_), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n770_), .B(KEYINPUT111), .Z(new_n771_));
  INV_X1    g570(.A(new_n604_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n665_), .A2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n678_), .A2(new_n568_), .A3(new_n773_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n774_), .A2(new_n767_), .A3(new_n318_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n771_), .A2(new_n775_), .ZN(G1332gat));
  OAI21_X1  g575(.A(G64gat), .B1(new_n774_), .B2(new_n715_), .ZN(new_n777_));
  XOR2_X1   g576(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n778_));
  XNOR2_X1  g577(.A(new_n777_), .B(new_n778_), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n715_), .A2(G64gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n779_), .B1(new_n769_), .B2(new_n780_), .ZN(G1333gat));
  OAI21_X1  g580(.A(G71gat), .B1(new_n774_), .B2(new_n477_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT49), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n477_), .A2(G71gat), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n783_), .B1(new_n769_), .B2(new_n784_), .ZN(G1334gat));
  OAI21_X1  g584(.A(G78gat), .B1(new_n774_), .B2(new_n447_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT50), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n447_), .A2(G78gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n769_), .B2(new_n788_), .ZN(G1335gat));
  NOR2_X1   g588(.A1(new_n714_), .A2(new_n722_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT113), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n792_), .B1(new_n714_), .B2(new_n722_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n674_), .A2(new_n700_), .A3(new_n603_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n791_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(G85gat), .B1(new_n795_), .B2(new_n318_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n768_), .A2(new_n721_), .A3(new_n702_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n669_), .A2(new_n481_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n796_), .B1(new_n797_), .B2(new_n798_), .ZN(G1336gat));
  NOR3_X1   g598(.A1(new_n795_), .A2(new_n482_), .A3(new_n715_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n482_), .B1(new_n797_), .B2(new_n715_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT114), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n800_), .A2(new_n802_), .ZN(G1337gat));
  OAI21_X1  g602(.A(G99gat), .B1(new_n795_), .B2(new_n477_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n805_));
  INV_X1    g604(.A(new_n500_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n797_), .A2(new_n806_), .A3(new_n477_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT115), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n804_), .A2(new_n805_), .A3(new_n808_), .ZN(new_n809_));
  OR2_X1    g608(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n809_), .B(new_n810_), .ZN(G1338gat));
  NAND2_X1  g610(.A1(new_n794_), .A2(new_n390_), .ZN(new_n812_));
  OAI21_X1  g611(.A(G106gat), .B1(new_n790_), .B2(new_n812_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n813_), .A2(KEYINPUT52), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n813_), .A2(KEYINPUT52), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n390_), .A2(new_n501_), .ZN(new_n816_));
  OAI22_X1  g615(.A1(new_n814_), .A2(new_n815_), .B1(new_n797_), .B2(new_n816_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g617(.A1(new_n538_), .A2(new_n550_), .A3(new_n553_), .A4(new_n560_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n819_), .A2(new_n603_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n538_), .A2(new_n550_), .A3(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n544_), .A2(new_n539_), .A3(new_n547_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n824_), .B1(KEYINPUT55), .B2(new_n548_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n560_), .B1(new_n822_), .B2(new_n825_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(KEYINPUT118), .A2(KEYINPUT56), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n820_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n827_), .ZN(new_n829_));
  AOI211_X1 g628(.A(new_n560_), .B(new_n829_), .C1(new_n822_), .C2(new_n825_), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT119), .B1(new_n828_), .B2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n823_), .B1(new_n537_), .B2(new_n821_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n544_), .A2(new_n547_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n549_), .B1(new_n833_), .B2(new_n480_), .ZN(new_n834_));
  AOI211_X1 g633(.A(KEYINPUT69), .B(new_n539_), .C1(new_n544_), .C2(new_n547_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n832_), .B1(new_n836_), .B2(new_n821_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n829_), .B1(new_n837_), .B2(new_n560_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT119), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n826_), .A2(new_n827_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n838_), .A2(new_n839_), .A3(new_n840_), .A4(new_n820_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n592_), .A2(new_n583_), .A3(new_n594_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n582_), .A2(new_n585_), .A3(new_n587_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n842_), .B(new_n600_), .C1(new_n843_), .C2(new_n583_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n602_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n563_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n831_), .A2(new_n841_), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n701_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT56), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n852_), .B1(new_n837_), .B2(new_n560_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n826_), .A2(KEYINPUT56), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(KEYINPUT120), .A3(new_n854_), .ZN(new_n855_));
  OR3_X1    g654(.A1(new_n826_), .A2(KEYINPUT120), .A3(KEYINPUT56), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n819_), .A2(new_n846_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n855_), .A2(new_n856_), .A3(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT58), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n855_), .A2(KEYINPUT58), .A3(new_n856_), .A4(new_n857_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n646_), .A3(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n848_), .A2(KEYINPUT57), .A3(new_n701_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n851_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n663_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n773_), .A2(new_n640_), .A3(new_n645_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n868_), .B2(new_n568_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n725_), .A2(new_n674_), .A3(new_n773_), .A4(new_n866_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n865_), .A2(new_n872_), .ZN(new_n873_));
  NOR4_X1   g672(.A1(new_n474_), .A2(new_n390_), .A3(new_n318_), .A4(new_n477_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(G113gat), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n876_), .A2(new_n877_), .A3(new_n603_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n871_), .B1(new_n864_), .B2(new_n665_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n874_), .B(KEYINPUT121), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n879_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(new_n875_), .B2(new_n879_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n883_), .A2(new_n772_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n878_), .B1(new_n884_), .B2(new_n877_), .ZN(G1340gat));
  INV_X1    g684(.A(G120gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n886_), .B1(new_n674_), .B2(KEYINPUT60), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n876_), .B(new_n887_), .C1(KEYINPUT60), .C2(new_n886_), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n883_), .A2(new_n568_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(new_n886_), .ZN(G1341gat));
  INV_X1    g689(.A(G127gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n876_), .A2(new_n891_), .A3(new_n700_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n663_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n883_), .A2(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n892_), .B1(new_n894_), .B2(new_n891_), .ZN(G1342gat));
  INV_X1    g694(.A(G134gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n876_), .A2(new_n896_), .A3(new_n677_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n883_), .A2(new_n646_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n898_), .B2(new_n896_), .ZN(G1343gat));
  NOR2_X1   g698(.A1(new_n447_), .A2(new_n273_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n900_), .A2(new_n715_), .A3(new_n669_), .ZN(new_n901_));
  XOR2_X1   g700(.A(new_n901_), .B(KEYINPUT122), .Z(new_n902_));
  NAND2_X1  g701(.A1(new_n873_), .A2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n603_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(new_n280_), .ZN(G1344gat));
  NOR2_X1   g705(.A1(new_n903_), .A2(new_n674_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(new_n281_), .ZN(G1345gat));
  NOR2_X1   g707(.A1(new_n903_), .A2(new_n665_), .ZN(new_n909_));
  XOR2_X1   g708(.A(KEYINPUT61), .B(G155gat), .Z(new_n910_));
  XNOR2_X1  g709(.A(new_n909_), .B(new_n910_), .ZN(G1346gat));
  INV_X1    g710(.A(G162gat), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n903_), .A2(new_n912_), .A3(new_n725_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n903_), .B2(new_n701_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  OAI211_X1 g715(.A(KEYINPUT123), .B(new_n912_), .C1(new_n903_), .C2(new_n701_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n913_), .B1(new_n916_), .B2(new_n917_), .ZN(G1347gat));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n474_), .A2(new_n716_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n390_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n880_), .A2(new_n904_), .A3(new_n922_), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n923_), .A2(KEYINPUT124), .A3(new_n211_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n848_), .A2(KEYINPUT57), .A3(new_n701_), .ZN(new_n926_));
  AOI21_X1  g725(.A(KEYINPUT57), .B1(new_n848_), .B2(new_n701_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n700_), .B1(new_n928_), .B2(new_n862_), .ZN(new_n929_));
  OAI211_X1 g728(.A(new_n603_), .B(new_n921_), .C1(new_n929_), .C2(new_n871_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n925_), .B1(new_n930_), .B2(G169gat), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n919_), .B1(new_n924_), .B2(new_n931_), .ZN(new_n932_));
  OAI21_X1  g731(.A(KEYINPUT124), .B1(new_n923_), .B2(new_n211_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n930_), .A2(new_n925_), .A3(G169gat), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n933_), .A2(KEYINPUT62), .A3(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n923_), .A2(new_n403_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n932_), .A2(new_n935_), .A3(new_n936_), .ZN(G1348gat));
  OAI21_X1  g736(.A(new_n921_), .B1(new_n929_), .B2(new_n871_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n402_), .B1(new_n938_), .B2(new_n674_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(KEYINPUT125), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n941_));
  OAI211_X1 g740(.A(new_n941_), .B(new_n402_), .C1(new_n938_), .C2(new_n674_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n871_), .B1(new_n864_), .B2(new_n663_), .ZN(new_n943_));
  OR3_X1    g742(.A1(new_n943_), .A2(KEYINPUT126), .A3(new_n390_), .ZN(new_n944_));
  OAI21_X1  g743(.A(KEYINPUT126), .B1(new_n943_), .B2(new_n390_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n674_), .A2(new_n203_), .A3(new_n920_), .ZN(new_n947_));
  AOI22_X1  g746(.A1(new_n940_), .A2(new_n942_), .B1(new_n946_), .B2(new_n947_), .ZN(G1349gat));
  NOR2_X1   g747(.A1(new_n920_), .A2(new_n665_), .ZN(new_n949_));
  AOI21_X1  g748(.A(G183gat), .B1(new_n946_), .B2(new_n949_), .ZN(new_n950_));
  AOI211_X1 g749(.A(new_n663_), .B(new_n938_), .C1(new_n232_), .C2(new_n234_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n950_), .A2(new_n951_), .ZN(G1350gat));
  OAI21_X1  g751(.A(G190gat), .B1(new_n938_), .B2(new_n725_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n677_), .A2(new_n235_), .A3(new_n237_), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n953_), .B1(new_n938_), .B2(new_n954_), .ZN(G1351gat));
  NAND3_X1  g754(.A1(new_n474_), .A2(new_n900_), .A3(new_n318_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n943_), .A2(new_n956_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n957_), .A2(new_n603_), .ZN(new_n958_));
  XNOR2_X1  g757(.A(new_n958_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g758(.A1(new_n957_), .A2(new_n568_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n960_), .B(G204gat), .ZN(G1353gat));
  NOR3_X1   g760(.A1(new_n943_), .A2(new_n663_), .A3(new_n956_), .ZN(new_n962_));
  NOR3_X1   g761(.A1(new_n962_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n963_));
  XOR2_X1   g762(.A(KEYINPUT63), .B(G211gat), .Z(new_n964_));
  AOI21_X1  g763(.A(new_n963_), .B1(new_n962_), .B2(new_n964_), .ZN(G1354gat));
  AOI21_X1  g764(.A(G218gat), .B1(new_n957_), .B2(new_n677_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n646_), .A2(G218gat), .ZN(new_n967_));
  XNOR2_X1  g766(.A(new_n967_), .B(KEYINPUT127), .ZN(new_n968_));
  AOI21_X1  g767(.A(new_n966_), .B1(new_n957_), .B2(new_n968_), .ZN(G1355gat));
endmodule


