//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 0 1 0 1 0 1 1 1 0 1 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n932_, new_n933_, new_n934_, new_n935_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n953_, new_n954_, new_n955_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(KEYINPUT36), .Z(new_n205_));
  XOR2_X1   g004(.A(KEYINPUT68), .B(KEYINPUT34), .Z(new_n206_));
  NAND2_X1  g005(.A1(G232gat), .A2(G233gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT35), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G99gat), .A3(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT7), .ZN(new_n217_));
  INV_X1    g016(.A(G99gat), .ZN(new_n218_));
  INV_X1    g017(.A(G106gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n215_), .A2(new_n216_), .A3(new_n220_), .ZN(new_n221_));
  OR2_X1    g020(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n222_));
  AND2_X1   g021(.A1(G85gat), .A2(G92gat), .ZN(new_n223_));
  AND2_X1   g022(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G85gat), .A2(G92gat), .ZN(new_n225_));
  NOR3_X1   g024(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  AND3_X1   g025(.A1(new_n221_), .A2(new_n222_), .A3(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n222_), .B1(new_n221_), .B2(new_n226_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G29gat), .B(G36gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G43gat), .B(G50gat), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n231_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT10), .B(G99gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n215_), .B1(new_n235_), .B2(G106gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(G92gat), .ZN(new_n238_));
  OAI22_X1  g037(.A1(new_n223_), .A2(new_n225_), .B1(KEYINPUT9), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G85gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(new_n238_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT9), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G85gat), .A2(G92gat), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n239_), .A2(new_n244_), .A3(KEYINPUT64), .ZN(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT64), .B1(new_n239_), .B2(new_n244_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n237_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n229_), .A2(new_n234_), .A3(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n208_), .A2(new_n209_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT15), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n234_), .A2(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n232_), .A2(KEYINPUT15), .A3(new_n233_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n254_), .B1(new_n247_), .B2(new_n229_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n210_), .B1(new_n250_), .B2(new_n255_), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n252_), .A2(new_n253_), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n212_), .A2(new_n214_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n220_), .A2(new_n216_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n226_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n222_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n221_), .A2(new_n222_), .A3(new_n226_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n247_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n257_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n210_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n265_), .A2(new_n248_), .A3(new_n266_), .A4(new_n249_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n256_), .A2(KEYINPUT69), .A3(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT69), .B1(new_n256_), .B2(new_n267_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n205_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT70), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT37), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n256_), .A2(new_n267_), .ZN(new_n273_));
  NOR3_X1   g072(.A1(new_n273_), .A2(KEYINPUT36), .A3(new_n204_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n276_), .B(new_n205_), .C1(new_n268_), .C2(new_n269_), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n271_), .A2(new_n272_), .A3(new_n275_), .A4(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n277_), .A2(new_n275_), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n281_), .A2(KEYINPUT71), .A3(new_n272_), .A4(new_n271_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n205_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n284_), .B1(new_n256_), .B2(new_n267_), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT37), .B1(new_n274_), .B2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n283_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G57gat), .B(G64gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G71gat), .B(G78gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n289_), .A2(new_n290_), .A3(KEYINPUT11), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(KEYINPUT11), .ZN(new_n292_));
  INV_X1    g091(.A(new_n290_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n289_), .A2(KEYINPUT11), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n291_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G15gat), .B(G22gat), .ZN(new_n298_));
  INV_X1    g097(.A(G1gat), .ZN(new_n299_));
  INV_X1    g098(.A(G8gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT14), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G1gat), .B(G8gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G127gat), .B(G155gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G183gat), .B(G211gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n308_), .A2(new_n309_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT17), .ZN(new_n313_));
  NOR3_X1   g112(.A1(new_n311_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT73), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n305_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(G231gat), .ZN(new_n317_));
  INV_X1    g116(.A(G233gat), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n312_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n320_), .A2(KEYINPUT17), .A3(new_n310_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n321_), .A2(KEYINPUT73), .A3(new_n304_), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n316_), .A2(new_n319_), .A3(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n319_), .B1(new_n316_), .B2(new_n322_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n297_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n316_), .A2(new_n322_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n319_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n316_), .A2(new_n319_), .A3(new_n322_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n328_), .A2(new_n296_), .A3(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n313_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n325_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT74), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT74), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n325_), .A2(new_n330_), .A3(new_n334_), .A4(new_n331_), .ZN(new_n335_));
  AND3_X1   g134(.A1(new_n333_), .A2(KEYINPUT75), .A3(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(KEYINPUT75), .B1(new_n333_), .B2(new_n335_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT66), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n296_), .B1(new_n229_), .B2(new_n247_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n339_), .B1(new_n340_), .B2(KEYINPUT12), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n262_), .A2(new_n263_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n239_), .A2(new_n244_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT64), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n239_), .A2(new_n244_), .A3(KEYINPUT64), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n236_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n297_), .B1(new_n342_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT12), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(KEYINPUT66), .A3(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n229_), .A2(new_n247_), .A3(new_n296_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(new_n348_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n297_), .A2(new_n349_), .ZN(new_n353_));
  AOI22_X1  g152(.A1(new_n341_), .A2(new_n350_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G230gat), .A2(G233gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n355_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n352_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G120gat), .B(G148gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT5), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G176gat), .B(G204gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n356_), .A2(new_n358_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n362_), .B(KEYINPUT67), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n366_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n364_), .A2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT13), .ZN(new_n369_));
  NOR3_X1   g168(.A1(new_n288_), .A2(new_n338_), .A3(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT83), .B(G43gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT31), .ZN(new_n372_));
  INV_X1    g171(.A(G169gat), .ZN(new_n373_));
  INV_X1    g172(.A(G176gat), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT22), .B(G169gat), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n377_), .A2(KEYINPUT80), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n373_), .A2(KEYINPUT22), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT80), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n374_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n376_), .B1(new_n378_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT81), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G183gat), .A2(G190gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT23), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT23), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(G183gat), .A3(G190gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT82), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT82), .B1(new_n385_), .B2(new_n386_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  XOR2_X1   g191(.A(KEYINPUT78), .B(G183gat), .Z(new_n393_));
  INV_X1    g192(.A(G190gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n392_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT81), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n397_), .B(new_n376_), .C1(new_n378_), .C2(new_n381_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n383_), .A2(new_n396_), .A3(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT26), .B(G190gat), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT25), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n393_), .A2(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n400_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(G169gat), .A2(G176gat), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT24), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n388_), .A2(new_n407_), .ZN(new_n408_));
  OR2_X1    g207(.A1(new_n408_), .A2(KEYINPUT79), .ZN(new_n409_));
  OR3_X1    g208(.A1(new_n375_), .A2(new_n406_), .A3(new_n405_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(KEYINPUT79), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n404_), .A2(new_n409_), .A3(new_n410_), .A4(new_n411_), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n399_), .A2(KEYINPUT30), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G227gat), .A2(G233gat), .ZN(new_n415_));
  XOR2_X1   g214(.A(new_n415_), .B(G15gat), .Z(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(G71gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(new_n218_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT30), .B1(new_n399_), .B2(new_n412_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n414_), .A2(new_n419_), .A3(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n418_), .B1(new_n413_), .B2(new_n420_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G127gat), .B(G134gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G113gat), .B(G120gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n424_), .A2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n422_), .A2(new_n423_), .A3(new_n427_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n372_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n429_), .A2(new_n372_), .A3(new_n430_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G141gat), .A2(G148gat), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT84), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(KEYINPUT84), .A2(G141gat), .A3(G148gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(G141gat), .ZN(new_n440_));
  INV_X1    g239(.A(G148gat), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n439_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G155gat), .A2(G162gat), .ZN(new_n443_));
  OR2_X1    g242(.A1(new_n443_), .A2(KEYINPUT1), .ZN(new_n444_));
  NOR2_X1   g243(.A1(G155gat), .A2(G162gat), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n444_), .B1(KEYINPUT86), .B2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n446_), .B1(KEYINPUT86), .B2(new_n444_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n443_), .A2(KEYINPUT1), .ZN(new_n448_));
  XOR2_X1   g247(.A(new_n448_), .B(KEYINPUT85), .Z(new_n449_));
  OAI21_X1  g248(.A(new_n442_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT87), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n451_), .B1(new_n439_), .B2(KEYINPUT2), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT2), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n437_), .A2(KEYINPUT87), .A3(new_n453_), .A4(new_n438_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n435_), .A2(new_n453_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT3), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n456_), .B1(G141gat), .B2(G148gat), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n440_), .A2(new_n441_), .A3(KEYINPUT3), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n455_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n452_), .A2(new_n454_), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n443_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n461_), .A2(new_n445_), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n460_), .A2(KEYINPUT88), .A3(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(KEYINPUT88), .B1(new_n460_), .B2(new_n462_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n450_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT29), .ZN(new_n466_));
  NOR2_X1   g265(.A1(KEYINPUT90), .A2(G228gat), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(KEYINPUT90), .A2(G228gat), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n318_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G211gat), .B(G218gat), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  OR2_X1    g272(.A1(G197gat), .A2(G204gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G197gat), .A2(G204gat), .ZN(new_n475_));
  AND2_X1   g274(.A1(KEYINPUT91), .A2(KEYINPUT21), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n474_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n473_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n474_), .A2(new_n475_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT21), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n472_), .A2(new_n474_), .A3(new_n475_), .A4(new_n476_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n478_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT92), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n478_), .A2(new_n482_), .A3(KEYINPUT92), .A4(new_n481_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n466_), .A2(new_n471_), .A3(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G78gat), .B(G106gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n490_), .B(KEYINPUT93), .Z(new_n491_));
  AOI21_X1  g290(.A(new_n483_), .B1(new_n465_), .B2(KEYINPUT29), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n489_), .B(new_n491_), .C1(new_n492_), .C2(new_n471_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT29), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n450_), .B(new_n495_), .C1(new_n463_), .C2(new_n464_), .ZN(new_n496_));
  XOR2_X1   g295(.A(G22gat), .B(G50gat), .Z(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n460_), .A2(new_n462_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT88), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n460_), .A2(KEYINPUT88), .A3(new_n462_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n497_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n503_), .A2(new_n495_), .A3(new_n450_), .A4(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n498_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n498_), .A2(new_n505_), .A3(new_n507_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n494_), .B1(new_n511_), .B2(KEYINPUT94), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n492_), .A2(new_n471_), .ZN(new_n513_));
  AOI211_X1 g312(.A(new_n470_), .B(new_n487_), .C1(new_n465_), .C2(KEYINPUT29), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n511_), .B(new_n490_), .C1(new_n513_), .C2(new_n514_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n498_), .A2(new_n505_), .A3(new_n507_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n507_), .B1(new_n498_), .B2(new_n505_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n491_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n519_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT94), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n518_), .A2(new_n520_), .A3(new_n521_), .A4(new_n493_), .ZN(new_n522_));
  AND3_X1   g321(.A1(new_n512_), .A2(new_n515_), .A3(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n399_), .A2(new_n487_), .A3(new_n412_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G226gat), .A2(G233gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT19), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT20), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n388_), .B1(G183gat), .B2(G190gat), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n375_), .B1(new_n377_), .B2(new_n374_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n392_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT25), .B(G183gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n400_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n410_), .A2(new_n407_), .A3(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n531_), .B1(new_n532_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n483_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n528_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n524_), .A2(new_n527_), .A3(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT96), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT96), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n524_), .A2(new_n541_), .A3(new_n538_), .A4(new_n527_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n487_), .B1(new_n412_), .B2(new_n399_), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n531_), .B(new_n483_), .C1(new_n532_), .C2(new_n535_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT20), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n526_), .B1(new_n543_), .B2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n540_), .A2(new_n542_), .A3(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G8gat), .B(G36gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT18), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G64gat), .B(G92gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n547_), .A2(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n527_), .B1(new_n524_), .B2(new_n538_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n545_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n399_), .A2(new_n412_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n527_), .B(new_n555_), .C1(new_n556_), .C2(new_n487_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n551_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n554_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n552_), .A2(KEYINPUT27), .A3(new_n559_), .ZN(new_n560_));
  NOR3_X1   g359(.A1(new_n543_), .A2(new_n545_), .A3(new_n526_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n551_), .B1(new_n561_), .B2(new_n553_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n559_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT27), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n465_), .A2(new_n428_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n503_), .A2(new_n450_), .A3(new_n427_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G225gat), .A2(G233gat), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n566_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n566_), .A2(new_n567_), .A3(KEYINPUT4), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT4), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n465_), .A2(new_n572_), .A3(new_n428_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n568_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n569_), .B1(new_n571_), .B2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G1gat), .B(G29gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(G85gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(KEYINPUT0), .B(G57gat), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n578_), .B(new_n579_), .Z(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n576_), .A2(new_n581_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n569_), .B(new_n580_), .C1(new_n571_), .C2(new_n575_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n560_), .A2(new_n565_), .A3(new_n582_), .A4(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n434_), .B1(new_n523_), .B2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n570_), .A2(new_n568_), .A3(new_n573_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n566_), .A2(new_n567_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n580_), .B1(new_n587_), .B2(new_n574_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n563_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT95), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT33), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n590_), .B1(new_n583_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n575_), .ZN(new_n593_));
  AOI22_X1  g392(.A1(new_n593_), .A2(new_n570_), .B1(new_n587_), .B2(new_n568_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n594_), .A2(KEYINPUT95), .A3(KEYINPUT33), .A4(new_n580_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n583_), .A2(new_n591_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n589_), .A2(new_n592_), .A3(new_n595_), .A4(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n582_), .A2(new_n583_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n558_), .A2(KEYINPUT32), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n561_), .A2(new_n553_), .A3(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n600_), .B1(new_n547_), .B2(new_n599_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n598_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n512_), .A2(new_n515_), .A3(new_n522_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n597_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n560_), .A2(new_n565_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n512_), .A2(new_n515_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n605_), .B1(new_n606_), .B2(new_n522_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n430_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n427_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n372_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n608_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n583_), .B(new_n582_), .C1(new_n611_), .C2(new_n431_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  AOI22_X1  g412(.A1(new_n585_), .A2(new_n604_), .B1(new_n607_), .B2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n257_), .A2(new_n304_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G229gat), .A2(G233gat), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n617_), .B1(new_n305_), .B2(new_n234_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n305_), .A2(new_n234_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n234_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(new_n304_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  AOI22_X1  g421(.A1(new_n615_), .A2(new_n618_), .B1(new_n622_), .B2(new_n617_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G113gat), .B(G141gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G169gat), .B(G197gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n623_), .B(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n614_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n370_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n633_), .A2(new_n299_), .A3(new_n598_), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n634_), .A2(KEYINPUT97), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(KEYINPUT97), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n635_), .A2(KEYINPUT38), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT98), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(KEYINPUT38), .B1(new_n635_), .B2(new_n636_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n281_), .A2(new_n271_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n614_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n333_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n335_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n647_), .A2(new_n369_), .A3(new_n630_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n643_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n299_), .B1(new_n650_), .B2(new_n598_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n640_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n639_), .A2(new_n652_), .ZN(G1324gat));
  NAND3_X1  g452(.A1(new_n633_), .A2(new_n300_), .A3(new_n605_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT39), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n650_), .A2(new_n605_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n655_), .B1(new_n656_), .B2(G8gat), .ZN(new_n657_));
  AOI211_X1 g456(.A(KEYINPUT39), .B(new_n300_), .C1(new_n650_), .C2(new_n605_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n654_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n659_), .B(new_n660_), .Z(G1325gat));
  INV_X1    g460(.A(new_n434_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n632_), .A2(G15gat), .A3(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT100), .ZN(new_n664_));
  OAI21_X1  g463(.A(G15gat), .B1(new_n649_), .B2(new_n662_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT41), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n665_), .A2(KEYINPUT41), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n664_), .A2(new_n666_), .A3(new_n667_), .ZN(G1326gat));
  OAI21_X1  g467(.A(G22gat), .B1(new_n649_), .B2(new_n603_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n603_), .A2(G22gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(new_n632_), .B2(new_n672_), .ZN(G1327gat));
  INV_X1    g472(.A(new_n338_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n674_), .A2(new_n641_), .A3(new_n369_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(new_n631_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n598_), .ZN(new_n677_));
  OR3_X1    g476(.A1(new_n676_), .A2(G29gat), .A3(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT102), .B1(new_n614_), .B2(new_n287_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n674_), .B1(new_n679_), .B2(KEYINPUT43), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n369_), .A2(new_n630_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n682_));
  OAI211_X1 g481(.A(KEYINPUT102), .B(new_n682_), .C1(new_n614_), .C2(new_n287_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n680_), .A2(KEYINPUT44), .A3(new_n681_), .A4(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n679_), .A2(KEYINPUT43), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n686_), .A2(new_n338_), .A3(new_n681_), .A4(new_n683_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(KEYINPUT103), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n687_), .A2(new_n691_), .A3(new_n688_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n685_), .B1(new_n690_), .B2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n693_), .A2(KEYINPUT104), .A3(new_n598_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(G29gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT104), .B1(new_n693_), .B2(new_n598_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n678_), .B1(new_n695_), .B2(new_n696_), .ZN(G1328gat));
  INV_X1    g496(.A(KEYINPUT105), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(KEYINPUT106), .B2(KEYINPUT46), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n684_), .A2(new_n605_), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n687_), .A2(new_n691_), .A3(new_n688_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n691_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n700_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(G36gat), .ZN(new_n704_));
  INV_X1    g503(.A(new_n676_), .ZN(new_n705_));
  INV_X1    g504(.A(G36gat), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n705_), .A2(new_n706_), .A3(new_n605_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT45), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n699_), .B1(new_n704_), .B2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n684_), .A2(new_n605_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n710_), .B1(new_n690_), .B2(new_n692_), .ZN(new_n711_));
  OAI211_X1 g510(.A(KEYINPUT105), .B(new_n708_), .C1(new_n711_), .C2(new_n706_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT106), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT46), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n709_), .B1(new_n713_), .B2(new_n714_), .ZN(G1329gat));
  NAND3_X1  g514(.A1(new_n693_), .A2(G43gat), .A3(new_n434_), .ZN(new_n716_));
  INV_X1    g515(.A(G43gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n717_), .B1(new_n676_), .B2(new_n662_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT47), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT47), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n716_), .A2(new_n721_), .A3(new_n718_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1330gat));
  AOI21_X1  g522(.A(G50gat), .B1(new_n705_), .B2(new_n523_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n523_), .A2(G50gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n693_), .B2(new_n725_), .ZN(G1331gat));
  INV_X1    g525(.A(G57gat), .ZN(new_n727_));
  INV_X1    g526(.A(new_n369_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n728_), .A2(new_n629_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n643_), .A2(new_n674_), .A3(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT107), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n727_), .B1(new_n731_), .B2(new_n598_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n729_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n733_), .A2(new_n614_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n338_), .B1(new_n286_), .B2(new_n283_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n736_), .A2(G57gat), .A3(new_n677_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n732_), .A2(new_n737_), .ZN(G1332gat));
  INV_X1    g537(.A(new_n736_), .ZN(new_n739_));
  INV_X1    g538(.A(G64gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(new_n740_), .A3(new_n605_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT48), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n731_), .A2(new_n605_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n743_), .B2(G64gat), .ZN(new_n744_));
  AOI211_X1 g543(.A(KEYINPUT48), .B(new_n740_), .C1(new_n731_), .C2(new_n605_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n741_), .B1(new_n744_), .B2(new_n745_), .ZN(G1333gat));
  OR3_X1    g545(.A1(new_n736_), .A2(G71gat), .A3(new_n662_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n731_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G71gat), .B1(new_n748_), .B2(new_n662_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n749_), .A2(KEYINPUT49), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(KEYINPUT49), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n747_), .B1(new_n750_), .B2(new_n751_), .ZN(G1334gat));
  INV_X1    g551(.A(G78gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n739_), .A2(new_n753_), .A3(new_n523_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n731_), .A2(new_n523_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(G78gat), .ZN(new_n757_));
  AOI211_X1 g556(.A(KEYINPUT50), .B(new_n753_), .C1(new_n731_), .C2(new_n523_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(G1335gat));
  NOR2_X1   g558(.A1(new_n674_), .A2(new_n641_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n734_), .A2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n240_), .B1(new_n761_), .B2(new_n677_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT108), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n680_), .A2(new_n683_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n764_), .A2(new_n733_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n677_), .A2(new_n240_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n763_), .B1(new_n765_), .B2(new_n766_), .ZN(G1336gat));
  INV_X1    g566(.A(new_n761_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n768_), .A2(new_n238_), .A3(new_n605_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n605_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n764_), .A2(new_n770_), .A3(new_n733_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n769_), .B1(new_n771_), .B2(new_n238_), .ZN(new_n772_));
  XOR2_X1   g571(.A(new_n772_), .B(KEYINPUT109), .Z(G1337gat));
  NOR3_X1   g572(.A1(new_n761_), .A2(new_n662_), .A3(new_n235_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n765_), .A2(new_n434_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(G99gat), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g576(.A1(new_n768_), .A2(new_n219_), .A3(new_n523_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n765_), .A2(new_n523_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n780_), .B2(G106gat), .ZN(new_n781_));
  AOI211_X1 g580(.A(KEYINPUT52), .B(new_n219_), .C1(new_n765_), .C2(new_n523_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT53), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n785_), .B(new_n778_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1339gat));
  NAND4_X1  g586(.A1(new_n287_), .A2(new_n674_), .A3(new_n630_), .A4(new_n728_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT54), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT54), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n735_), .A2(new_n790_), .A3(new_n630_), .A4(new_n728_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n623_), .A2(new_n628_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n628_), .B1(new_n622_), .B2(new_n616_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n615_), .A2(new_n619_), .A3(new_n617_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n793_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(new_n364_), .B2(new_n367_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n363_), .A2(new_n629_), .ZN(new_n800_));
  AND4_X1   g599(.A1(new_n247_), .A2(new_n262_), .A3(new_n296_), .A4(new_n263_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n353_), .B1(new_n340_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n803_), .B1(new_n357_), .B2(KEYINPUT110), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n803_), .B2(new_n357_), .ZN(new_n805_));
  AOI211_X1 g604(.A(new_n339_), .B(KEYINPUT12), .C1(new_n264_), .C2(new_n297_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT66), .B1(new_n348_), .B2(new_n349_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n802_), .B(new_n805_), .C1(new_n806_), .C2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n804_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n808_), .B(new_n365_), .C1(new_n354_), .C2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT56), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT111), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n810_), .A2(new_n811_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n810_), .A2(KEYINPUT111), .A3(new_n811_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n800_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n799_), .B1(new_n817_), .B2(KEYINPUT112), .ZN(new_n818_));
  INV_X1    g617(.A(new_n800_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n802_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n366_), .B1(new_n820_), .B2(new_n804_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n821_), .A2(KEYINPUT56), .A3(new_n808_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT56), .B1(new_n821_), .B2(new_n808_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n823_), .B2(KEYINPUT111), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n819_), .B(KEYINPUT112), .C1(new_n824_), .C2(new_n815_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n641_), .B1(new_n818_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT57), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT112), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n815_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n800_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(new_n825_), .A3(new_n799_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(new_n833_), .A3(new_n641_), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT113), .B1(new_n364_), .B2(new_n797_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT113), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n363_), .A2(new_n836_), .A3(new_n798_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n835_), .B(new_n837_), .C1(new_n813_), .C2(new_n823_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(KEYINPUT58), .ZN(new_n839_));
  AOI22_X1  g638(.A1(new_n828_), .A2(new_n834_), .B1(new_n288_), .B2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n792_), .B1(new_n840_), .B2(new_n646_), .ZN(new_n841_));
  NOR4_X1   g640(.A1(new_n662_), .A2(new_n523_), .A3(new_n605_), .A4(new_n677_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(G113gat), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(new_n845_), .A3(new_n629_), .ZN(new_n846_));
  OAI21_X1  g645(.A(KEYINPUT115), .B1(new_n840_), .B2(new_n674_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n839_), .A2(new_n288_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n799_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n819_), .B1(new_n824_), .B2(new_n815_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(new_n829_), .ZN(new_n851_));
  AOI211_X1 g650(.A(KEYINPUT57), .B(new_n642_), .C1(new_n851_), .C2(new_n825_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n833_), .B1(new_n832_), .B2(new_n641_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n848_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n854_), .A2(new_n855_), .A3(new_n338_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n847_), .A2(new_n856_), .A3(new_n792_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT114), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n842_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n842_), .A2(new_n858_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n859_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n857_), .A2(KEYINPUT116), .A3(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT116), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n865_), .B1(new_n843_), .B2(KEYINPUT59), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n789_), .A2(new_n791_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n854_), .A2(new_n338_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n868_), .B2(KEYINPUT115), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n862_), .B1(new_n869_), .B2(new_n856_), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n629_), .B(new_n864_), .C1(new_n866_), .C2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n846_), .B1(new_n872_), .B2(new_n845_), .ZN(G1340gat));
  INV_X1    g672(.A(G120gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n874_), .B1(new_n728_), .B2(KEYINPUT60), .ZN(new_n875_));
  OR2_X1    g674(.A1(new_n874_), .A2(KEYINPUT60), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n841_), .A2(new_n842_), .A3(new_n875_), .A4(new_n876_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(KEYINPUT117), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n369_), .B(new_n864_), .C1(new_n866_), .C2(new_n870_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n878_), .B1(new_n880_), .B2(new_n874_), .ZN(G1341gat));
  INV_X1    g680(.A(G127gat), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n844_), .A2(new_n882_), .A3(new_n674_), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n646_), .B(new_n864_), .C1(new_n866_), .C2(new_n870_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n883_), .B1(new_n885_), .B2(new_n882_), .ZN(G1342gat));
  INV_X1    g685(.A(G134gat), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n844_), .A2(new_n887_), .A3(new_n642_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n288_), .B(new_n864_), .C1(new_n866_), .C2(new_n870_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n888_), .B1(new_n890_), .B2(new_n887_), .ZN(G1343gat));
  NOR4_X1   g690(.A1(new_n603_), .A2(new_n434_), .A3(new_n677_), .A4(new_n605_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n841_), .A2(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n893_), .A2(new_n630_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(new_n440_), .ZN(G1344gat));
  NOR2_X1   g694(.A1(new_n893_), .A2(new_n728_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(new_n441_), .ZN(G1345gat));
  NOR2_X1   g696(.A1(new_n893_), .A2(new_n338_), .ZN(new_n898_));
  XOR2_X1   g697(.A(KEYINPUT61), .B(G155gat), .Z(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(G1346gat));
  OAI21_X1  g699(.A(G162gat), .B1(new_n893_), .B2(new_n287_), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n641_), .A2(G162gat), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n893_), .B2(new_n902_), .ZN(G1347gat));
  NOR2_X1   g702(.A1(new_n612_), .A2(new_n770_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n629_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(KEYINPUT118), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n906_), .A2(new_n523_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n373_), .B1(new_n857_), .B2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n904_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(new_n523_), .ZN(new_n912_));
  AND2_X1   g711(.A1(new_n857_), .A2(new_n912_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n913_), .A2(new_n629_), .A3(new_n377_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n910_), .A2(new_n914_), .ZN(G1348gat));
  NAND2_X1  g714(.A1(new_n841_), .A2(new_n603_), .ZN(new_n916_));
  NOR4_X1   g715(.A1(new_n916_), .A2(new_n374_), .A3(new_n728_), .A4(new_n911_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n913_), .A2(new_n369_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(new_n918_), .B2(new_n374_), .ZN(G1349gat));
  NOR2_X1   g718(.A1(new_n647_), .A2(new_n533_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n857_), .A2(new_n912_), .A3(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(KEYINPUT119), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT119), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n857_), .A2(new_n923_), .A3(new_n912_), .A4(new_n920_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n674_), .A2(new_n904_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n393_), .B1(new_n916_), .B2(new_n925_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n922_), .A2(new_n924_), .A3(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(KEYINPUT120), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT120), .ZN(new_n929_));
  NAND4_X1  g728(.A1(new_n922_), .A2(new_n929_), .A3(new_n924_), .A4(new_n926_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n928_), .A2(new_n930_), .ZN(G1350gat));
  NAND2_X1  g730(.A1(new_n642_), .A2(new_n400_), .ZN(new_n932_));
  XOR2_X1   g731(.A(new_n932_), .B(KEYINPUT121), .Z(new_n933_));
  NAND2_X1  g732(.A1(new_n913_), .A2(new_n933_), .ZN(new_n934_));
  AND2_X1   g733(.A1(new_n913_), .A2(new_n288_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n935_), .B2(new_n394_), .ZN(G1351gat));
  INV_X1    g735(.A(KEYINPUT123), .ZN(new_n937_));
  AOI22_X1  g736(.A1(new_n854_), .A2(new_n647_), .B1(new_n789_), .B2(new_n791_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n662_), .A2(new_n523_), .A3(new_n677_), .ZN(new_n939_));
  INV_X1    g738(.A(new_n939_), .ZN(new_n940_));
  OR2_X1    g739(.A1(new_n940_), .A2(KEYINPUT122), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(KEYINPUT122), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n941_), .A2(new_n605_), .A3(new_n942_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n937_), .B1(new_n938_), .B2(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(new_n943_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n828_), .A2(new_n834_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n646_), .B1(new_n946_), .B2(new_n848_), .ZN(new_n947_));
  OAI211_X1 g746(.A(new_n945_), .B(KEYINPUT123), .C1(new_n947_), .C2(new_n867_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n944_), .A2(new_n948_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n949_), .A2(new_n629_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(KEYINPUT124), .B(G197gat), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n950_), .B(new_n951_), .ZN(G1352gat));
  NAND2_X1  g751(.A1(new_n949_), .A2(new_n369_), .ZN(new_n953_));
  INV_X1    g752(.A(G204gat), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n954_), .A2(KEYINPUT125), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n953_), .B(new_n955_), .ZN(G1353gat));
  NAND2_X1  g755(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n957_));
  AOI21_X1  g756(.A(KEYINPUT126), .B1(new_n646_), .B2(new_n957_), .ZN(new_n958_));
  AND3_X1   g757(.A1(new_n646_), .A2(KEYINPUT126), .A3(new_n957_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n949_), .B1(new_n958_), .B2(new_n959_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n961_));
  XOR2_X1   g760(.A(new_n960_), .B(new_n961_), .Z(G1354gat));
  INV_X1    g761(.A(G218gat), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n963_), .B1(new_n949_), .B2(new_n288_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n641_), .A2(G218gat), .ZN(new_n965_));
  INV_X1    g764(.A(new_n965_), .ZN(new_n966_));
  AOI21_X1  g765(.A(new_n966_), .B1(new_n944_), .B2(new_n948_), .ZN(new_n967_));
  OAI21_X1  g766(.A(KEYINPUT127), .B1(new_n964_), .B2(new_n967_), .ZN(new_n968_));
  INV_X1    g767(.A(new_n967_), .ZN(new_n969_));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n970_));
  AOI21_X1  g769(.A(new_n287_), .B1(new_n944_), .B2(new_n948_), .ZN(new_n971_));
  OAI211_X1 g770(.A(new_n969_), .B(new_n970_), .C1(new_n963_), .C2(new_n971_), .ZN(new_n972_));
  AND2_X1   g771(.A1(new_n968_), .A2(new_n972_), .ZN(G1355gat));
endmodule


