//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 0 0 1 0 0 0' ..
//Module:
 module locked_locked_c1355( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat,
    G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat,
    G85gat, G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat,
    G141gat, G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat,
    G197gat, G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat,
    G229gat, G230gat, G231gat, G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  , KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64);
input KEYINPUT64;
input KEYINPUT65;
input KEYINPUT66;
input KEYINPUT67;
input KEYINPUT68;
input KEYINPUT69;
input KEYINPUT70;
input KEYINPUT71;
input KEYINPUT72;
input KEYINPUT73;
input KEYINPUT74;
input KEYINPUT75;
input KEYINPUT76;
input KEYINPUT77;
input KEYINPUT78;
input KEYINPUT79;
input KEYINPUT80;
input KEYINPUT81;
input KEYINPUT82;
input KEYINPUT83;
input KEYINPUT84;
input KEYINPUT85;
input KEYINPUT86;
input KEYINPUT87;
input KEYINPUT88;
input KEYINPUT89;
input KEYINPUT90;
input KEYINPUT91;
input KEYINPUT92;
input KEYINPUT93;
input KEYINPUT94;
input KEYINPUT95;
input KEYINPUT96;
input KEYINPUT97;
input KEYINPUT98;
input KEYINPUT99;
input KEYINPUT100;
input KEYINPUT101;
input KEYINPUT102;
input KEYINPUT103;
input KEYINPUT104;
input KEYINPUT105;
input KEYINPUT106;
input KEYINPUT107;
input KEYINPUT108;
input KEYINPUT109;
input KEYINPUT110;
input KEYINPUT111;
input KEYINPUT112;
input KEYINPUT113;
input KEYINPUT114;
input KEYINPUT115;
input KEYINPUT116;
input KEYINPUT117;
input KEYINPUT118;
input KEYINPUT119;
input KEYINPUT120;
input KEYINPUT121;
input KEYINPUT122;
input KEYINPUT123;
input KEYINPUT124;
input KEYINPUT125;
input KEYINPUT126;
input KEYINPUT127;
//Header:
   input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat,
    G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat,
    G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, G113gat, G120gat,
    G127gat, G134gat, G141gat, G148gat, G155gat, G162gat, G169gat, G176gat,
    G183gat, G190gat, G197gat, G204gat, G211gat, G218gat, G225gat, G226gat,
    G227gat, G228gat, G229gat, G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n477_, new_n478_, new_n480_, new_n481_,
    new_n482_, new_n484_, new_n485_, new_n486_, new_n487_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n516_, new_n517_, new_n518_, new_n519_, new_n521_, new_n522_,
    new_n523_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n534_, new_n535_, new_n536_,
    new_n538_, new_n539_, new_n540_, new_n542_, new_n543_, new_n544_,
    new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n552_, new_n554_, new_n555_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n626_, new_n627_, new_n628_, new_n630_,
    new_n631_, new_n632_, new_n634_, new_n635_, new_n636_, new_n638_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n659_, new_n660_, new_n662_,
    new_n663_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_;
wire RLL_wire_A_64;
wire RLL_wire_A_65;
wire RLL_wire_A_66;
wire RLL_wire_A_67;
wire RLL_wire_A_68;
wire RLL_wire_A_69;
wire RLL_wire_A_70;
wire RLL_wire_A_71;
wire RLL_wire_A_72;
wire RLL_wire_A_73;
wire RLL_wire_A_74;
wire RLL_wire_A_75;
wire RLL_wire_A_76;
wire RLL_wire_A_77;
wire RLL_wire_A_78;
wire RLL_wire_A_79;
wire RLL_wire_A_80;
wire RLL_wire_A_81;
wire RLL_wire_A_82;
wire RLL_wire_A_83;
wire RLL_wire_A_84;
wire RLL_wire_A_85;
wire RLL_wire_A_86;
wire RLL_wire_A_87;
wire RLL_wire_A_88;
wire RLL_wire_A_89;
wire RLL_wire_A_90;
wire RLL_wire_A_91;
wire RLL_wire_A_92;
wire RLL_wire_A_93;
wire RLL_wire_A_94;
wire RLL_wire_A_95;
wire RLL_wire_A_96;
wire RLL_wire_A_97;
wire RLL_wire_A_98;
wire RLL_wire_A_99;
wire RLL_wire_A_100;
wire RLL_wire_A_101;
wire RLL_wire_A_102;
wire RLL_wire_A_103;
wire RLL_wire_A_104;
wire RLL_wire_A_105;
wire RLL_wire_A_106;
wire RLL_wire_A_107;
wire RLL_wire_A_108;
wire RLL_wire_A_109;
wire RLL_wire_A_110;
wire RLL_wire_A_111;
wire RLL_wire_A_112;
wire RLL_wire_A_113;
wire RLL_wire_A_114;
wire RLL_wire_A_115;
wire RLL_wire_A_116;
wire RLL_wire_A_117;
wire RLL_wire_A_118;
wire RLL_wire_A_119;
wire RLL_wire_A_120;
wire RLL_wire_A_121;
wire RLL_wire_A_122;
wire RLL_wire_A_123;
wire RLL_wire_A_124;
wire RLL_wire_A_125;
wire RLL_wire_A_126;
wire RLL_wire_A_127;

//Body:
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n138_));
  INV_X1    g001(.A(new_n138_), .ZN(new_n139_));
  XOR2_X1   g002(.A(KEYINPUT10), .B(G99gat), .Z(new_n140_));
  INV_X1    g003(.A(G106gat), .ZN(new_n141_));
  NAND2_X1  g004(.A1(new_n140_), .A2(new_n141_), .ZN(new_n142_));
  INV_X1    g005(.A(KEYINPUT9), .ZN(new_n143_));
  INV_X1    g006(.A(G85gat), .ZN(new_n144_));
  INV_X1    g007(.A(G92gat), .ZN(RLL_wire_A_64));
  XNOR2_X1 RLL_XNOR_64 (.A(RLL_wire_A_64), .B(KEYINPUT64), .ZN(new_n145_) );
  OAI21_X1  g008(.A(new_n143_), .B1(new_n144_), .B2(new_n145_), .ZN(new_n146_));
  NAND3_X1  g009(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n147_));
  OAI211_X1 g010(.A(new_n146_), .B(new_n147_), .C1(G85gat), .C2(G92gat), .ZN(new_n148_));
  NAND2_X1  g011(.A1(G99gat), .A2(G106gat), .ZN(new_n149_));
  XNOR2_X1  g012(.A(new_n149_), .B(KEYINPUT6), .ZN(new_n150_));
  AND3_X1   g013(.A1(new_n142_), .A2(new_n148_), .A3(new_n150_), .ZN(new_n151_));
  OAI21_X1  g014(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(RLL_wire_A_65));
  XNOR2_X1 RLL_XNOR_65 (.A(RLL_wire_A_65), .B(KEYINPUT65), .ZN(new_n152_) );
  NOR2_X1   g015(.A1(G99gat), .A2(G106gat), .ZN(new_n153_));
  INV_X1    g016(.A(KEYINPUT7), .ZN(new_n154_));
  NAND2_X1  g017(.A1(new_n153_), .A2(new_n154_), .ZN(new_n155_));
  NAND3_X1  g018(.A1(new_n150_), .A2(new_n152_), .A3(new_n155_), .ZN(new_n156_));
  INV_X1    g019(.A(KEYINPUT8), .ZN(new_n157_));
  XOR2_X1   g020(.A(G85gat), .B(G92gat), .Z(new_n158_));
  NAND3_X1  g021(.A1(new_n156_), .A2(new_n157_), .A3(new_n158_), .ZN(RLL_wire_A_66));
  XNOR2_X1 RLL_XNOR_66 (.A(RLL_wire_A_66), .B(KEYINPUT66), .ZN(new_n159_) );
  INV_X1    g022(.A(KEYINPUT6), .ZN(new_n160_));
  XNOR2_X1  g023(.A(new_n149_), .B(new_n160_), .ZN(new_n161_));
  NAND2_X1  g024(.A1(new_n155_), .A2(new_n152_), .ZN(RLL_wire_A_67));
  XOR2_X1 RLL_XOR_67 (.A(RLL_wire_A_67), .B(KEYINPUT67), .Z(new_n162_) );
  OAI21_X1  g025(.A(new_n158_), .B1(new_n161_), .B2(new_n162_), .ZN(new_n163_));
  NAND2_X1  g026(.A1(new_n163_), .A2(KEYINPUT8), .ZN(new_n164_));
  AOI21_X1  g027(.A(new_n151_), .B1(new_n159_), .B2(new_n164_), .ZN(RLL_wire_A_68));
  XNOR2_X1 RLL_XNOR_68 (.A(RLL_wire_A_68), .B(KEYINPUT68), .ZN(new_n165_) );
  XOR2_X1   g028(.A(G71gat), .B(G78gat), .Z(new_n166_));
  XNOR2_X1  g029(.A(G57gat), .B(G64gat), .ZN(new_n167_));
  OAI21_X1  g030(.A(new_n166_), .B1(KEYINPUT11), .B2(new_n167_), .ZN(RLL_wire_A_69));
  XNOR2_X1 RLL_XNOR_69 (.A(RLL_wire_A_69), .B(KEYINPUT69), .ZN(new_n168_) );
  NAND2_X1  g031(.A1(new_n167_), .A2(KEYINPUT11), .ZN(new_n169_));
  XOR2_X1   g032(.A(new_n168_), .B(new_n169_), .Z(new_n170_));
  NAND2_X1  g033(.A1(new_n165_), .A2(new_n170_), .ZN(new_n171_));
  INV_X1    g034(.A(new_n171_), .ZN(new_n172_));
  NOR2_X1   g035(.A1(new_n165_), .A2(new_n170_), .ZN(new_n173_));
  OAI21_X1  g036(.A(new_n139_), .B1(new_n172_), .B2(new_n173_), .ZN(new_n174_));
  NAND2_X1  g037(.A1(new_n159_), .A2(new_n164_), .ZN(RLL_wire_A_70));
  XNOR2_X1 RLL_XNOR_70 (.A(RLL_wire_A_70), .B(KEYINPUT70), .ZN(new_n175_) );
  INV_X1    g038(.A(new_n151_), .ZN(new_n176_));
  NAND2_X1  g039(.A1(new_n175_), .A2(new_n176_), .ZN(new_n177_));
  XNOR2_X1  g040(.A(new_n168_), .B(new_n169_), .ZN(new_n178_));
  NAND3_X1  g041(.A1(new_n177_), .A2(KEYINPUT12), .A3(new_n178_), .ZN(new_n179_));
  INV_X1    g042(.A(KEYINPUT12), .ZN(new_n180_));
  OAI21_X1  g043(.A(new_n180_), .B1(new_n165_), .B2(new_n170_), .ZN(RLL_wire_A_71));
  XOR2_X1 RLL_XOR_71 (.A(RLL_wire_A_71), .B(KEYINPUT71), .Z(new_n181_) );
  AOI21_X1  g044(.A(new_n139_), .B1(new_n165_), .B2(new_n170_), .ZN(new_n182_));
  NAND3_X1  g045(.A1(new_n179_), .A2(new_n181_), .A3(new_n182_), .ZN(new_n183_));
  NAND2_X1  g046(.A1(new_n174_), .A2(new_n183_), .ZN(new_n184_));
  XOR2_X1   g047(.A(G120gat), .B(G148gat), .Z(new_n185_));
  XNOR2_X1  g048(.A(new_n185_), .B(KEYINPUT5), .ZN(new_n186_));
  XNOR2_X1  g049(.A(G176gat), .B(G204gat), .ZN(new_n187_));
  XOR2_X1   g050(.A(new_n186_), .B(new_n187_), .Z(new_n188_));
  INV_X1    g051(.A(new_n188_), .ZN(RLL_wire_A_72));
  XNOR2_X1 RLL_XNOR_72 (.A(RLL_wire_A_72), .B(KEYINPUT72), .ZN(new_n189_) );
  NAND2_X1  g052(.A1(new_n184_), .A2(new_n189_), .ZN(new_n190_));
  NAND3_X1  g053(.A1(new_n174_), .A2(new_n183_), .A3(new_n188_), .ZN(new_n191_));
  NAND2_X1  g054(.A1(new_n190_), .A2(new_n191_), .ZN(new_n192_));
  OR2_X1    g055(.A1(new_n192_), .A2(KEYINPUT13), .ZN(new_n193_));
  NAND2_X1  g056(.A1(new_n192_), .A2(KEYINPUT13), .ZN(new_n194_));
  NAND2_X1  g057(.A1(new_n193_), .A2(new_n194_), .ZN(new_n195_));
  INV_X1    g058(.A(new_n195_), .ZN(new_n196_));
  NAND2_X1  g059(.A1(G232gat), .A2(G233gat), .ZN(new_n197_));
  XOR2_X1   g060(.A(new_n197_), .B(KEYINPUT34), .Z(RLL_wire_A_73));
  XNOR2_X1 RLL_XNOR_73 (.A(RLL_wire_A_73), .B(KEYINPUT73), .ZN(new_n198_) );
  INV_X1    g061(.A(KEYINPUT35), .ZN(new_n199_));
  NOR2_X1   g062(.A1(new_n198_), .A2(new_n199_), .ZN(new_n200_));
  XNOR2_X1  g063(.A(G29gat), .B(G36gat), .ZN(new_n201_));
  XNOR2_X1  g064(.A(G43gat), .B(G50gat), .ZN(new_n202_));
  XNOR2_X1  g065(.A(new_n201_), .B(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g066(.A(new_n203_), .B(KEYINPUT15), .ZN(new_n204_));
  NAND2_X1  g067(.A1(new_n177_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g068(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g069(.A1(new_n165_), .A2(new_n203_), .ZN(new_n207_));
  NAND2_X1  g070(.A1(new_n198_), .A2(new_n199_), .ZN(new_n208_));
  NAND2_X1  g071(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  OAI21_X1  g072(.A(new_n200_), .B1(new_n206_), .B2(new_n209_), .ZN(new_n210_));
  XOR2_X1   g073(.A(G190gat), .B(G218gat), .Z(new_n211_));
  XNOR2_X1  g074(.A(G134gat), .B(G162gat), .ZN(new_n212_));
  XNOR2_X1  g075(.A(new_n211_), .B(new_n212_), .ZN(RLL_wire_A_74));
  XNOR2_X1 RLL_XNOR_74 (.A(RLL_wire_A_74), .B(KEYINPUT74), .ZN(new_n213_) );
  INV_X1    g076(.A(KEYINPUT36), .ZN(new_n214_));
  NAND2_X1  g077(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g078(.A(new_n215_), .ZN(new_n216_));
  INV_X1    g079(.A(new_n200_), .ZN(new_n217_));
  NAND4_X1  g080(.A1(new_n205_), .A2(new_n207_), .A3(new_n217_), .A4(new_n208_), .ZN(new_n218_));
  NAND3_X1  g081(.A1(new_n210_), .A2(new_n216_), .A3(new_n218_), .ZN(RLL_wire_A_75));
  XOR2_X1 RLL_XOR_75 (.A(RLL_wire_A_75), .B(KEYINPUT75), .Z(new_n219_) );
  INV_X1    g082(.A(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g083(.A(new_n213_), .B(KEYINPUT36), .ZN(new_n221_));
  INV_X1    g084(.A(new_n221_), .ZN(new_n222_));
  AOI21_X1  g085(.A(new_n222_), .B1(new_n210_), .B2(new_n218_), .ZN(new_n223_));
  OAI21_X1  g086(.A(KEYINPUT37), .B1(new_n220_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g087(.A1(new_n210_), .A2(new_n218_), .ZN(new_n225_));
  NAND2_X1  g088(.A1(new_n225_), .A2(new_n221_), .ZN(new_n226_));
  INV_X1    g089(.A(KEYINPUT37), .ZN(new_n227_));
  NAND3_X1  g090(.A1(new_n226_), .A2(new_n227_), .A3(new_n219_), .ZN(new_n228_));
  NAND2_X1  g091(.A1(new_n224_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g092(.A(G15gat), .B(G22gat), .ZN(new_n230_));
  INV_X1    g093(.A(G1gat), .ZN(new_n231_));
  INV_X1    g094(.A(G8gat), .ZN(new_n232_));
  OAI21_X1  g095(.A(KEYINPUT14), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g096(.A1(new_n230_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g097(.A(G1gat), .B(G8gat), .ZN(new_n235_));
  XNOR2_X1  g098(.A(new_n234_), .B(new_n235_), .ZN(RLL_wire_A_76));
  XOR2_X1 RLL_XOR_76 (.A(RLL_wire_A_76), .B(KEYINPUT76), .Z(new_n236_) );
  NAND2_X1  g099(.A1(G231gat), .A2(G233gat), .ZN(new_n237_));
  XNOR2_X1  g100(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g101(.A(new_n238_), .B(new_n178_), .ZN(new_n239_));
  XOR2_X1   g102(.A(G127gat), .B(G155gat), .Z(new_n240_));
  XNOR2_X1  g103(.A(new_n240_), .B(KEYINPUT16), .ZN(new_n241_));
  XNOR2_X1  g104(.A(G183gat), .B(G211gat), .ZN(new_n242_));
  XNOR2_X1  g105(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  INV_X1    g106(.A(KEYINPUT17), .ZN(new_n244_));
  NOR2_X1   g107(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g108(.A1(new_n239_), .A2(new_n245_), .ZN(RLL_wire_A_77));
  XOR2_X1 RLL_XOR_77 (.A(RLL_wire_A_77), .B(KEYINPUT77), .Z(new_n246_) );
  XNOR2_X1  g109(.A(new_n238_), .B(new_n170_), .ZN(new_n247_));
  XNOR2_X1  g110(.A(new_n243_), .B(KEYINPUT17), .ZN(new_n248_));
  NAND2_X1  g111(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g112(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g113(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g114(.A1(new_n229_), .A2(new_n251_), .ZN(new_n252_));
  NOR2_X1   g115(.A1(new_n196_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g116(.A(new_n203_), .ZN(RLL_wire_A_78));
  XNOR2_X1 RLL_XNOR_78 (.A(RLL_wire_A_78), .B(KEYINPUT78), .ZN(new_n254_) );
  OR2_X1    g117(.A1(new_n236_), .A2(new_n254_), .ZN(RLL_wire_A_79));
  XNOR2_X1 RLL_XNOR_79 (.A(RLL_wire_A_79), .B(KEYINPUT79), .ZN(new_n255_) );
  NAND2_X1  g118(.A1(new_n236_), .A2(new_n254_), .ZN(new_n256_));
  NAND2_X1  g119(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g120(.A1(new_n257_), .A2(G229gat), .A3(G233gat), .ZN(new_n258_));
  NAND2_X1  g121(.A1(new_n204_), .A2(new_n236_), .ZN(new_n259_));
  NAND2_X1  g122(.A1(G229gat), .A2(G233gat), .ZN(new_n260_));
  NAND3_X1  g123(.A1(new_n259_), .A2(new_n260_), .A3(new_n255_), .ZN(new_n261_));
  NAND2_X1  g124(.A1(new_n258_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g125(.A(G113gat), .B(G141gat), .ZN(new_n263_));
  XNOR2_X1  g126(.A(G169gat), .B(G197gat), .ZN(new_n264_));
  XOR2_X1   g127(.A(new_n263_), .B(new_n264_), .Z(new_n265_));
  INV_X1    g128(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g129(.A1(new_n262_), .A2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g130(.A1(new_n258_), .A2(new_n261_), .A3(new_n265_), .ZN(new_n268_));
  NAND2_X1  g131(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g132(.A(new_n269_), .ZN(RLL_wire_A_80));
  XOR2_X1 RLL_XOR_80 (.A(RLL_wire_A_80), .B(KEYINPUT80), .Z(new_n270_) );
  INV_X1    g133(.A(G183gat), .ZN(new_n271_));
  NAND2_X1  g134(.A1(new_n271_), .A2(KEYINPUT25), .ZN(new_n272_));
  INV_X1    g135(.A(KEYINPUT25), .ZN(new_n273_));
  NAND2_X1  g136(.A1(new_n273_), .A2(G183gat), .ZN(new_n274_));
  INV_X1    g137(.A(G190gat), .ZN(new_n275_));
  NAND2_X1  g138(.A1(new_n275_), .A2(KEYINPUT26), .ZN(new_n276_));
  INV_X1    g139(.A(KEYINPUT26), .ZN(new_n277_));
  NAND2_X1  g140(.A1(new_n277_), .A2(G190gat), .ZN(new_n278_));
  NAND4_X1  g141(.A1(new_n272_), .A2(new_n274_), .A3(new_n276_), .A4(new_n278_), .ZN(new_n279_));
  NOR2_X1   g142(.A1(G169gat), .A2(G176gat), .ZN(new_n280_));
  INV_X1    g143(.A(new_n280_), .ZN(RLL_wire_A_81));
  XNOR2_X1 RLL_XNOR_81 (.A(RLL_wire_A_81), .B(KEYINPUT81), .ZN(new_n281_) );
  NAND2_X1  g144(.A1(G169gat), .A2(G176gat), .ZN(new_n282_));
  NAND3_X1  g145(.A1(new_n281_), .A2(KEYINPUT24), .A3(new_n282_), .ZN(new_n283_));
  NAND2_X1  g146(.A1(new_n279_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g147(.A(KEYINPUT23), .ZN(new_n285_));
  AOI21_X1  g148(.A(new_n285_), .B1(G183gat), .B2(G190gat), .ZN(new_n286_));
  NAND2_X1  g149(.A1(G183gat), .A2(G190gat), .ZN(new_n287_));
  NOR2_X1   g150(.A1(new_n287_), .A2(KEYINPUT23), .ZN(new_n288_));
  OAI22_X1  g151(.A1(new_n286_), .A2(new_n288_), .B1(new_n281_), .B2(KEYINPUT24), .ZN(new_n289_));
  INV_X1    g152(.A(G169gat), .ZN(new_n290_));
  NAND2_X1  g153(.A1(new_n290_), .A2(KEYINPUT22), .ZN(new_n291_));
  INV_X1    g154(.A(KEYINPUT22), .ZN(new_n292_));
  NAND2_X1  g155(.A1(new_n292_), .A2(G169gat), .ZN(new_n293_));
  INV_X1    g156(.A(G176gat), .ZN(new_n294_));
  NAND3_X1  g157(.A1(new_n291_), .A2(new_n293_), .A3(new_n294_), .ZN(RLL_wire_A_82));
  XOR2_X1 RLL_XOR_82 (.A(RLL_wire_A_82), .B(KEYINPUT82), .Z(new_n295_) );
  NAND2_X1  g158(.A1(new_n295_), .A2(new_n282_), .ZN(new_n296_));
  NAND2_X1  g159(.A1(new_n287_), .A2(KEYINPUT23), .ZN(new_n297_));
  NAND3_X1  g160(.A1(new_n285_), .A2(G183gat), .A3(G190gat), .ZN(new_n298_));
  AOI22_X1  g161(.A1(new_n297_), .A2(new_n298_), .B1(new_n271_), .B2(new_n275_), .ZN(new_n299_));
  OAI22_X1  g162(.A1(new_n284_), .A2(new_n289_), .B1(new_n296_), .B2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g163(.A(new_n300_), .B(KEYINPUT30), .ZN(RLL_wire_A_83));
  XOR2_X1 RLL_XOR_83 (.A(RLL_wire_A_83), .B(KEYINPUT83), .Z(new_n301_) );
  XOR2_X1   g164(.A(G15gat), .B(G43gat), .Z(RLL_wire_A_84));
  XOR2_X1 RLL_XOR_84 (.A(RLL_wire_A_84), .B(KEYINPUT84), .Z(new_n302_) );
  NAND2_X1  g165(.A1(G227gat), .A2(G233gat), .ZN(new_n303_));
  XNOR2_X1  g166(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g167(.A(G71gat), .B(G99gat), .ZN(RLL_wire_A_85));
  XOR2_X1 RLL_XOR_85 (.A(RLL_wire_A_85), .B(KEYINPUT85), .Z(new_n305_) );
  XNOR2_X1  g168(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  OR2_X1    g169(.A1(new_n301_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g170(.A1(new_n301_), .A2(new_n306_), .ZN(new_n308_));
  NAND2_X1  g171(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g172(.A(G127gat), .B(G134gat), .ZN(new_n310_));
  XNOR2_X1  g173(.A(G113gat), .B(G120gat), .ZN(new_n311_));
  AND2_X1   g174(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NOR2_X1   g175(.A1(new_n310_), .A2(new_n311_), .ZN(new_n313_));
  NOR2_X1   g176(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g177(.A(new_n314_), .B(KEYINPUT31), .ZN(new_n315_));
  INV_X1    g178(.A(new_n315_), .ZN(new_n316_));
  NAND2_X1  g179(.A1(new_n309_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g180(.A1(new_n307_), .A2(new_n315_), .A3(new_n308_), .ZN(RLL_wire_A_86));
  XOR2_X1 RLL_XOR_86 (.A(RLL_wire_A_86), .B(KEYINPUT86), .Z(new_n318_) );
  NAND2_X1  g181(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g182(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g183(.A1(G141gat), .A2(G148gat), .ZN(new_n321_));
  OR2_X1    g184(.A1(G141gat), .A2(G148gat), .ZN(RLL_wire_A_87));
  XNOR2_X1 RLL_XNOR_87 (.A(RLL_wire_A_87), .B(KEYINPUT87), .ZN(new_n322_) );
  NOR2_X1   g185(.A1(G155gat), .A2(G162gat), .ZN(new_n323_));
  INV_X1    g186(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g187(.A1(G155gat), .A2(G162gat), .ZN(new_n325_));
  NAND2_X1  g188(.A1(new_n325_), .A2(KEYINPUT1), .ZN(new_n326_));
  NAND2_X1  g189(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  NOR2_X1   g190(.A1(new_n325_), .A2(KEYINPUT1), .ZN(new_n328_));
  OAI211_X1 g191(.A(new_n321_), .B(new_n322_), .C1(new_n327_), .C2(new_n328_), .ZN(new_n329_));
  NOR2_X1   g192(.A1(G141gat), .A2(G148gat), .ZN(new_n330_));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n331_));
  NAND2_X1  g194(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g195(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n333_));
  INV_X1    g196(.A(KEYINPUT2), .ZN(new_n334_));
  NAND2_X1  g197(.A1(new_n321_), .A2(new_n334_), .ZN(new_n335_));
  NAND3_X1  g198(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n336_));
  NAND4_X1  g199(.A1(new_n332_), .A2(new_n333_), .A3(new_n335_), .A4(new_n336_), .ZN(new_n337_));
  AND2_X1   g200(.A1(new_n324_), .A2(new_n325_), .ZN(new_n338_));
  NAND2_X1  g201(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g202(.A1(new_n329_), .A2(new_n339_), .ZN(new_n340_));
  NOR2_X1   g203(.A1(new_n340_), .A2(KEYINPUT29), .ZN(new_n341_));
  XOR2_X1   g204(.A(G22gat), .B(G50gat), .Z(new_n342_));
  XNOR2_X1  g205(.A(new_n342_), .B(KEYINPUT28), .ZN(RLL_wire_A_88));
  XOR2_X1 RLL_XOR_88 (.A(RLL_wire_A_88), .B(KEYINPUT88), .Z(new_n343_) );
  XNOR2_X1  g206(.A(new_n341_), .B(new_n343_), .ZN(RLL_wire_A_89));
  XOR2_X1 RLL_XOR_89 (.A(RLL_wire_A_89), .B(KEYINPUT89), .Z(new_n344_) );
  INV_X1    g207(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g208(.A1(new_n340_), .A2(KEYINPUT29), .ZN(new_n346_));
  INV_X1    g209(.A(G228gat), .ZN(new_n347_));
  INV_X1    g210(.A(G233gat), .ZN(new_n348_));
  NOR2_X1   g211(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g212(.A(new_n349_), .ZN(new_n350_));
  INV_X1    g213(.A(G197gat), .ZN(new_n351_));
  NOR2_X1   g214(.A1(new_n351_), .A2(G204gat), .ZN(RLL_wire_A_90));
  XOR2_X1 RLL_XOR_90 (.A(RLL_wire_A_90), .B(KEYINPUT90), .Z(new_n352_) );
  INV_X1    g215(.A(G204gat), .ZN(new_n353_));
  NOR2_X1   g216(.A1(new_n353_), .A2(G197gat), .ZN(new_n354_));
  OAI21_X1  g217(.A(KEYINPUT21), .B1(new_n352_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g218(.A1(new_n353_), .A2(G197gat), .ZN(RLL_wire_A_91));
  XNOR2_X1 RLL_XNOR_91 (.A(RLL_wire_A_91), .B(KEYINPUT91), .ZN(new_n356_) );
  NAND2_X1  g219(.A1(new_n351_), .A2(G204gat), .ZN(new_n357_));
  INV_X1    g220(.A(KEYINPUT21), .ZN(new_n358_));
  NAND3_X1  g221(.A1(new_n356_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g222(.A(G211gat), .B(G218gat), .ZN(new_n360_));
  NAND3_X1  g223(.A1(new_n355_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g224(.A(new_n360_), .ZN(new_n362_));
  NAND2_X1  g225(.A1(new_n356_), .A2(new_n357_), .ZN(new_n363_));
  NAND3_X1  g226(.A1(new_n362_), .A2(KEYINPUT21), .A3(new_n363_), .ZN(RLL_wire_A_92));
  XOR2_X1 RLL_XOR_92 (.A(RLL_wire_A_92), .B(KEYINPUT92), .Z(new_n364_) );
  NAND2_X1  g227(.A1(new_n361_), .A2(new_n364_), .ZN(RLL_wire_A_93));
  XOR2_X1 RLL_XOR_93 (.A(RLL_wire_A_93), .B(KEYINPUT93), .Z(new_n365_) );
  NAND3_X1  g228(.A1(new_n346_), .A2(new_n350_), .A3(new_n365_), .ZN(RLL_wire_A_94));
  XNOR2_X1 RLL_XNOR_94 (.A(RLL_wire_A_94), .B(KEYINPUT94), .ZN(new_n366_) );
  INV_X1    g229(.A(KEYINPUT29), .ZN(new_n367_));
  AOI21_X1  g230(.A(new_n367_), .B1(new_n329_), .B2(new_n339_), .ZN(new_n368_));
  AND2_X1   g231(.A1(new_n361_), .A2(new_n364_), .ZN(new_n369_));
  OAI21_X1  g232(.A(new_n349_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g233(.A(G78gat), .B(G106gat), .ZN(new_n371_));
  INV_X1    g234(.A(new_n371_), .ZN(new_n372_));
  AND3_X1   g235(.A1(new_n366_), .A2(new_n370_), .A3(new_n372_), .ZN(RLL_wire_A_95));
  XNOR2_X1 RLL_XNOR_95 (.A(RLL_wire_A_95), .B(KEYINPUT95), .ZN(new_n373_) );
  AOI21_X1  g236(.A(new_n372_), .B1(new_n366_), .B2(new_n370_), .ZN(RLL_wire_A_96));
  XOR2_X1 RLL_XOR_96 (.A(RLL_wire_A_96), .B(KEYINPUT96), .Z(new_n374_) );
  OAI21_X1  g237(.A(new_n345_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g238(.A1(new_n366_), .A2(new_n370_), .ZN(new_n376_));
  NAND2_X1  g239(.A1(new_n376_), .A2(new_n371_), .ZN(new_n377_));
  NAND3_X1  g240(.A1(new_n366_), .A2(new_n370_), .A3(new_n372_), .ZN(new_n378_));
  NAND3_X1  g241(.A1(new_n377_), .A2(new_n344_), .A3(new_n378_), .ZN(RLL_wire_A_97));
  XOR2_X1 RLL_XOR_97 (.A(RLL_wire_A_97), .B(KEYINPUT97), .Z(new_n379_) );
  NAND2_X1  g242(.A1(new_n375_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g243(.A1(G226gat), .A2(G233gat), .ZN(new_n381_));
  XOR2_X1   g244(.A(new_n381_), .B(KEYINPUT19), .Z(new_n382_));
  INV_X1    g245(.A(new_n382_), .ZN(new_n383_));
  OAI21_X1  g246(.A(KEYINPUT20), .B1(new_n300_), .B2(new_n365_), .ZN(new_n384_));
  XNOR2_X1  g247(.A(KEYINPUT25), .B(G183gat), .ZN(new_n385_));
  XNOR2_X1  g248(.A(KEYINPUT26), .B(G190gat), .ZN(new_n386_));
  INV_X1    g249(.A(KEYINPUT24), .ZN(new_n387_));
  AOI21_X1  g250(.A(new_n387_), .B1(G169gat), .B2(G176gat), .ZN(RLL_wire_A_98));
  XNOR2_X1 RLL_XNOR_98 (.A(RLL_wire_A_98), .B(KEYINPUT98), .ZN(new_n388_) );
  AOI22_X1  g251(.A1(new_n385_), .A2(new_n386_), .B1(new_n388_), .B2(new_n281_), .ZN(new_n389_));
  AOI22_X1  g252(.A1(new_n297_), .A2(new_n298_), .B1(new_n387_), .B2(new_n280_), .ZN(RLL_wire_A_99));
  XNOR2_X1 RLL_XNOR_99 (.A(RLL_wire_A_99), .B(KEYINPUT99), .ZN(new_n390_) );
  NAND2_X1  g253(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g254(.A(new_n282_), .ZN(new_n392_));
  XNOR2_X1  g255(.A(KEYINPUT22), .B(G169gat), .ZN(new_n393_));
  AOI21_X1  g256(.A(new_n392_), .B1(new_n393_), .B2(new_n294_), .ZN(RLL_wire_A_100));
  XNOR2_X1 RLL_XNOR_100 (.A(RLL_wire_A_100), .B(KEYINPUT100), .ZN(new_n394_) );
  OAI22_X1  g257(.A1(new_n286_), .A2(new_n288_), .B1(G183gat), .B2(G190gat), .ZN(new_n395_));
  NAND2_X1  g258(.A1(new_n394_), .A2(new_n395_), .ZN(RLL_wire_A_101));
  XOR2_X1 RLL_XOR_101 (.A(RLL_wire_A_101), .B(KEYINPUT101), .Z(new_n396_) );
  AOI22_X1  g259(.A1(new_n391_), .A2(new_n396_), .B1(new_n364_), .B2(new_n361_), .ZN(new_n397_));
  OAI21_X1  g260(.A(new_n383_), .B1(new_n384_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g261(.A1(new_n300_), .A2(new_n365_), .ZN(new_n399_));
  NAND4_X1  g262(.A1(new_n391_), .A2(new_n396_), .A3(new_n364_), .A4(new_n361_), .ZN(new_n400_));
  NAND4_X1  g263(.A1(new_n399_), .A2(new_n400_), .A3(KEYINPUT20), .A4(new_n382_), .ZN(new_n401_));
  XOR2_X1   g264(.A(G8gat), .B(G36gat), .Z(new_n402_));
  XNOR2_X1  g265(.A(new_n402_), .B(KEYINPUT18), .ZN(new_n403_));
  XNOR2_X1  g266(.A(G64gat), .B(G92gat), .ZN(new_n404_));
  XNOR2_X1  g267(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  AND3_X1   g268(.A1(new_n398_), .A2(new_n401_), .A3(new_n405_), .ZN(new_n406_));
  AOI21_X1  g269(.A(new_n405_), .B1(new_n398_), .B2(new_n401_), .ZN(new_n407_));
  NOR2_X1   g270(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g271(.A1(new_n340_), .A2(new_n314_), .ZN(RLL_wire_A_102));
  XNOR2_X1 RLL_XNOR_102 (.A(RLL_wire_A_102), .B(KEYINPUT102), .ZN(new_n409_) );
  XNOR2_X1  g272(.A(new_n310_), .B(new_n311_), .ZN(new_n410_));
  NAND3_X1  g273(.A1(new_n410_), .A2(new_n329_), .A3(new_n339_), .ZN(new_n411_));
  NAND3_X1  g274(.A1(new_n409_), .A2(new_n411_), .A3(KEYINPUT4), .ZN(new_n412_));
  NAND2_X1  g275(.A1(G225gat), .A2(G233gat), .ZN(new_n413_));
  INV_X1    g276(.A(new_n413_), .ZN(new_n414_));
  INV_X1    g277(.A(KEYINPUT4), .ZN(new_n415_));
  NAND3_X1  g278(.A1(new_n340_), .A2(new_n415_), .A3(new_n314_), .ZN(new_n416_));
  NAND3_X1  g279(.A1(new_n412_), .A2(new_n414_), .A3(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g280(.A(G1gat), .B(G29gat), .ZN(new_n418_));
  XNOR2_X1  g281(.A(new_n418_), .B(KEYINPUT0), .ZN(new_n419_));
  XOR2_X1   g282(.A(G57gat), .B(G85gat), .Z(new_n420_));
  XNOR2_X1  g283(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  NAND3_X1  g284(.A1(new_n409_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n422_));
  NAND4_X1  g285(.A1(new_n417_), .A2(KEYINPUT33), .A3(new_n421_), .A4(new_n422_), .ZN(new_n423_));
  NAND3_X1  g286(.A1(new_n417_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n424_));
  INV_X1    g287(.A(KEYINPUT33), .ZN(new_n425_));
  NAND2_X1  g288(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  AND2_X1   g289(.A1(new_n409_), .A2(new_n411_), .ZN(new_n427_));
  AOI21_X1  g290(.A(new_n421_), .B1(new_n427_), .B2(new_n414_), .ZN(new_n428_));
  NAND3_X1  g291(.A1(new_n412_), .A2(new_n413_), .A3(new_n416_), .ZN(new_n429_));
  NAND2_X1  g292(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND4_X1  g293(.A1(new_n408_), .A2(new_n423_), .A3(new_n426_), .A4(new_n430_), .ZN(new_n431_));
  NAND2_X1  g294(.A1(new_n405_), .A2(KEYINPUT32), .ZN(new_n432_));
  NAND3_X1  g295(.A1(new_n432_), .A2(new_n401_), .A3(new_n398_), .ZN(RLL_wire_A_103));
  XNOR2_X1 RLL_XNOR_103 (.A(RLL_wire_A_103), .B(KEYINPUT103), .ZN(new_n433_) );
  INV_X1    g296(.A(KEYINPUT20), .ZN(new_n434_));
  AOI22_X1  g297(.A1(new_n390_), .A2(new_n389_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n435_));
  AOI21_X1  g298(.A(new_n434_), .B1(new_n369_), .B2(new_n435_), .ZN(RLL_wire_A_104));
  XNOR2_X1 RLL_XNOR_104 (.A(RLL_wire_A_104), .B(KEYINPUT104), .ZN(new_n436_) );
  AOI21_X1  g299(.A(new_n382_), .B1(new_n436_), .B2(new_n399_), .ZN(new_n437_));
  NOR3_X1   g300(.A1(new_n384_), .A2(new_n397_), .A3(new_n383_), .ZN(new_n438_));
  OAI211_X1 g301(.A(KEYINPUT32), .B(new_n405_), .C1(new_n437_), .C2(new_n438_), .ZN(new_n439_));
  AND3_X1   g302(.A1(new_n417_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n440_));
  AOI21_X1  g303(.A(new_n421_), .B1(new_n417_), .B2(new_n422_), .ZN(new_n441_));
  OAI211_X1 g304(.A(new_n433_), .B(new_n439_), .C1(new_n440_), .C2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g305(.A(new_n380_), .B1(new_n431_), .B2(new_n442_), .ZN(new_n443_));
  NOR2_X1   g306(.A1(new_n440_), .A2(new_n441_), .ZN(new_n444_));
  INV_X1    g307(.A(new_n405_), .ZN(new_n445_));
  OAI21_X1  g308(.A(new_n445_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n446_));
  NAND3_X1  g309(.A1(new_n398_), .A2(new_n401_), .A3(new_n405_), .ZN(new_n447_));
  NAND3_X1  g310(.A1(new_n446_), .A2(KEYINPUT27), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g311(.A(KEYINPUT27), .ZN(new_n449_));
  OAI21_X1  g312(.A(new_n449_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n450_));
  AND4_X1   g313(.A1(new_n380_), .A2(new_n444_), .A3(new_n448_), .A4(new_n450_), .ZN(RLL_wire_A_105));
  XOR2_X1 RLL_XOR_105 (.A(RLL_wire_A_105), .B(KEYINPUT105), .Z(new_n451_) );
  OAI21_X1  g314(.A(new_n320_), .B1(new_n443_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g315(.A1(new_n450_), .A2(new_n448_), .ZN(new_n453_));
  NOR2_X1   g316(.A1(new_n453_), .A2(new_n380_), .ZN(new_n454_));
  NAND3_X1  g317(.A1(new_n454_), .A2(new_n444_), .A3(new_n319_), .ZN(RLL_wire_A_106));
  XNOR2_X1 RLL_XNOR_106 (.A(RLL_wire_A_106), .B(KEYINPUT106), .ZN(new_n455_) );
  AOI21_X1  g318(.A(new_n270_), .B1(new_n452_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g319(.A1(new_n253_), .A2(new_n456_), .ZN(RLL_wire_A_107));
  XOR2_X1 RLL_XOR_107 (.A(RLL_wire_A_107), .B(KEYINPUT107), .Z(new_n457_) );
  INV_X1    g320(.A(new_n457_), .ZN(new_n458_));
  INV_X1    g321(.A(new_n444_), .ZN(new_n459_));
  NAND3_X1  g322(.A1(new_n458_), .A2(new_n231_), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g323(.A(KEYINPUT38), .ZN(new_n461_));
  OR2_X1    g324(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g325(.A1(new_n195_), .A2(new_n269_), .ZN(new_n463_));
  NOR2_X1   g326(.A1(new_n463_), .A2(new_n250_), .ZN(new_n464_));
  NAND2_X1  g327(.A1(new_n226_), .A2(new_n219_), .ZN(new_n465_));
  INV_X1    g328(.A(new_n465_), .ZN(RLL_wire_A_108));
  XOR2_X1 RLL_XOR_108 (.A(RLL_wire_A_108), .B(KEYINPUT108), .Z(new_n466_) );
  AOI21_X1  g329(.A(new_n466_), .B1(new_n452_), .B2(new_n455_), .ZN(new_n467_));
  NAND2_X1  g330(.A1(new_n464_), .A2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g331(.A(G1gat), .B1(new_n468_), .B2(new_n444_), .ZN(new_n469_));
  NAND2_X1  g332(.A1(new_n460_), .A2(new_n461_), .ZN(new_n470_));
  NAND3_X1  g333(.A1(new_n462_), .A2(new_n469_), .A3(new_n470_), .ZN(G1324gat));
  NAND3_X1  g334(.A1(new_n458_), .A2(new_n232_), .A3(new_n453_), .ZN(new_n472_));
  NAND3_X1  g335(.A1(new_n464_), .A2(new_n453_), .A3(new_n467_), .ZN(RLL_wire_A_109));
  XOR2_X1 RLL_XOR_109 (.A(RLL_wire_A_109), .B(KEYINPUT109), .Z(new_n473_) );
  NAND2_X1  g336(.A1(new_n473_), .A2(G8gat), .ZN(new_n474_));
  AND2_X1   g337(.A1(new_n474_), .A2(KEYINPUT39), .ZN(new_n475_));
  NOR2_X1   g338(.A1(new_n474_), .A2(KEYINPUT39), .ZN(new_n476_));
  OAI21_X1  g339(.A(new_n472_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g340(.A(KEYINPUT40), .ZN(new_n478_));
  XNOR2_X1  g341(.A(new_n477_), .B(new_n478_), .ZN(G1325gat));
  OAI21_X1  g342(.A(G15gat), .B1(new_n468_), .B2(new_n320_), .ZN(RLL_wire_A_110));
  XNOR2_X1 RLL_XNOR_110 (.A(RLL_wire_A_110), .B(KEYINPUT110), .ZN(new_n480_) );
  XNOR2_X1  g343(.A(new_n480_), .B(KEYINPUT41), .ZN(new_n481_));
  NOR3_X1   g344(.A1(new_n457_), .A2(G15gat), .A3(new_n320_), .ZN(new_n482_));
  OR2_X1    g345(.A1(new_n481_), .A2(new_n482_), .ZN(G1326gat));
  INV_X1    g346(.A(new_n380_), .ZN(new_n484_));
  OAI21_X1  g347(.A(G22gat), .B1(new_n468_), .B2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g348(.A(new_n485_), .B(KEYINPUT42), .ZN(new_n486_));
  OR2_X1    g349(.A1(new_n484_), .A2(G22gat), .ZN(new_n487_));
  OAI21_X1  g350(.A(new_n486_), .B1(new_n457_), .B2(new_n487_), .ZN(G1327gat));
  NOR2_X1   g351(.A1(new_n463_), .A2(new_n251_), .ZN(new_n489_));
  INV_X1    g352(.A(KEYINPUT43), .ZN(new_n490_));
  NAND2_X1  g353(.A1(new_n452_), .A2(new_n455_), .ZN(new_n491_));
  INV_X1    g354(.A(new_n229_), .ZN(new_n492_));
  AOI21_X1  g355(.A(new_n490_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  AOI211_X1 g356(.A(KEYINPUT43), .B(new_n229_), .C1(new_n452_), .C2(new_n455_), .ZN(new_n494_));
  OAI21_X1  g357(.A(new_n489_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g358(.A(KEYINPUT44), .ZN(new_n496_));
  NAND2_X1  g359(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  OAI211_X1 g360(.A(KEYINPUT44), .B(new_n489_), .C1(new_n493_), .C2(new_n494_), .ZN(new_n498_));
  NAND3_X1  g361(.A1(new_n497_), .A2(new_n459_), .A3(new_n498_), .ZN(RLL_wire_A_111));
  XOR2_X1 RLL_XOR_111 (.A(RLL_wire_A_111), .B(KEYINPUT111), .Z(new_n499_) );
  NAND2_X1  g362(.A1(new_n499_), .A2(G29gat), .ZN(new_n500_));
  NOR2_X1   g363(.A1(new_n465_), .A2(new_n251_), .ZN(new_n501_));
  NAND3_X1  g364(.A1(new_n456_), .A2(new_n195_), .A3(new_n501_), .ZN(new_n502_));
  OR2_X1    g365(.A1(new_n444_), .A2(G29gat), .ZN(new_n503_));
  OAI21_X1  g366(.A(new_n500_), .B1(new_n502_), .B2(new_n503_), .ZN(G1328gat));
  NAND3_X1  g367(.A1(new_n497_), .A2(new_n453_), .A3(new_n498_), .ZN(new_n505_));
  NAND2_X1  g368(.A1(new_n505_), .A2(G36gat), .ZN(RLL_wire_A_112));
  XNOR2_X1 RLL_XNOR_112 (.A(RLL_wire_A_112), .B(KEYINPUT112), .ZN(new_n506_) );
  INV_X1    g369(.A(new_n453_), .ZN(new_n507_));
  NOR3_X1   g370(.A1(new_n502_), .A2(G36gat), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g371(.A(KEYINPUT45), .ZN(new_n509_));
  XNOR2_X1  g372(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  NAND2_X1  g373(.A1(new_n506_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g374(.A(KEYINPUT46), .ZN(new_n512_));
  NAND2_X1  g375(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g376(.A1(new_n506_), .A2(KEYINPUT46), .A3(new_n510_), .ZN(new_n514_));
  NAND2_X1  g377(.A1(new_n513_), .A2(new_n514_), .ZN(G1329gat));
  NAND4_X1  g378(.A1(new_n497_), .A2(G43gat), .A3(new_n319_), .A4(new_n498_), .ZN(new_n516_));
  INV_X1    g379(.A(G43gat), .ZN(new_n517_));
  OAI21_X1  g380(.A(new_n517_), .B1(new_n502_), .B2(new_n320_), .ZN(new_n518_));
  NAND2_X1  g381(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g382(.A(new_n519_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g383(.A1(new_n497_), .A2(new_n380_), .A3(new_n498_), .ZN(new_n521_));
  NAND2_X1  g384(.A1(new_n521_), .A2(G50gat), .ZN(new_n522_));
  OR2_X1    g385(.A1(new_n484_), .A2(G50gat), .ZN(new_n523_));
  OAI21_X1  g386(.A(new_n522_), .B1(new_n502_), .B2(new_n523_), .ZN(G1331gat));
  NOR2_X1   g387(.A1(new_n252_), .A2(new_n195_), .ZN(new_n525_));
  AOI21_X1  g388(.A(new_n269_), .B1(new_n452_), .B2(new_n455_), .ZN(new_n526_));
  NAND2_X1  g389(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g390(.A(new_n527_), .ZN(RLL_wire_A_113));
  XNOR2_X1 RLL_XNOR_113 (.A(RLL_wire_A_113), .B(KEYINPUT113), .ZN(new_n528_) );
  AOI21_X1  g391(.A(G57gat), .B1(new_n528_), .B2(new_n459_), .ZN(new_n529_));
  NAND4_X1  g392(.A1(new_n467_), .A2(new_n270_), .A3(new_n196_), .A4(new_n251_), .ZN(new_n530_));
  INV_X1    g393(.A(G57gat), .ZN(new_n531_));
  NOR3_X1   g394(.A1(new_n530_), .A2(new_n531_), .A3(new_n444_), .ZN(new_n532_));
  NOR2_X1   g395(.A1(new_n529_), .A2(new_n532_), .ZN(RLL_wire_A_114));
  XOR2_X1 RLL_XOR_114 (.A(RLL_wire_A_114), .B(KEYINPUT114), .Z(G1332gat) );
  OAI21_X1  g396(.A(G64gat), .B1(new_n530_), .B2(new_n507_), .ZN(new_n534_));
  XNOR2_X1  g397(.A(new_n534_), .B(KEYINPUT48), .ZN(new_n535_));
  OR2_X1    g398(.A1(new_n507_), .A2(G64gat), .ZN(new_n536_));
  OAI21_X1  g399(.A(new_n535_), .B1(new_n527_), .B2(new_n536_), .ZN(G1333gat));
  OAI21_X1  g400(.A(G71gat), .B1(new_n530_), .B2(new_n320_), .ZN(new_n538_));
  XNOR2_X1  g401(.A(new_n538_), .B(KEYINPUT49), .ZN(new_n539_));
  OR2_X1    g402(.A1(new_n320_), .A2(G71gat), .ZN(new_n540_));
  OAI21_X1  g403(.A(new_n539_), .B1(new_n527_), .B2(new_n540_), .ZN(G1334gat));
  OAI21_X1  g404(.A(G78gat), .B1(new_n530_), .B2(new_n484_), .ZN(RLL_wire_A_115));
  XNOR2_X1 RLL_XNOR_115 (.A(RLL_wire_A_115), .B(KEYINPUT115), .ZN(new_n542_) );
  XNOR2_X1  g405(.A(new_n542_), .B(KEYINPUT50), .ZN(new_n543_));
  OR2_X1    g406(.A1(new_n484_), .A2(G78gat), .ZN(new_n544_));
  OAI21_X1  g407(.A(new_n543_), .B1(new_n527_), .B2(new_n544_), .ZN(G1335gat));
  AND3_X1   g408(.A1(new_n526_), .A2(new_n196_), .A3(new_n501_), .ZN(new_n546_));
  AOI21_X1  g409(.A(G85gat), .B1(new_n546_), .B2(new_n459_), .ZN(new_n547_));
  OR2_X1    g410(.A1(new_n493_), .A2(new_n494_), .ZN(new_n548_));
  NOR3_X1   g411(.A1(new_n195_), .A2(new_n269_), .A3(new_n251_), .ZN(new_n549_));
  NAND2_X1  g412(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g413(.A(new_n550_), .ZN(new_n551_));
  NOR2_X1   g414(.A1(new_n444_), .A2(new_n144_), .ZN(RLL_wire_A_116));
  XNOR2_X1 RLL_XNOR_116 (.A(RLL_wire_A_116), .B(KEYINPUT116), .ZN(new_n552_) );
  AOI21_X1  g415(.A(new_n547_), .B1(new_n551_), .B2(new_n552_), .ZN(G1336gat));
  AOI21_X1  g416(.A(G92gat), .B1(new_n546_), .B2(new_n453_), .ZN(new_n554_));
  NOR2_X1   g417(.A1(new_n507_), .A2(new_n145_), .ZN(new_n555_));
  AOI21_X1  g418(.A(new_n554_), .B1(new_n551_), .B2(new_n555_), .ZN(G1337gat));
  OAI21_X1  g419(.A(G99gat), .B1(new_n550_), .B2(new_n320_), .ZN(new_n557_));
  NAND3_X1  g420(.A1(new_n546_), .A2(new_n319_), .A3(new_n140_), .ZN(RLL_wire_A_117));
  XOR2_X1 RLL_XOR_117 (.A(RLL_wire_A_117), .B(KEYINPUT117), .Z(new_n558_) );
  NAND2_X1  g421(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g422(.A1(new_n559_), .A2(KEYINPUT51), .ZN(RLL_wire_A_118));
  XOR2_X1 RLL_XOR_118 (.A(RLL_wire_A_118), .B(KEYINPUT118), .Z(new_n560_) );
  INV_X1    g423(.A(KEYINPUT51), .ZN(new_n561_));
  NAND3_X1  g424(.A1(new_n557_), .A2(new_n561_), .A3(new_n558_), .ZN(new_n562_));
  NAND2_X1  g425(.A1(new_n560_), .A2(new_n562_), .ZN(G1338gat));
  NAND3_X1  g426(.A1(new_n546_), .A2(new_n141_), .A3(new_n380_), .ZN(new_n564_));
  OAI211_X1 g427(.A(new_n380_), .B(new_n549_), .C1(new_n493_), .C2(new_n494_), .ZN(new_n565_));
  INV_X1    g428(.A(KEYINPUT52), .ZN(new_n566_));
  AND3_X1   g429(.A1(new_n565_), .A2(new_n566_), .A3(G106gat), .ZN(new_n567_));
  AOI21_X1  g430(.A(new_n566_), .B1(new_n565_), .B2(G106gat), .ZN(new_n568_));
  OAI21_X1  g431(.A(new_n564_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g432(.A(new_n569_), .B(KEYINPUT53), .ZN(RLL_wire_A_119));
  XNOR2_X1 RLL_XNOR_119 (.A(RLL_wire_A_119), .B(KEYINPUT119), .ZN(G1339gat) );
  NAND2_X1  g433(.A1(new_n251_), .A2(new_n270_), .ZN(RLL_wire_A_120));
  XNOR2_X1 RLL_XNOR_120 (.A(RLL_wire_A_120), .B(KEYINPUT120), .ZN(new_n571_) );
  AOI21_X1  g434(.A(new_n571_), .B1(new_n193_), .B2(new_n194_), .ZN(new_n572_));
  INV_X1    g435(.A(KEYINPUT54), .ZN(new_n573_));
  AND3_X1   g436(.A1(new_n572_), .A2(new_n573_), .A3(new_n229_), .ZN(new_n574_));
  AOI21_X1  g437(.A(new_n573_), .B1(new_n572_), .B2(new_n229_), .ZN(new_n575_));
  NOR2_X1   g438(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g439(.A1(new_n269_), .A2(new_n191_), .ZN(new_n577_));
  INV_X1    g440(.A(KEYINPUT55), .ZN(new_n578_));
  NAND2_X1  g441(.A1(new_n183_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g442(.A1(new_n179_), .A2(new_n181_), .A3(new_n171_), .ZN(new_n580_));
  NAND2_X1  g443(.A1(new_n580_), .A2(new_n139_), .ZN(new_n581_));
  NAND4_X1  g444(.A1(new_n179_), .A2(new_n181_), .A3(new_n182_), .A4(KEYINPUT55), .ZN(new_n582_));
  NAND3_X1  g445(.A1(new_n579_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  NAND2_X1  g446(.A1(new_n583_), .A2(new_n189_), .ZN(new_n584_));
  INV_X1    g447(.A(KEYINPUT56), .ZN(new_n585_));
  NAND2_X1  g448(.A1(new_n584_), .A2(new_n585_), .ZN(RLL_wire_A_121));
  XNOR2_X1 RLL_XNOR_121 (.A(RLL_wire_A_121), .B(KEYINPUT121), .ZN(new_n586_) );
  NAND3_X1  g449(.A1(new_n583_), .A2(KEYINPUT56), .A3(new_n189_), .ZN(new_n587_));
  AOI21_X1  g450(.A(new_n577_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  AOI21_X1  g451(.A(new_n265_), .B1(new_n257_), .B2(new_n260_), .ZN(new_n589_));
  NAND2_X1  g452(.A1(new_n259_), .A2(new_n255_), .ZN(new_n590_));
  OAI21_X1  g453(.A(new_n589_), .B1(new_n590_), .B2(new_n260_), .ZN(new_n591_));
  AND2_X1   g454(.A1(new_n591_), .A2(new_n268_), .ZN(new_n592_));
  AND2_X1   g455(.A1(new_n192_), .A2(new_n592_), .ZN(new_n593_));
  OAI21_X1  g456(.A(new_n465_), .B1(new_n588_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g457(.A(KEYINPUT57), .ZN(new_n595_));
  NAND2_X1  g458(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  AND2_X1   g459(.A1(new_n592_), .A2(new_n191_), .ZN(new_n597_));
  AND3_X1   g460(.A1(new_n583_), .A2(KEYINPUT56), .A3(new_n189_), .ZN(new_n598_));
  AOI21_X1  g461(.A(KEYINPUT56), .B1(new_n583_), .B2(new_n189_), .ZN(new_n599_));
  OAI21_X1  g462(.A(new_n597_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g463(.A(KEYINPUT58), .ZN(new_n601_));
  AOI21_X1  g464(.A(new_n229_), .B1(new_n600_), .B2(new_n601_), .ZN(RLL_wire_A_122));
  XOR2_X1 RLL_XOR_122 (.A(RLL_wire_A_122), .B(KEYINPUT122), .Z(new_n602_) );
  OAI211_X1 g465(.A(KEYINPUT58), .B(new_n597_), .C1(new_n598_), .C2(new_n599_), .ZN(new_n603_));
  NAND2_X1  g466(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  OAI211_X1 g467(.A(new_n465_), .B(KEYINPUT57), .C1(new_n588_), .C2(new_n593_), .ZN(RLL_wire_A_123));
  XOR2_X1 RLL_XOR_123 (.A(RLL_wire_A_123), .B(KEYINPUT123), .Z(new_n605_) );
  NAND3_X1  g468(.A1(new_n596_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n606_));
  AOI21_X1  g469(.A(new_n576_), .B1(new_n606_), .B2(new_n250_), .ZN(new_n607_));
  NAND3_X1  g470(.A1(new_n454_), .A2(new_n459_), .A3(new_n319_), .ZN(new_n608_));
  NOR2_X1   g471(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  AOI21_X1  g472(.A(G113gat), .B1(new_n609_), .B2(new_n269_), .ZN(new_n610_));
  OAI21_X1  g473(.A(KEYINPUT59), .B1(new_n607_), .B2(new_n608_), .ZN(new_n611_));
  INV_X1    g474(.A(KEYINPUT59), .ZN(new_n612_));
  INV_X1    g475(.A(new_n608_), .ZN(new_n613_));
  AOI22_X1  g476(.A1(new_n595_), .A2(new_n594_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n614_));
  AOI21_X1  g477(.A(new_n251_), .B1(new_n614_), .B2(new_n605_), .ZN(new_n615_));
  OAI211_X1 g478(.A(new_n612_), .B(new_n613_), .C1(new_n615_), .C2(new_n576_), .ZN(new_n616_));
  AND2_X1   g479(.A1(new_n611_), .A2(new_n616_), .ZN(RLL_wire_A_124));
  XNOR2_X1 RLL_XNOR_124 (.A(RLL_wire_A_124), .B(KEYINPUT124), .ZN(new_n617_) );
  INV_X1    g480(.A(G113gat), .ZN(new_n618_));
  NOR2_X1   g481(.A1(new_n270_), .A2(new_n618_), .ZN(new_n619_));
  AOI21_X1  g482(.A(new_n610_), .B1(new_n617_), .B2(new_n619_), .ZN(G1340gat));
  INV_X1    g483(.A(G120gat), .ZN(new_n621_));
  OAI21_X1  g484(.A(new_n621_), .B1(new_n195_), .B2(KEYINPUT60), .ZN(RLL_wire_A_125));
  XOR2_X1 RLL_XOR_125 (.A(RLL_wire_A_125), .B(KEYINPUT125), .Z(new_n622_) );
  OAI211_X1 g485(.A(new_n609_), .B(new_n622_), .C1(KEYINPUT60), .C2(new_n621_), .ZN(new_n623_));
  AND3_X1   g486(.A1(new_n611_), .A2(new_n196_), .A3(new_n616_), .ZN(new_n624_));
  OAI21_X1  g487(.A(new_n623_), .B1(new_n624_), .B2(new_n621_), .ZN(G1341gat));
  AOI21_X1  g488(.A(G127gat), .B1(new_n609_), .B2(new_n251_), .ZN(new_n626_));
  INV_X1    g489(.A(G127gat), .ZN(new_n627_));
  NOR2_X1   g490(.A1(new_n250_), .A2(new_n627_), .ZN(new_n628_));
  AOI21_X1  g491(.A(new_n626_), .B1(new_n617_), .B2(new_n628_), .ZN(G1342gat));
  AOI21_X1  g492(.A(G134gat), .B1(new_n609_), .B2(new_n466_), .ZN(new_n630_));
  INV_X1    g493(.A(G134gat), .ZN(new_n631_));
  NOR2_X1   g494(.A1(new_n229_), .A2(new_n631_), .ZN(new_n632_));
  AOI21_X1  g495(.A(new_n630_), .B1(new_n617_), .B2(new_n632_), .ZN(G1343gat));
  NAND4_X1  g496(.A1(new_n507_), .A2(new_n320_), .A3(new_n380_), .A4(new_n459_), .ZN(new_n634_));
  NOR2_X1   g497(.A1(new_n607_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g498(.A1(new_n635_), .A2(new_n269_), .ZN(new_n636_));
  XNOR2_X1  g499(.A(new_n636_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g500(.A1(new_n635_), .A2(new_n196_), .ZN(new_n638_));
  XNOR2_X1  g501(.A(new_n638_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g502(.A1(new_n635_), .A2(new_n251_), .ZN(new_n640_));
  XNOR2_X1  g503(.A(KEYINPUT61), .B(G155gat), .ZN(new_n641_));
  XNOR2_X1  g504(.A(new_n640_), .B(new_n641_), .ZN(G1346gat));
  AOI21_X1  g505(.A(G162gat), .B1(new_n635_), .B2(new_n466_), .ZN(new_n643_));
  AND2_X1   g506(.A1(new_n492_), .A2(G162gat), .ZN(new_n644_));
  AOI21_X1  g507(.A(new_n643_), .B1(new_n635_), .B2(new_n644_), .ZN(G1347gat));
  NOR3_X1   g508(.A1(new_n507_), .A2(new_n320_), .A3(new_n459_), .ZN(new_n646_));
  AND2_X1   g509(.A1(new_n646_), .A2(new_n269_), .ZN(RLL_wire_A_126));
  XOR2_X1 RLL_XOR_126 (.A(RLL_wire_A_126), .B(KEYINPUT126), .Z(new_n647_) );
  OAI211_X1 g510(.A(new_n484_), .B(new_n647_), .C1(new_n615_), .C2(new_n576_), .ZN(new_n648_));
  INV_X1    g511(.A(KEYINPUT62), .ZN(new_n649_));
  AND3_X1   g512(.A1(new_n648_), .A2(new_n649_), .A3(G169gat), .ZN(new_n650_));
  AOI21_X1  g513(.A(new_n649_), .B1(new_n648_), .B2(G169gat), .ZN(new_n651_));
  OAI211_X1 g514(.A(new_n484_), .B(new_n646_), .C1(new_n615_), .C2(new_n576_), .ZN(new_n652_));
  NAND2_X1  g515(.A1(new_n269_), .A2(new_n393_), .ZN(new_n653_));
  OAI22_X1  g516(.A1(new_n650_), .A2(new_n651_), .B1(new_n652_), .B2(new_n653_), .ZN(G1348gat));
  OAI21_X1  g517(.A(new_n294_), .B1(new_n652_), .B2(new_n195_), .ZN(new_n655_));
  NOR2_X1   g518(.A1(new_n607_), .A2(new_n380_), .ZN(new_n656_));
  NAND4_X1  g519(.A1(new_n656_), .A2(G176gat), .A3(new_n196_), .A4(new_n646_), .ZN(new_n657_));
  AND2_X1   g520(.A1(new_n655_), .A2(new_n657_), .ZN(G1349gat));
  NOR3_X1   g521(.A1(new_n652_), .A2(new_n385_), .A3(new_n250_), .ZN(new_n659_));
  NAND3_X1  g522(.A1(new_n656_), .A2(new_n251_), .A3(new_n646_), .ZN(new_n660_));
  AOI21_X1  g523(.A(new_n659_), .B1(new_n271_), .B2(new_n660_), .ZN(G1350gat));
  OAI21_X1  g524(.A(G190gat), .B1(new_n652_), .B2(new_n229_), .ZN(new_n662_));
  NAND2_X1  g525(.A1(new_n466_), .A2(new_n386_), .ZN(RLL_wire_A_127));
  XOR2_X1 RLL_XOR_127 (.A(RLL_wire_A_127), .B(KEYINPUT127), .Z(new_n663_) );
  OAI21_X1  g526(.A(new_n662_), .B1(new_n652_), .B2(new_n663_), .ZN(G1351gat));
  NAND3_X1  g527(.A1(new_n320_), .A2(new_n380_), .A3(new_n444_), .ZN(new_n665_));
  NOR3_X1   g528(.A1(new_n607_), .A2(new_n507_), .A3(new_n665_), .ZN(new_n666_));
  AND3_X1   g529(.A1(new_n666_), .A2(G197gat), .A3(new_n269_), .ZN(new_n667_));
  AOI21_X1  g530(.A(G197gat), .B1(new_n666_), .B2(new_n269_), .ZN(new_n668_));
  NOR2_X1   g531(.A1(new_n667_), .A2(new_n668_), .ZN(G1352gat));
  NAND2_X1  g532(.A1(new_n666_), .A2(new_n196_), .ZN(new_n670_));
  NAND2_X1  g533(.A1(new_n670_), .A2(G204gat), .ZN(new_n671_));
  NAND3_X1  g534(.A1(new_n666_), .A2(new_n353_), .A3(new_n196_), .ZN(new_n672_));
  NAND2_X1  g535(.A1(new_n671_), .A2(new_n672_), .ZN(G1353gat));
  AOI21_X1  g536(.A(new_n250_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n674_));
  OR2_X1    g537(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n675_));
  AND3_X1   g538(.A1(new_n666_), .A2(new_n674_), .A3(new_n675_), .ZN(new_n676_));
  AOI21_X1  g539(.A(new_n675_), .B1(new_n666_), .B2(new_n674_), .ZN(new_n677_));
  NOR2_X1   g540(.A1(new_n676_), .A2(new_n677_), .ZN(G1354gat));
  NAND2_X1  g541(.A1(new_n666_), .A2(new_n466_), .ZN(new_n679_));
  INV_X1    g542(.A(G218gat), .ZN(new_n680_));
  NOR2_X1   g543(.A1(new_n229_), .A2(new_n680_), .ZN(new_n681_));
  AOI22_X1  g544(.A1(new_n679_), .A2(new_n680_), .B1(new_n666_), .B2(new_n681_), .ZN(G1355gat));

endmodule
