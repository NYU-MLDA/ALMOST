//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n854_, new_n856_, new_n857_,
    new_n859_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n904_, new_n905_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_;
  INV_X1    g000(.A(KEYINPUT66), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT65), .ZN(new_n203_));
  INV_X1    g002(.A(G64gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G57gat), .ZN(new_n205_));
  INV_X1    g004(.A(G57gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G64gat), .ZN(new_n207_));
  AOI21_X1  g006(.A(KEYINPUT11), .B1(new_n205_), .B2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G71gat), .B(G78gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n203_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  AND2_X1   g009(.A1(G71gat), .A2(G78gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G71gat), .A2(G78gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G57gat), .B(G64gat), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n213_), .B(KEYINPUT65), .C1(new_n214_), .C2(KEYINPUT11), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(KEYINPUT11), .ZN(new_n216_));
  AND3_X1   g015(.A1(new_n210_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n216_), .B1(new_n210_), .B2(new_n215_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT7), .ZN(new_n220_));
  INV_X1    g019(.A(G99gat), .ZN(new_n221_));
  INV_X1    g020(.A(G106gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G99gat), .A2(G106gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT6), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n223_), .A2(new_n226_), .A3(new_n227_), .A4(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230_));
  INV_X1    g029(.A(G85gat), .ZN(new_n231_));
  INV_X1    g030(.A(G92gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(G85gat), .A2(G92gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n229_), .A2(new_n230_), .A3(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n230_), .B1(new_n229_), .B2(new_n235_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n226_), .A2(new_n227_), .ZN(new_n239_));
  XOR2_X1   g038(.A(KEYINPUT10), .B(G99gat), .Z(new_n240_));
  AOI21_X1  g039(.A(new_n239_), .B1(new_n240_), .B2(new_n222_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n243_), .B1(G85gat), .B2(G92gat), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n232_), .A2(KEYINPUT64), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n232_), .A2(KEYINPUT64), .ZN(new_n246_));
  OAI21_X1  g045(.A(G85gat), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT9), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n244_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  OAI22_X1  g048(.A1(new_n237_), .A2(new_n238_), .B1(new_n242_), .B2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n202_), .B1(new_n219_), .B2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n219_), .A2(new_n250_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n210_), .A2(new_n215_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n216_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n210_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n238_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n244_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT64), .B(G92gat), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n260_), .A2(new_n231_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n259_), .B1(new_n261_), .B2(KEYINPUT9), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n258_), .A2(new_n236_), .B1(new_n262_), .B2(new_n241_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n257_), .A2(new_n263_), .A3(KEYINPUT66), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n251_), .A2(new_n252_), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G230gat), .A2(G233gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n267_), .B1(new_n257_), .B2(new_n263_), .ZN(new_n269_));
  NOR3_X1   g068(.A1(new_n257_), .A2(new_n263_), .A3(KEYINPUT12), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT12), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n271_), .B1(new_n219_), .B2(new_n250_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n269_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n268_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G120gat), .B(G148gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT5), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G176gat), .B(G204gat), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n276_), .B(new_n277_), .Z(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n278_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n268_), .A2(new_n273_), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n282_), .A2(KEYINPUT13), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n283_), .B(KEYINPUT67), .Z(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(KEYINPUT13), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n285_), .B(KEYINPUT68), .Z(new_n286_));
  NOR2_X1   g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n287_), .A2(KEYINPUT69), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(KEYINPUT69), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT76), .B(G1gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(G8gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT14), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G15gat), .B(G22gat), .ZN(new_n294_));
  XOR2_X1   g093(.A(G1gat), .B(G8gat), .Z(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n293_), .A2(new_n294_), .A3(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT14), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n298_), .B1(new_n291_), .B2(G8gat), .ZN(new_n299_));
  INV_X1    g098(.A(new_n294_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n295_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n297_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G29gat), .B(G36gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G43gat), .B(G50gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n305_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n307_), .A2(new_n297_), .A3(new_n301_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G229gat), .A2(G233gat), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n307_), .A2(KEYINPUT15), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT15), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n305_), .A2(new_n314_), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n313_), .A2(new_n297_), .A3(new_n315_), .A4(new_n301_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n306_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n310_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G113gat), .B(G141gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G169gat), .B(G197gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n312_), .A2(new_n318_), .A3(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n321_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n310_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n324_), .B1(new_n316_), .B2(new_n306_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n323_), .B1(new_n325_), .B2(new_n311_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n322_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G8gat), .B(G36gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT18), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G64gat), .B(G92gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G226gat), .A2(G233gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G211gat), .B(G218gat), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT86), .ZN(new_n336_));
  INV_X1    g135(.A(G197gat), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n336_), .B1(new_n337_), .B2(G204gat), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n335_), .A2(KEYINPUT21), .A3(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G197gat), .B(G204gat), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n340_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n335_), .A2(KEYINPUT21), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G169gat), .A2(G176gat), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT22), .B(G169gat), .ZN(new_n348_));
  INV_X1    g147(.A(G176gat), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n347_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n350_), .B(KEYINPUT92), .Z(new_n351_));
  NAND2_X1  g150(.A1(G183gat), .A2(G190gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT23), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT79), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT79), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n352_), .A2(new_n355_), .A3(KEYINPUT23), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT23), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n357_), .A2(G183gat), .A3(G190gat), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n354_), .A2(new_n356_), .A3(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n359_), .B1(G183gat), .B2(G190gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n351_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT90), .B(KEYINPUT24), .ZN(new_n362_));
  OR3_X1    g161(.A1(new_n362_), .A2(KEYINPUT91), .A3(new_n347_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT91), .B1(new_n362_), .B2(new_n347_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n363_), .B(new_n364_), .C1(G169gat), .C2(G176gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n353_), .A2(new_n358_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(G169gat), .A2(G176gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n362_), .A2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT26), .B(G190gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT25), .B(G183gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n365_), .A2(new_n366_), .A3(new_n368_), .A4(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n345_), .B1(new_n361_), .B2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n346_), .A2(KEYINPUT24), .ZN(new_n374_));
  MUX2_X1   g173(.A(new_n374_), .B(KEYINPUT24), .S(new_n367_), .Z(new_n375_));
  INV_X1    g174(.A(new_n369_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT78), .B(G183gat), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n377_), .B1(new_n378_), .B2(KEYINPUT25), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n375_), .B(new_n359_), .C1(new_n376_), .C2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n366_), .B1(new_n378_), .B2(G190gat), .ZN(new_n381_));
  AOI21_X1  g180(.A(G176gat), .B1(KEYINPUT80), .B2(KEYINPUT22), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(G169gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n380_), .A2(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n385_), .A2(new_n344_), .ZN(new_n386_));
  OAI211_X1 g185(.A(KEYINPUT20), .B(new_n334_), .C1(new_n373_), .C2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT20), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n361_), .A2(new_n372_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n389_), .B1(new_n390_), .B2(new_n345_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n345_), .A2(new_n385_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n334_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n331_), .B1(new_n388_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n331_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n344_), .B1(new_n361_), .B2(new_n372_), .ZN(new_n397_));
  NOR3_X1   g196(.A1(new_n397_), .A2(new_n392_), .A3(new_n389_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n387_), .B(new_n396_), .C1(new_n398_), .C2(new_n334_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n395_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT27), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(G155gat), .A2(G162gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G155gat), .A2(G162gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(G141gat), .A2(G148gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT3), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G141gat), .A2(G148gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT2), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n406_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n405_), .A2(KEYINPUT1), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n405_), .A2(KEYINPUT1), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(new_n414_), .A3(new_n404_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n407_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n415_), .A2(new_n409_), .A3(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n412_), .A2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G127gat), .B(G134gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G113gat), .B(G120gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n418_), .A2(new_n422_), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n415_), .A2(new_n409_), .A3(new_n416_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n424_), .A2(new_n411_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(new_n421_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n423_), .A2(new_n426_), .A3(KEYINPUT4), .ZN(new_n427_));
  OR3_X1    g226(.A1(new_n425_), .A2(KEYINPUT4), .A3(new_n421_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G225gat), .A2(G233gat), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n427_), .A2(new_n428_), .A3(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n423_), .A2(new_n426_), .A3(new_n429_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G1gat), .B(G29gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT0), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(new_n206_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(G85gat), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n431_), .A2(new_n432_), .A3(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT94), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n431_), .A2(new_n436_), .A3(KEYINPUT94), .A4(new_n432_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n431_), .A2(new_n432_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n435_), .B(new_n231_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n439_), .A2(new_n440_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n334_), .ZN(new_n445_));
  OAI211_X1 g244(.A(KEYINPUT20), .B(new_n445_), .C1(new_n373_), .C2(new_n386_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n446_), .B(new_n331_), .C1(new_n398_), .C2(new_n445_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n399_), .A2(new_n447_), .A3(KEYINPUT27), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n402_), .A2(new_n444_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT87), .ZN(new_n450_));
  INV_X1    g249(.A(G233gat), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n451_), .A2(KEYINPUT85), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(KEYINPUT85), .ZN(new_n453_));
  OAI21_X1  g252(.A(G228gat), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT29), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n456_), .B1(new_n412_), .B2(new_n417_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n455_), .B1(new_n457_), .B2(new_n344_), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT29), .B1(new_n424_), .B2(new_n411_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n345_), .A2(new_n459_), .A3(new_n454_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G78gat), .B(G106gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n462_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n458_), .A2(new_n460_), .A3(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n450_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT83), .B1(new_n418_), .B2(KEYINPUT29), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G22gat), .B(G50gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT28), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT83), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n425_), .A2(new_n470_), .A3(new_n456_), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n467_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n469_), .B1(new_n467_), .B2(new_n471_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT88), .B1(new_n466_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n465_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n464_), .B1(new_n458_), .B2(new_n460_), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT87), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n474_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT88), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n463_), .A2(new_n465_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT84), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT87), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n475_), .A2(new_n481_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n484_), .B1(new_n475_), .B2(new_n481_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT30), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n385_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n380_), .A2(KEYINPUT30), .A3(new_n384_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G15gat), .B(G43gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G71gat), .B(G99gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G227gat), .A2(G233gat), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n495_), .B(KEYINPUT81), .Z(new_n496_));
  XNOR2_X1  g295(.A(new_n494_), .B(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n491_), .B(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT82), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n421_), .B(KEYINPUT31), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n500_), .B(new_n502_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n486_), .A2(new_n487_), .A3(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n500_), .B(new_n501_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n484_), .ZN(new_n506_));
  NOR3_X1   g305(.A1(new_n466_), .A2(KEYINPUT88), .A3(new_n474_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n480_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n506_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n505_), .B1(new_n509_), .B2(new_n485_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n449_), .B1(new_n504_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n396_), .A2(KEYINPUT32), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n446_), .B(new_n513_), .C1(new_n398_), .C2(new_n445_), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n387_), .B(new_n512_), .C1(new_n398_), .C2(new_n334_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT95), .B1(new_n444_), .B2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n439_), .A2(new_n440_), .A3(new_n443_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT95), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n518_), .A2(new_n519_), .A3(new_n514_), .A4(new_n515_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n395_), .A2(KEYINPUT93), .A3(new_n399_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n423_), .A2(new_n426_), .A3(new_n430_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(new_n442_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT33), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n524_), .B1(new_n437_), .B2(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n526_), .B1(new_n525_), .B2(new_n437_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n521_), .A2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(KEYINPUT93), .B1(new_n395_), .B2(new_n399_), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n517_), .B(new_n520_), .C1(new_n528_), .C2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n503_), .B1(new_n509_), .B2(new_n485_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n511_), .A2(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(G190gat), .B(G218gat), .Z(new_n534_));
  XOR2_X1   g333(.A(G134gat), .B(G162gat), .Z(new_n535_));
  XOR2_X1   g334(.A(new_n534_), .B(new_n535_), .Z(new_n536_));
  XOR2_X1   g335(.A(new_n536_), .B(KEYINPUT36), .Z(new_n537_));
  NAND2_X1  g336(.A1(G232gat), .A2(G233gat), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n538_), .B(KEYINPUT34), .Z(new_n539_));
  XNOR2_X1  g338(.A(KEYINPUT70), .B(KEYINPUT35), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n540_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT72), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n543_), .B1(new_n305_), .B2(new_n263_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n541_), .B1(new_n544_), .B2(KEYINPUT71), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n250_), .A2(new_n313_), .A3(new_n315_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n545_), .A2(new_n547_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n537_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  XOR2_X1   g350(.A(KEYINPUT75), .B(KEYINPUT37), .Z(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n548_), .A2(new_n549_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(KEYINPUT73), .B(KEYINPUT36), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n536_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT74), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n551_), .B(new_n553_), .C1(new_n554_), .C2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n554_), .A2(new_n558_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n552_), .B1(new_n560_), .B2(new_n550_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G231gat), .A2(G233gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n257_), .B(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(new_n302_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT77), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G127gat), .B(G155gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT16), .ZN(new_n569_));
  XOR2_X1   g368(.A(G183gat), .B(G211gat), .Z(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n572_), .A2(KEYINPUT17), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n567_), .A2(new_n573_), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n565_), .A2(KEYINPUT17), .A3(new_n572_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n567_), .A2(new_n573_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n562_), .A2(new_n578_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n290_), .A2(new_n327_), .A3(new_n533_), .A4(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT96), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n444_), .A2(new_n291_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT38), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n327_), .B1(new_n284_), .B2(new_n286_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n578_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n560_), .A2(new_n550_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(KEYINPUT97), .B1(new_n533_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT97), .ZN(new_n591_));
  AOI211_X1 g390(.A(new_n591_), .B(new_n588_), .C1(new_n511_), .C2(new_n532_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n586_), .B(new_n587_), .C1(new_n590_), .C2(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(G1gat), .B1(new_n593_), .B2(new_n444_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n584_), .A2(new_n594_), .ZN(G1324gat));
  OAI21_X1  g394(.A(new_n503_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n509_), .A2(new_n505_), .A3(new_n485_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  AOI22_X1  g397(.A1(new_n598_), .A2(new_n449_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n591_), .B1(new_n599_), .B2(new_n588_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n533_), .A2(KEYINPUT97), .A3(new_n589_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n578_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT98), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n402_), .A2(new_n448_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n602_), .A2(new_n603_), .A3(new_n586_), .A4(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n605_), .A2(G8gat), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT39), .ZN(new_n607_));
  INV_X1    g406(.A(new_n604_), .ZN(new_n608_));
  OAI21_X1  g407(.A(KEYINPUT98), .B1(new_n593_), .B2(new_n608_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n606_), .A2(KEYINPUT99), .A3(new_n607_), .A4(new_n609_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n609_), .A2(new_n607_), .A3(G8gat), .A4(new_n605_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT99), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n605_), .A2(G8gat), .ZN(new_n614_));
  AOI211_X1 g413(.A(new_n585_), .B(new_n578_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n603_), .B1(new_n615_), .B2(new_n604_), .ZN(new_n616_));
  OAI21_X1  g415(.A(KEYINPUT39), .B1(new_n614_), .B2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n610_), .A2(new_n613_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(G8gat), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n581_), .A2(new_n619_), .A3(new_n604_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT40), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n618_), .A2(KEYINPUT40), .A3(new_n620_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1325gat));
  INV_X1    g424(.A(G15gat), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n581_), .A2(new_n626_), .A3(new_n503_), .ZN(new_n627_));
  OAI21_X1  g426(.A(G15gat), .B1(new_n593_), .B2(new_n505_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(KEYINPUT41), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n628_), .A2(KEYINPUT41), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n627_), .A2(new_n629_), .A3(new_n630_), .ZN(G1326gat));
  INV_X1    g430(.A(G22gat), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n486_), .A2(new_n487_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n581_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n633_), .ZN(new_n635_));
  OAI21_X1  g434(.A(G22gat), .B1(new_n593_), .B2(new_n635_), .ZN(new_n636_));
  XOR2_X1   g435(.A(KEYINPUT100), .B(KEYINPUT42), .Z(new_n637_));
  OR2_X1    g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n637_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n634_), .A2(new_n638_), .A3(new_n639_), .ZN(G1327gat));
  NAND2_X1  g439(.A1(new_n578_), .A2(new_n588_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n585_), .A2(new_n599_), .A3(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(G29gat), .B1(new_n642_), .B2(new_n518_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n562_), .ZN(new_n644_));
  OAI21_X1  g443(.A(KEYINPUT43), .B1(new_n599_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT43), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n533_), .A2(new_n646_), .A3(new_n562_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n648_), .A2(new_n586_), .A3(new_n578_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n651_), .A2(G29gat), .A3(new_n518_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n587_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n653_), .A2(KEYINPUT44), .A3(new_n586_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n643_), .B1(new_n652_), .B2(new_n654_), .ZN(G1328gat));
  INV_X1    g454(.A(KEYINPUT102), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(KEYINPUT46), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n651_), .A2(new_n604_), .A3(new_n654_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(G36gat), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(KEYINPUT101), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n658_), .A2(new_n661_), .A3(G36gat), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n656_), .A2(KEYINPUT46), .ZN(new_n664_));
  INV_X1    g463(.A(G36gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n642_), .A2(new_n665_), .A3(new_n604_), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n666_), .A2(KEYINPUT45), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(KEYINPUT45), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n664_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n657_), .B1(new_n663_), .B2(new_n669_), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n658_), .A2(new_n661_), .A3(G36gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n661_), .B1(new_n658_), .B2(G36gat), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n669_), .B(new_n657_), .C1(new_n671_), .C2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n670_), .A2(new_n674_), .ZN(G1329gat));
  NAND4_X1  g474(.A1(new_n651_), .A2(G43gat), .A3(new_n503_), .A4(new_n654_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n642_), .A2(new_n503_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n676_), .B1(G43gat), .B2(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g478(.A(G50gat), .B1(new_n642_), .B2(new_n633_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n651_), .A2(G50gat), .A3(new_n633_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n681_), .B2(new_n654_), .ZN(G1331gat));
  NOR3_X1   g481(.A1(new_n284_), .A2(new_n286_), .A3(new_n327_), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n683_), .A2(new_n533_), .A3(new_n579_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(new_n206_), .A3(new_n518_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n290_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n327_), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n686_), .A2(new_n687_), .A3(new_n602_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n688_), .A2(new_n518_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n685_), .B1(new_n689_), .B2(new_n206_), .ZN(G1332gat));
  NAND3_X1  g489(.A1(new_n684_), .A2(new_n204_), .A3(new_n604_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n688_), .ZN(new_n692_));
  OAI21_X1  g491(.A(G64gat), .B1(new_n692_), .B2(new_n608_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n693_), .A2(KEYINPUT48), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n693_), .A2(KEYINPUT48), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n691_), .B1(new_n694_), .B2(new_n695_), .ZN(G1333gat));
  INV_X1    g495(.A(G71gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n684_), .A2(new_n697_), .A3(new_n503_), .ZN(new_n698_));
  OAI21_X1  g497(.A(G71gat), .B1(new_n692_), .B2(new_n505_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n699_), .A2(KEYINPUT49), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(KEYINPUT49), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n698_), .B1(new_n700_), .B2(new_n701_), .ZN(G1334gat));
  INV_X1    g501(.A(G78gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n684_), .A2(new_n703_), .A3(new_n633_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G78gat), .B1(new_n692_), .B2(new_n635_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n705_), .A2(KEYINPUT50), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n705_), .A2(KEYINPUT50), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n704_), .B1(new_n706_), .B2(new_n707_), .ZN(G1335gat));
  AND2_X1   g507(.A1(new_n653_), .A2(new_n683_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(G85gat), .B1(new_n710_), .B2(new_n444_), .ZN(new_n711_));
  NOR4_X1   g510(.A1(new_n290_), .A2(new_n327_), .A3(new_n599_), .A4(new_n641_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n712_), .A2(new_n231_), .A3(new_n518_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1336gat));
  AOI21_X1  g513(.A(G92gat), .B1(new_n712_), .B2(new_n604_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT103), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n608_), .A2(new_n260_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT104), .Z(new_n718_));
  AOI21_X1  g517(.A(new_n716_), .B1(new_n709_), .B2(new_n718_), .ZN(G1337gat));
  OAI21_X1  g518(.A(G99gat), .B1(new_n710_), .B2(new_n505_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n712_), .A2(new_n240_), .A3(new_n503_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(KEYINPUT105), .A2(KEYINPUT51), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n720_), .A2(new_n721_), .A3(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(KEYINPUT105), .A2(KEYINPUT51), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n723_), .B(new_n724_), .ZN(G1338gat));
  NAND3_X1  g524(.A1(new_n712_), .A2(new_n222_), .A3(new_n633_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n653_), .A2(new_n633_), .A3(new_n683_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT52), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n727_), .A2(new_n728_), .A3(G106gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n727_), .B2(G106gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n726_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT107), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n733_), .B(new_n726_), .C1(new_n729_), .C2(new_n730_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(KEYINPUT106), .B(KEYINPUT53), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n732_), .A2(new_n734_), .A3(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n732_), .B2(new_n734_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n736_), .A2(new_n737_), .ZN(G1339gat));
  NOR2_X1   g537(.A1(new_n604_), .A2(new_n444_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n510_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n740_), .A2(KEYINPUT59), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n562_), .A2(new_n578_), .A3(new_n327_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n742_), .B1(new_n284_), .B2(new_n286_), .ZN(new_n743_));
  XOR2_X1   g542(.A(KEYINPUT108), .B(KEYINPUT54), .Z(new_n744_));
  XOR2_X1   g543(.A(new_n743_), .B(new_n744_), .Z(new_n745_));
  NAND2_X1  g544(.A1(new_n309_), .A2(new_n310_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT112), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n746_), .A2(new_n747_), .A3(new_n321_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n324_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n749_));
  OAI21_X1  g548(.A(KEYINPUT112), .B1(new_n749_), .B2(new_n323_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n316_), .A2(new_n324_), .A3(new_n306_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n748_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT113), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT113), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n748_), .A2(new_n750_), .A3(new_n754_), .A4(new_n751_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n755_), .A2(new_n326_), .ZN(new_n756_));
  AND4_X1   g555(.A1(KEYINPUT114), .A2(new_n282_), .A3(new_n753_), .A4(new_n756_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n753_), .A2(new_n326_), .A3(new_n755_), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT114), .B1(new_n758_), .B2(new_n282_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n757_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n327_), .A2(new_n281_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT109), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT110), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n266_), .B1(new_n219_), .B2(new_n250_), .ZN(new_n764_));
  OAI21_X1  g563(.A(KEYINPUT12), .B1(new_n257_), .B2(new_n263_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n219_), .A2(new_n271_), .A3(new_n250_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n764_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n763_), .B1(new_n767_), .B2(KEYINPUT55), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n273_), .A2(KEYINPUT110), .A3(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n251_), .B(new_n264_), .C1(new_n270_), .C2(new_n272_), .ZN(new_n772_));
  AOI22_X1  g571(.A1(new_n267_), .A2(new_n772_), .B1(new_n767_), .B2(KEYINPUT55), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n280_), .B1(new_n771_), .B2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(KEYINPUT111), .B1(new_n774_), .B2(KEYINPUT56), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT56), .ZN(new_n776_));
  AOI211_X1 g575(.A(new_n776_), .B(new_n280_), .C1(new_n771_), .C2(new_n773_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n762_), .B1(new_n775_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT111), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n774_), .A2(new_n779_), .A3(KEYINPUT56), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n760_), .B1(new_n778_), .B2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n782_), .A2(KEYINPUT57), .A3(new_n589_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT115), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT110), .B1(new_n273_), .B2(new_n769_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n765_), .A2(new_n766_), .ZN(new_n787_));
  AOI211_X1 g586(.A(new_n763_), .B(KEYINPUT55), .C1(new_n787_), .C2(new_n269_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n773_), .B1(new_n786_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n278_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n776_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n774_), .A2(KEYINPUT56), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(KEYINPUT111), .A3(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n793_), .A2(new_n780_), .A3(new_n762_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n588_), .B1(new_n794_), .B2(new_n760_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n795_), .A2(KEYINPUT115), .A3(KEYINPUT57), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n785_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n782_), .A2(new_n589_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT57), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n758_), .A2(new_n281_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n774_), .A2(KEYINPUT56), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n800_), .B(KEYINPUT58), .C1(new_n777_), .C2(new_n801_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n802_), .A2(new_n562_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n800_), .B1(new_n801_), .B2(new_n777_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT58), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n798_), .A2(new_n799_), .B1(new_n803_), .B2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n587_), .B1(new_n797_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n745_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT115), .B1(new_n795_), .B2(KEYINPUT57), .ZN(new_n811_));
  AND4_X1   g610(.A1(KEYINPUT115), .A2(new_n782_), .A3(KEYINPUT57), .A4(new_n589_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n807_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n813_), .A2(new_n809_), .A3(new_n578_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n741_), .B1(new_n810_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n740_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n743_), .B(new_n744_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n808_), .B2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT59), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n816_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(G113gat), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n821_), .A2(new_n822_), .A3(new_n687_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n819_), .B2(new_n687_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n824_), .A2(KEYINPUT116), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n824_), .A2(KEYINPUT116), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n823_), .A2(new_n825_), .A3(new_n826_), .ZN(G1340gat));
  XNOR2_X1  g626(.A(KEYINPUT118), .B(G120gat), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n806_), .A2(new_n562_), .A3(new_n802_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n795_), .B2(KEYINPUT57), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n830_), .B1(new_n785_), .B2(new_n796_), .ZN(new_n831_));
  OAI21_X1  g630(.A(KEYINPUT117), .B1(new_n831_), .B2(new_n587_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(new_n745_), .A3(new_n814_), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n833_), .A2(new_n741_), .B1(KEYINPUT59), .B2(new_n819_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n828_), .B1(new_n834_), .B2(new_n686_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n819_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT60), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n287_), .A2(new_n837_), .A3(new_n828_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n837_), .B2(new_n828_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n836_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT119), .B1(new_n835_), .B2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n816_), .A2(new_n686_), .A3(new_n820_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n828_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n846_), .A3(new_n840_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n842_), .A2(new_n847_), .ZN(G1341gat));
  OAI21_X1  g647(.A(G127gat), .B1(new_n821_), .B2(new_n578_), .ZN(new_n849_));
  OR2_X1    g648(.A1(new_n578_), .A2(G127gat), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n819_), .B2(new_n850_), .ZN(G1342gat));
  AOI21_X1  g650(.A(G134gat), .B1(new_n836_), .B2(new_n588_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n562_), .A2(G134gat), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(KEYINPUT120), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n852_), .B1(new_n834_), .B2(new_n854_), .ZN(G1343gat));
  OAI211_X1 g654(.A(new_n504_), .B(new_n739_), .C1(new_n808_), .C2(new_n818_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(new_n687_), .ZN(new_n857_));
  XOR2_X1   g656(.A(new_n857_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g657(.A1(new_n856_), .A2(new_n290_), .ZN(new_n859_));
  XOR2_X1   g658(.A(new_n859_), .B(G148gat), .Z(G1345gat));
  OR3_X1    g659(.A1(new_n856_), .A2(KEYINPUT121), .A3(new_n578_), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT121), .B1(new_n856_), .B2(new_n578_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  XOR2_X1   g662(.A(KEYINPUT61), .B(G155gat), .Z(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(KEYINPUT122), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n863_), .B(new_n866_), .ZN(G1346gat));
  INV_X1    g666(.A(G162gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n868_), .B1(new_n856_), .B2(new_n589_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(KEYINPUT123), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n808_), .A2(new_n818_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(new_n597_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n872_), .A2(G162gat), .A3(new_n562_), .A4(new_n739_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT123), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n874_), .B(new_n868_), .C1(new_n856_), .C2(new_n589_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n870_), .A2(new_n873_), .A3(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT124), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT124), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n870_), .A2(new_n873_), .A3(new_n878_), .A4(new_n875_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n879_), .ZN(G1347gat));
  NOR2_X1   g679(.A1(new_n608_), .A2(new_n518_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n510_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n833_), .A2(new_n883_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n884_), .A2(new_n327_), .A3(new_n348_), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n327_), .B(new_n883_), .C1(new_n810_), .C2(new_n815_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n886_), .A2(new_n887_), .A3(G169gat), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n886_), .B2(G169gat), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT125), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n888_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  AOI211_X1 g690(.A(KEYINPUT125), .B(new_n887_), .C1(new_n886_), .C2(G169gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n885_), .B1(new_n891_), .B2(new_n892_), .ZN(G1348gat));
  AOI21_X1  g692(.A(G176gat), .B1(new_n884_), .B2(new_n287_), .ZN(new_n894_));
  NOR4_X1   g693(.A1(new_n871_), .A2(new_n349_), .A3(new_n290_), .A4(new_n882_), .ZN(new_n895_));
  OR2_X1    g694(.A1(new_n895_), .A2(KEYINPUT126), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(KEYINPUT126), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n894_), .B1(new_n896_), .B2(new_n897_), .ZN(G1349gat));
  NOR2_X1   g697(.A1(new_n578_), .A2(new_n370_), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n587_), .B(new_n883_), .C1(new_n808_), .C2(new_n818_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n378_), .ZN(new_n901_));
  AOI22_X1  g700(.A1(new_n884_), .A2(new_n899_), .B1(new_n900_), .B2(new_n901_), .ZN(G1350gat));
  NAND2_X1  g701(.A1(new_n884_), .A2(new_n562_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(G190gat), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n884_), .A2(new_n588_), .A3(new_n369_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1351gat));
  NAND2_X1  g705(.A1(new_n872_), .A2(new_n881_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n687_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT127), .B(G197gat), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(G1352gat));
  NAND3_X1  g709(.A1(new_n872_), .A2(new_n686_), .A3(new_n881_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g711(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n587_), .A2(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n907_), .A2(new_n914_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n915_), .B(new_n916_), .ZN(G1354gat));
  OAI21_X1  g716(.A(G218gat), .B1(new_n907_), .B2(new_n644_), .ZN(new_n918_));
  OR2_X1    g717(.A1(new_n589_), .A2(G218gat), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n907_), .B2(new_n919_), .ZN(G1355gat));
endmodule


