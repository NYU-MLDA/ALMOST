//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n866_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  XOR2_X1   g001(.A(G85gat), .B(G92gat), .Z(new_n203_));
  NAND2_X1  g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT6), .ZN(new_n205_));
  OR2_X1    g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n205_), .B1(KEYINPUT7), .B2(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n203_), .B1(new_n207_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(KEYINPUT10), .B(G99gat), .Z(new_n214_));
  INV_X1    g013(.A(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n203_), .A2(KEYINPUT9), .ZN(new_n217_));
  INV_X1    g016(.A(G85gat), .ZN(new_n218_));
  INV_X1    g017(.A(G92gat), .ZN(new_n219_));
  OR3_X1    g018(.A1(new_n218_), .A2(new_n219_), .A3(KEYINPUT9), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n216_), .A2(new_n217_), .A3(new_n220_), .A4(new_n205_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n213_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G57gat), .B(G64gat), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n224_), .A2(KEYINPUT11), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(KEYINPUT11), .ZN(new_n226_));
  XOR2_X1   g025(.A(G71gat), .B(G78gat), .Z(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n226_), .A2(new_n227_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n223_), .A2(new_n230_), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n229_), .B(new_n228_), .C1(new_n213_), .C2(new_n222_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT12), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n231_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n232_), .A2(new_n233_), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n235_), .A2(KEYINPUT66), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(KEYINPUT66), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n234_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G230gat), .A2(G233gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n231_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n232_), .ZN(new_n242_));
  OAI211_X1 g041(.A(G230gat), .B(G233gat), .C1(new_n241_), .C2(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G120gat), .B(G148gat), .Z(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G176gat), .B(G204gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n240_), .A2(new_n243_), .A3(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n248_), .B(KEYINPUT68), .Z(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n251_), .B1(new_n240_), .B2(new_n243_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n202_), .B1(new_n249_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n240_), .A2(new_n243_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(new_n250_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n240_), .A2(new_n243_), .A3(new_n248_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(KEYINPUT13), .A3(new_n256_), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n253_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G231gat), .A2(G233gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n230_), .B(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G1gat), .B(G8gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT73), .ZN(new_n262_));
  OR2_X1    g061(.A1(G15gat), .A2(G22gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G15gat), .A2(G22gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G1gat), .A2(G8gat), .ZN(new_n265_));
  AOI22_X1  g064(.A1(new_n263_), .A2(new_n264_), .B1(KEYINPUT14), .B2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n262_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n260_), .B(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT17), .ZN(new_n270_));
  XOR2_X1   g069(.A(G127gat), .B(G155gat), .Z(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT16), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G183gat), .B(G211gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  OR3_X1    g073(.A1(new_n269_), .A2(new_n270_), .A3(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(KEYINPUT17), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n269_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT37), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G232gat), .A2(G233gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT34), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n281_), .B1(new_n283_), .B2(KEYINPUT35), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G29gat), .B(G36gat), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n285_), .A2(KEYINPUT69), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n285_), .A2(KEYINPUT69), .ZN(new_n287_));
  XOR2_X1   g086(.A(G43gat), .B(G50gat), .Z(new_n288_));
  OR3_X1    g087(.A1(new_n286_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n288_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT15), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n212_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n211_), .B(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(new_n221_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n284_), .B1(new_n293_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n291_), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT70), .B1(new_n223_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT70), .ZN(new_n300_));
  NOR4_X1   g099(.A1(new_n213_), .A2(new_n300_), .A3(new_n291_), .A4(new_n222_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n297_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n283_), .A2(KEYINPUT35), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n303_), .B(new_n297_), .C1(new_n299_), .C2(new_n301_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G190gat), .B(G218gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G134gat), .B(G162gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n311_), .A2(KEYINPUT36), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n308_), .A2(new_n313_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .A4(new_n312_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n311_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT36), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n320_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n280_), .B1(new_n316_), .B2(new_n322_), .ZN(new_n323_));
  AOI211_X1 g122(.A(KEYINPUT37), .B(new_n321_), .C1(new_n314_), .C2(new_n315_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n258_), .A2(new_n279_), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n298_), .A2(new_n267_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT74), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G229gat), .A2(G233gat), .ZN(new_n331_));
  INV_X1    g130(.A(new_n267_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n293_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n330_), .A2(new_n331_), .A3(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n291_), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n330_), .A2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n334_), .B1(new_n336_), .B2(new_n331_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G113gat), .B(G141gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT75), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G169gat), .B(G197gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT76), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n337_), .A2(KEYINPUT77), .A3(new_n342_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n334_), .B(new_n341_), .C1(new_n336_), .C2(new_n331_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(KEYINPUT77), .B1(new_n337_), .B2(new_n342_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT78), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n337_), .A2(new_n342_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT78), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n350_), .A2(new_n351_), .A3(new_n344_), .A4(new_n343_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n347_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT25), .B(G183gat), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT26), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(G190gat), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT26), .B(G190gat), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n355_), .B(new_n359_), .C1(new_n360_), .C2(new_n358_), .ZN(new_n361_));
  NOR3_X1   g160(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G169gat), .A2(G176gat), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n362_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G183gat), .A2(G190gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT23), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT80), .B(KEYINPUT23), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n370_), .B1(new_n371_), .B2(new_n368_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n361_), .A2(new_n366_), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(G183gat), .ZN(new_n374_));
  INV_X1    g173(.A(G190gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n367_), .A2(new_n369_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n376_), .B(new_n377_), .C1(new_n371_), .C2(new_n367_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(G169gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n373_), .A2(new_n381_), .ZN(new_n382_));
  AND2_X1   g181(.A1(G197gat), .A2(G204gat), .ZN(new_n383_));
  NOR2_X1   g182(.A1(G197gat), .A2(G204gat), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT85), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G211gat), .B(G218gat), .ZN(new_n386_));
  AOI21_X1  g185(.A(KEYINPUT21), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n386_), .ZN(new_n388_));
  INV_X1    g187(.A(G218gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(G211gat), .ZN(new_n390_));
  INV_X1    g189(.A(G211gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(G218gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(G197gat), .ZN(new_n394_));
  INV_X1    g193(.A(G204gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G197gat), .A2(G204gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n393_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n388_), .A2(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n387_), .B1(new_n400_), .B2(KEYINPUT21), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n382_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT90), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT90), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n382_), .A2(new_n401_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G226gat), .A2(G233gat), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n407_), .B(KEYINPUT19), .Z(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT20), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT80), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n410_), .A2(KEYINPUT23), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n369_), .A2(KEYINPUT80), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n368_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n375_), .A2(KEYINPUT26), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n374_), .A2(KEYINPUT25), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT25), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(G183gat), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n357_), .A2(new_n414_), .A3(new_n415_), .A4(new_n417_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n413_), .A2(new_n418_), .A3(new_n377_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n369_), .A2(KEYINPUT80), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n410_), .A2(KEYINPUT23), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n368_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n367_), .A2(KEYINPUT23), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n376_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n419_), .A2(new_n366_), .B1(new_n424_), .B2(new_n380_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT85), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n426_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n427_), .A2(new_n393_), .ZN(new_n428_));
  AOI22_X1  g227(.A1(new_n390_), .A2(new_n392_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT21), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n387_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n409_), .B1(new_n425_), .B2(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT91), .B1(new_n406_), .B2(new_n433_), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n382_), .A2(new_n401_), .A3(new_n404_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n404_), .B1(new_n382_), .B2(new_n401_), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n433_), .B(KEYINPUT91), .C1(new_n435_), .C2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT20), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n366_), .A2(new_n413_), .A3(new_n377_), .A4(new_n418_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n367_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n441_));
  AOI22_X1  g240(.A1(new_n441_), .A2(new_n370_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n380_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n440_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n439_), .B1(new_n444_), .B2(new_n401_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT21), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n446_), .B1(new_n388_), .B2(new_n399_), .ZN(new_n447_));
  OAI211_X1 g246(.A(new_n373_), .B(new_n381_), .C1(new_n447_), .C2(new_n387_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n445_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n408_), .ZN(new_n450_));
  AOI21_X1  g249(.A(KEYINPUT89), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT89), .ZN(new_n452_));
  AOI211_X1 g251(.A(new_n452_), .B(new_n408_), .C1(new_n445_), .C2(new_n448_), .ZN(new_n453_));
  OAI22_X1  g252(.A1(new_n434_), .A2(new_n438_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n454_));
  XOR2_X1   g253(.A(G8gat), .B(G36gat), .Z(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G64gat), .B(G92gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n454_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n449_), .A2(new_n450_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n452_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n449_), .A2(KEYINPUT89), .A3(new_n450_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n433_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT91), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(new_n437_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n459_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n464_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n460_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT27), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n449_), .A2(new_n450_), .ZN(new_n474_));
  XOR2_X1   g273(.A(KEYINPUT97), .B(KEYINPUT20), .Z(new_n475_));
  OAI21_X1  g274(.A(new_n475_), .B1(new_n444_), .B2(new_n401_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT98), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  OAI211_X1 g277(.A(KEYINPUT98), .B(new_n475_), .C1(new_n444_), .C2(new_n401_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n406_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n474_), .B1(new_n480_), .B2(new_n450_), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT100), .B1(new_n481_), .B2(new_n469_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n479_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n476_), .A2(new_n477_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n450_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n474_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT100), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(new_n488_), .A3(new_n459_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n482_), .A2(new_n489_), .A3(KEYINPUT27), .A4(new_n470_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n473_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(G233gat), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n492_), .A2(KEYINPUT84), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(KEYINPUT84), .ZN(new_n494_));
  OAI21_X1  g293(.A(G228gat), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT29), .ZN(new_n496_));
  NOR2_X1   g295(.A1(G141gat), .A2(G148gat), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT3), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G141gat), .A2(G148gat), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT2), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n499_), .A2(new_n502_), .A3(new_n503_), .A4(new_n504_), .ZN(new_n505_));
  OR2_X1    g304(.A1(G155gat), .A2(G162gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G155gat), .A2(G162gat), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(KEYINPUT1), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT1), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n510_), .A2(G155gat), .A3(G162gat), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n509_), .A2(new_n511_), .A3(new_n506_), .ZN(new_n512_));
  XOR2_X1   g311(.A(G141gat), .B(G148gat), .Z(new_n513_));
  AOI22_X1  g312(.A1(new_n505_), .A2(new_n508_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n401_), .B(new_n495_), .C1(new_n496_), .C2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G78gat), .B(G106gat), .ZN(new_n516_));
  XOR2_X1   g315(.A(KEYINPUT86), .B(KEYINPUT29), .Z(new_n517_));
  OR2_X1    g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n495_), .B1(new_n518_), .B2(new_n401_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT87), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  AOI211_X1 g320(.A(KEYINPUT87), .B(new_n495_), .C1(new_n518_), .C2(new_n401_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n515_), .B(new_n516_), .C1(new_n521_), .C2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT83), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n514_), .A2(new_n517_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n432_), .A2(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(KEYINPUT87), .B1(new_n527_), .B2(new_n495_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n519_), .A2(new_n520_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n516_), .B1(new_n530_), .B2(new_n515_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G22gat), .B(G50gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n505_), .A2(new_n508_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n512_), .A2(new_n513_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT28), .B1(new_n535_), .B2(KEYINPUT29), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT28), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n514_), .A2(new_n537_), .A3(new_n496_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT88), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT88), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n536_), .A2(new_n541_), .A3(new_n538_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n532_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n540_), .A2(new_n532_), .A3(new_n542_), .ZN(new_n544_));
  OAI22_X1  g343(.A1(new_n525_), .A2(new_n531_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n515_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n516_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n544_), .A2(new_n543_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n548_), .A2(new_n549_), .A3(new_n524_), .A4(new_n523_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n545_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G71gat), .B(G99gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(G43gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n382_), .B(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G113gat), .B(G120gat), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT82), .ZN(new_n556_));
  INV_X1    g355(.A(G120gat), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(G113gat), .ZN(new_n558_));
  INV_X1    g357(.A(G113gat), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(G120gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT82), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(G127gat), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n564_), .A2(G134gat), .ZN(new_n565_));
  INV_X1    g364(.A(G134gat), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n566_), .A2(G127gat), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT81), .B1(new_n565_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(G127gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n564_), .A2(G134gat), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT81), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n569_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  AND4_X1   g371(.A1(new_n556_), .A2(new_n563_), .A3(new_n568_), .A4(new_n572_), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n556_), .A2(new_n563_), .B1(new_n568_), .B2(new_n572_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n554_), .B(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G227gat), .A2(G233gat), .ZN(new_n577_));
  INV_X1    g376(.A(G15gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT30), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT31), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n576_), .B(new_n581_), .Z(new_n582_));
  OAI21_X1  g381(.A(new_n514_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n555_), .A2(KEYINPUT82), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n558_), .A2(new_n560_), .A3(KEYINPUT82), .ZN(new_n585_));
  INV_X1    g384(.A(new_n572_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n571_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n587_));
  OAI22_X1  g386(.A1(new_n584_), .A2(new_n585_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n563_), .A2(new_n556_), .A3(new_n568_), .A4(new_n572_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n535_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G225gat), .A2(G233gat), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n583_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT4), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n535_), .A2(new_n588_), .A3(new_n589_), .A4(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT94), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n583_), .A2(KEYINPUT4), .A3(new_n590_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n591_), .B(KEYINPUT93), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n592_), .B1(new_n595_), .B2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G1gat), .B(G29gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G57gat), .B(G85gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n599_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT99), .ZN(new_n606_));
  INV_X1    g405(.A(new_n604_), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n592_), .B(new_n607_), .C1(new_n595_), .C2(new_n598_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n605_), .A2(new_n606_), .A3(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n599_), .A2(KEYINPUT99), .A3(new_n604_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n582_), .A2(new_n611_), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n491_), .A2(new_n551_), .A3(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n469_), .A2(KEYINPUT32), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n487_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n464_), .A2(new_n468_), .A3(new_n614_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n609_), .A2(new_n616_), .A3(new_n617_), .A4(new_n610_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n608_), .A2(KEYINPUT96), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT33), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n596_), .A2(new_n591_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n595_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n583_), .A2(new_n590_), .A3(new_n597_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n623_), .A2(new_n604_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n608_), .A2(KEYINPUT96), .A3(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n620_), .A2(new_n625_), .A3(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n618_), .B1(new_n628_), .B2(new_n471_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n551_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  AOI22_X1  g430(.A1(new_n545_), .A2(new_n550_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n473_), .A2(new_n632_), .A3(new_n490_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n582_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n613_), .B1(new_n634_), .B2(KEYINPUT101), .ZN(new_n635_));
  INV_X1    g434(.A(new_n582_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n473_), .A2(new_n632_), .A3(new_n490_), .ZN(new_n637_));
  AOI22_X1  g436(.A1(new_n619_), .A2(KEYINPUT33), .B1(new_n622_), .B2(new_n624_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n638_), .A2(new_n470_), .A3(new_n460_), .A4(new_n627_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n551_), .B1(new_n639_), .B2(new_n618_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n636_), .B1(new_n637_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT101), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n354_), .B1(new_n635_), .B2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n327_), .A2(new_n644_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n645_), .A2(G1gat), .A3(new_n611_), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n646_), .A2(KEYINPUT38), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n258_), .A2(new_n353_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT102), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n258_), .A2(KEYINPUT102), .A3(new_n353_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n650_), .A2(new_n279_), .A3(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n321_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n654_), .B1(new_n635_), .B2(new_n643_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n652_), .A2(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G1gat), .B1(new_n656_), .B2(new_n611_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n646_), .A2(KEYINPUT38), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n647_), .A2(new_n657_), .A3(new_n658_), .ZN(G1324gat));
  INV_X1    g458(.A(new_n491_), .ZN(new_n660_));
  OR3_X1    g459(.A1(new_n645_), .A2(G8gat), .A3(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G8gat), .B1(new_n656_), .B2(new_n660_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n662_), .A2(KEYINPUT39), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(KEYINPUT39), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n661_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n665_), .B(new_n666_), .Z(G1325gat));
  OAI21_X1  g466(.A(G15gat), .B1(new_n656_), .B2(new_n636_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT41), .Z(new_n669_));
  NAND2_X1  g468(.A1(new_n582_), .A2(new_n578_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n669_), .B1(new_n645_), .B2(new_n670_), .ZN(G1326gat));
  OAI21_X1  g470(.A(G22gat), .B1(new_n656_), .B2(new_n630_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT42), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n630_), .A2(G22gat), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n673_), .B1(new_n645_), .B2(new_n674_), .ZN(G1327gat));
  NAND3_X1  g474(.A1(new_n650_), .A2(new_n278_), .A3(new_n651_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT104), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n325_), .B1(new_n635_), .B2(new_n643_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n678_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n653_), .B(new_n280_), .ZN(new_n682_));
  OAI211_X1 g481(.A(KEYINPUT101), .B(new_n636_), .C1(new_n637_), .C2(new_n640_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n613_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n634_), .A2(KEYINPUT101), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n682_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n687_), .A2(KEYINPUT105), .A3(KEYINPUT43), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n681_), .A2(new_n688_), .ZN(new_n689_));
  OAI211_X1 g488(.A(new_n680_), .B(new_n682_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT106), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n635_), .A2(new_n643_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n692_), .A2(new_n693_), .A3(new_n680_), .A4(new_n682_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n691_), .A2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n689_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n677_), .A2(new_n696_), .ZN(new_n697_));
  XOR2_X1   g496(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n611_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n677_), .A2(KEYINPUT44), .A3(new_n696_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n700_), .A2(G29gat), .A3(new_n701_), .A4(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(G29gat), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n653_), .A2(new_n279_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n258_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(new_n644_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n704_), .B1(new_n707_), .B2(new_n611_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n703_), .A2(new_n708_), .ZN(G1328gat));
  NOR3_X1   g508(.A1(new_n707_), .A2(G36gat), .A3(new_n660_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT45), .Z(new_n711_));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n711_), .B1(new_n712_), .B2(KEYINPUT46), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n700_), .A2(new_n491_), .A3(new_n702_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n714_), .B2(G36gat), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT46), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n716_), .A2(KEYINPUT108), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n715_), .B(new_n717_), .ZN(G1329gat));
  NAND2_X1  g517(.A1(new_n700_), .A2(new_n702_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n582_), .A2(G43gat), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n707_), .A2(new_n636_), .ZN(new_n721_));
  OAI22_X1  g520(.A1(new_n719_), .A2(new_n720_), .B1(G43gat), .B2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g522(.A(G50gat), .B1(new_n719_), .B2(new_n630_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n630_), .A2(G50gat), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT109), .Z(new_n726_));
  OAI21_X1  g525(.A(new_n724_), .B1(new_n707_), .B2(new_n726_), .ZN(G1331gat));
  INV_X1    g526(.A(new_n258_), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n655_), .A2(new_n354_), .A3(new_n728_), .A4(new_n279_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G57gat), .B1(new_n729_), .B2(new_n611_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n692_), .A2(KEYINPUT110), .A3(new_n354_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(KEYINPUT110), .B1(new_n692_), .B2(new_n354_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n732_), .A2(new_n258_), .A3(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(new_n279_), .A3(new_n325_), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n611_), .A2(G57gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n730_), .B1(new_n735_), .B2(new_n736_), .ZN(G1332gat));
  OAI21_X1  g536(.A(G64gat), .B1(new_n729_), .B2(new_n660_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT48), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n660_), .A2(G64gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n735_), .B2(new_n740_), .ZN(G1333gat));
  OAI21_X1  g540(.A(G71gat), .B1(new_n729_), .B2(new_n636_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT49), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n636_), .A2(G71gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n735_), .B2(new_n744_), .ZN(G1334gat));
  OAI21_X1  g544(.A(G78gat), .B1(new_n729_), .B2(new_n630_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT50), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n630_), .A2(G78gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n735_), .B2(new_n748_), .ZN(G1335gat));
  NAND2_X1  g548(.A1(new_n734_), .A2(new_n705_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n751_), .A2(new_n218_), .A3(new_n701_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n258_), .A2(new_n353_), .A3(new_n279_), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n689_), .A2(KEYINPUT111), .A3(new_n695_), .ZN(new_n754_));
  AOI21_X1  g553(.A(KEYINPUT111), .B1(new_n689_), .B2(new_n695_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n753_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  OAI211_X1 g557(.A(KEYINPUT112), .B(new_n753_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n758_), .A2(new_n701_), .A3(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n752_), .B1(new_n760_), .B2(new_n218_), .ZN(G1336gat));
  NAND3_X1  g560(.A1(new_n751_), .A2(new_n219_), .A3(new_n491_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n758_), .A2(new_n491_), .A3(new_n759_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(new_n219_), .ZN(G1337gat));
  NAND3_X1  g563(.A1(new_n758_), .A2(new_n582_), .A3(new_n759_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(G99gat), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n582_), .A2(new_n214_), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT113), .B1(new_n751_), .B2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n766_), .A2(new_n768_), .A3(new_n770_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(G1338gat));
  AND2_X1   g573(.A1(new_n753_), .A2(new_n551_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n215_), .B1(new_n696_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT117), .ZN(new_n777_));
  XOR2_X1   g576(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n778_));
  OR3_X1    g577(.A1(new_n776_), .A2(new_n777_), .A3(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n776_), .A2(new_n778_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT116), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n777_), .B1(new_n776_), .B2(new_n778_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n776_), .A2(KEYINPUT116), .A3(new_n778_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n779_), .A2(new_n782_), .A3(new_n783_), .A4(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n751_), .A2(new_n215_), .A3(new_n551_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n785_), .A2(new_n786_), .A3(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(G1339gat));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n791_), .B1(new_n327_), .B2(new_n354_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n326_), .A2(KEYINPUT54), .A3(new_n353_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n353_), .A2(new_n256_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT55), .B1(new_n238_), .B2(new_n239_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n240_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n238_), .A2(KEYINPUT55), .A3(new_n239_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT56), .B1(new_n799_), .B2(new_n250_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT56), .ZN(new_n802_));
  AOI211_X1 g601(.A(new_n802_), .B(new_n251_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n795_), .B1(new_n801_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n336_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n341_), .B1(new_n806_), .B2(new_n331_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n330_), .A2(new_n333_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n809_));
  OAI211_X1 g608(.A(G229gat), .B(G233gat), .C1(new_n808_), .C2(new_n809_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n808_), .A2(new_n809_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n807_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n344_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n653_), .B1(new_n805_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  OAI211_X1 g616(.A(KEYINPUT57), .B(new_n653_), .C1(new_n805_), .C2(new_n814_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n813_), .A2(new_n249_), .ZN(new_n819_));
  OAI211_X1 g618(.A(KEYINPUT58), .B(new_n819_), .C1(new_n800_), .C2(new_n803_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n820_), .A2(new_n682_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n819_), .B1(new_n800_), .B2(new_n803_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT58), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n821_), .A2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n817_), .A2(new_n818_), .A3(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n794_), .B1(new_n826_), .B2(new_n278_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n491_), .A2(new_n551_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n828_), .A2(new_n582_), .A3(new_n701_), .ZN(new_n829_));
  OAI21_X1  g628(.A(KEYINPUT120), .B1(new_n827_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT120), .ZN(new_n831_));
  INV_X1    g630(.A(new_n829_), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n815_), .A2(new_n816_), .B1(new_n821_), .B2(new_n824_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n279_), .B1(new_n833_), .B2(new_n818_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n831_), .B(new_n832_), .C1(new_n834_), .C2(new_n794_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n830_), .A2(new_n835_), .A3(new_n559_), .A4(new_n353_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT59), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(new_n827_), .B2(new_n829_), .ZN(new_n838_));
  OAI211_X1 g637(.A(KEYINPUT59), .B(new_n832_), .C1(new_n834_), .C2(new_n794_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n354_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n836_), .B1(new_n840_), .B2(new_n559_), .ZN(G1340gat));
  OAI21_X1  g640(.A(new_n557_), .B1(new_n258_), .B2(KEYINPUT60), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n557_), .A2(KEYINPUT60), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(KEYINPUT121), .B2(new_n843_), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n842_), .A2(KEYINPUT121), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n830_), .A2(new_n835_), .A3(new_n844_), .A4(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n258_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n847_), .B2(new_n557_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT122), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  OAI211_X1 g649(.A(KEYINPUT122), .B(new_n846_), .C1(new_n847_), .C2(new_n557_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1341gat));
  NAND3_X1  g651(.A1(new_n830_), .A2(new_n835_), .A3(new_n279_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n838_), .A2(new_n839_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n279_), .A2(G127gat), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT123), .ZN(new_n856_));
  AOI22_X1  g655(.A1(new_n853_), .A2(new_n564_), .B1(new_n854_), .B2(new_n856_), .ZN(G1342gat));
  NAND4_X1  g656(.A1(new_n830_), .A2(new_n835_), .A3(new_n566_), .A4(new_n654_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n325_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n859_), .B2(new_n566_), .ZN(G1343gat));
  NAND3_X1  g659(.A1(new_n636_), .A2(new_n551_), .A3(new_n701_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n827_), .A2(new_n491_), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n353_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n728_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(KEYINPUT124), .B(G148gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1345gat));
  NAND2_X1  g666(.A1(new_n862_), .A2(new_n279_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(KEYINPUT61), .B(G155gat), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n868_), .B(new_n869_), .ZN(G1346gat));
  AOI21_X1  g669(.A(G162gat), .B1(new_n862_), .B2(new_n654_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n682_), .A2(G162gat), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(KEYINPUT125), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n871_), .B1(new_n862_), .B2(new_n873_), .ZN(G1347gat));
  NOR2_X1   g673(.A1(new_n827_), .A2(new_n551_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n660_), .A2(new_n612_), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(KEYINPUT22), .B(G169gat), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n877_), .A2(new_n353_), .A3(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(G169gat), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n353_), .A2(new_n876_), .ZN(new_n881_));
  XOR2_X1   g680(.A(new_n881_), .B(KEYINPUT126), .Z(new_n882_));
  AOI21_X1  g681(.A(new_n880_), .B1(new_n875_), .B2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n883_), .A2(new_n884_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n879_), .B1(new_n885_), .B2(new_n886_), .ZN(G1348gat));
  NAND2_X1  g686(.A1(new_n877_), .A2(new_n728_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g688(.A1(new_n875_), .A2(new_n279_), .A3(new_n876_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n355_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n891_), .B1(new_n374_), .B2(new_n890_), .ZN(G1350gat));
  NAND3_X1  g691(.A1(new_n877_), .A2(new_n360_), .A3(new_n654_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n877_), .A2(new_n682_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(new_n375_), .ZN(G1351gat));
  INV_X1    g694(.A(new_n827_), .ZN(new_n896_));
  AND3_X1   g695(.A1(new_n491_), .A2(new_n636_), .A3(new_n632_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n354_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n394_), .ZN(G1352gat));
  NOR2_X1   g699(.A1(new_n898_), .A2(new_n258_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(new_n395_), .ZN(G1353gat));
  NOR2_X1   g701(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n903_));
  AND2_X1   g702(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n904_));
  NOR4_X1   g703(.A1(new_n898_), .A2(new_n278_), .A3(new_n903_), .A4(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n898_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n279_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n905_), .B1(new_n907_), .B2(new_n903_), .ZN(G1354gat));
  AOI21_X1  g707(.A(G218gat), .B1(new_n906_), .B2(new_n654_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n325_), .A2(new_n389_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(KEYINPUT127), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n909_), .B1(new_n906_), .B2(new_n911_), .ZN(G1355gat));
endmodule


