//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 0 1 0 0 0 1 1 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n778_,
    new_n779_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n816_, new_n817_, new_n818_, new_n820_, new_n821_,
    new_n822_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n924_,
    new_n926_, new_n927_, new_n928_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_, new_n951_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n958_, new_n959_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n986_, new_n987_, new_n988_,
    new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_,
    new_n995_, new_n996_, new_n997_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT78), .ZN(new_n203_));
  XOR2_X1   g002(.A(G71gat), .B(G99gat), .Z(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT25), .B(G183gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT26), .B(G190gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT74), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT74), .A2(G169gat), .A3(G176gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n211_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n209_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT75), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT75), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n209_), .A2(new_n216_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT23), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT23), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(G183gat), .A3(G190gat), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  NOR3_X1   g024(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n218_), .A2(new_n220_), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(G169gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT22), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT22), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(G169gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n233_), .A2(G176gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n214_), .A2(new_n215_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT76), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n235_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT76), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n237_), .B(new_n238_), .C1(G176gat), .C2(new_n233_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n224_), .A2(KEYINPUT77), .ZN(new_n240_));
  INV_X1    g039(.A(G183gat), .ZN(new_n241_));
  INV_X1    g040(.A(G190gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n222_), .A2(new_n224_), .A3(KEYINPUT77), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n240_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n236_), .A2(new_n239_), .A3(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n228_), .A2(KEYINPUT30), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT30), .B1(new_n228_), .B2(new_n246_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n206_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n249_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n251_), .A2(new_n247_), .A3(new_n205_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G15gat), .B(G43gat), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT79), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n250_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT31), .ZN(new_n260_));
  INV_X1    g059(.A(G134gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(G127gat), .ZN(new_n262_));
  INV_X1    g061(.A(G127gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(G134gat), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n262_), .A2(new_n264_), .A3(KEYINPUT80), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT80), .B1(new_n262_), .B2(new_n264_), .ZN(new_n267_));
  OAI21_X1  g066(.A(G113gat), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT80), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n263_), .A2(G134gat), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n261_), .A2(G127gat), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n269_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(G113gat), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(new_n273_), .A3(new_n265_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n268_), .A2(new_n274_), .A3(G120gat), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(G120gat), .B1(new_n268_), .B2(new_n274_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n260_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NOR3_X1   g078(.A1(new_n276_), .A2(new_n277_), .A3(new_n260_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT81), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n259_), .A2(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n257_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n281_), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n256_), .A2(new_n258_), .ZN(new_n287_));
  OAI22_X1  g086(.A1(new_n284_), .A2(new_n285_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT98), .B(KEYINPUT27), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT20), .ZN(new_n290_));
  NOR2_X1   g089(.A1(G197gat), .A2(G204gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT89), .ZN(new_n292_));
  INV_X1    g091(.A(G204gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n291_), .B1(new_n296_), .B2(G197gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G211gat), .B(G218gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT21), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n298_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n296_), .A2(G197gat), .ZN(new_n304_));
  INV_X1    g103(.A(new_n291_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(KEYINPUT90), .B(KEYINPUT21), .Z(new_n307_));
  AOI21_X1  g106(.A(new_n303_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(G197gat), .B1(new_n294_), .B2(new_n295_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT88), .ZN(new_n310_));
  INV_X1    g109(.A(G197gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n310_), .B1(new_n311_), .B2(G204gat), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n293_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT21), .B1(new_n309_), .B2(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n302_), .B1(new_n308_), .B2(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n226_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n317_));
  AND3_X1   g116(.A1(new_n317_), .A2(new_n240_), .A3(new_n244_), .ZN(new_n318_));
  XOR2_X1   g117(.A(KEYINPUT25), .B(G183gat), .Z(new_n319_));
  INV_X1    g118(.A(KEYINPUT91), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n207_), .A2(KEYINPUT91), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT92), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n242_), .A2(KEYINPUT26), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n242_), .A2(KEYINPUT26), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n323_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n208_), .A2(KEYINPUT92), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n321_), .A2(new_n322_), .A3(new_n326_), .A4(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n243_), .ZN(new_n329_));
  OR2_X1    g128(.A1(new_n225_), .A2(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n234_), .A2(new_n235_), .ZN(new_n331_));
  AOI22_X1  g130(.A1(new_n318_), .A2(new_n328_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n290_), .B1(new_n316_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n228_), .A2(new_n246_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n307_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n315_), .B(new_n298_), .C1(new_n297_), .C2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n301_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n334_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G226gat), .A2(G233gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT19), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  AND3_X1   g140(.A1(new_n333_), .A2(new_n338_), .A3(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n318_), .A2(new_n328_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n330_), .A2(new_n331_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n290_), .B1(new_n345_), .B2(new_n337_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n316_), .A2(new_n228_), .A3(new_n246_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n341_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(G92gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G8gat), .B(G36gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT18), .ZN(new_n351_));
  INV_X1    g150(.A(G64gat), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT18), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n350_), .B(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n355_), .A2(G64gat), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n349_), .B1(new_n353_), .B2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(G64gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n351_), .A2(new_n352_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n358_), .A2(new_n359_), .A3(G92gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  NOR3_X1   g160(.A1(new_n342_), .A2(new_n348_), .A3(new_n361_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n357_), .A2(new_n360_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n334_), .A2(new_n337_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT20), .B1(new_n316_), .B2(new_n332_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n340_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n333_), .A2(new_n338_), .A3(new_n341_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n363_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n289_), .B1(new_n362_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n361_), .A2(KEYINPUT97), .ZN(new_n370_));
  OR2_X1    g169(.A1(new_n361_), .A2(KEYINPUT97), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n346_), .A2(new_n341_), .A3(new_n347_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n341_), .B1(new_n333_), .B2(new_n338_), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n370_), .B(new_n371_), .C1(new_n372_), .C2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n366_), .A2(new_n363_), .A3(new_n367_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(KEYINPUT27), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n369_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G228gat), .A2(G233gat), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT29), .ZN(new_n380_));
  INV_X1    g179(.A(G155gat), .ZN(new_n381_));
  INV_X1    g180(.A(G162gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G155gat), .A2(G162gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n385_), .A2(KEYINPUT1), .ZN(new_n386_));
  OR2_X1    g185(.A1(G141gat), .A2(G148gat), .ZN(new_n387_));
  NAND3_X1  g186(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G141gat), .A2(G148gat), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n387_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT82), .B1(new_n386_), .B2(new_n390_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n387_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT82), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n392_), .B(new_n393_), .C1(KEYINPUT1), .C2(new_n385_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n391_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n385_), .B(KEYINPUT84), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n387_), .A2(KEYINPUT83), .A3(KEYINPUT3), .ZN(new_n397_));
  NOR2_X1   g196(.A1(G141gat), .A2(G148gat), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT3), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT2), .ZN(new_n400_));
  AOI22_X1  g199(.A1(new_n398_), .A2(new_n399_), .B1(new_n389_), .B2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT83), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n403_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n397_), .A2(new_n401_), .A3(new_n402_), .A4(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n396_), .A2(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n380_), .B1(new_n395_), .B2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n379_), .B1(new_n407_), .B2(new_n316_), .ZN(new_n408_));
  AOI22_X1  g207(.A1(new_n391_), .A2(new_n394_), .B1(new_n396_), .B2(new_n405_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n337_), .B(new_n378_), .C1(new_n409_), .C2(new_n380_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G78gat), .B(G106gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n395_), .A2(new_n406_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n415_), .B1(new_n416_), .B2(KEYINPUT29), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n409_), .A2(new_n380_), .A3(new_n414_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G22gat), .B(G50gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT86), .B(KEYINPUT87), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n417_), .A2(new_n418_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n421_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n414_), .B1(new_n409_), .B2(new_n380_), .ZN(new_n424_));
  AND4_X1   g223(.A1(new_n380_), .A2(new_n395_), .A3(new_n406_), .A4(new_n414_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n423_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n412_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n408_), .A2(new_n410_), .A3(new_n427_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n413_), .A2(new_n422_), .A3(new_n426_), .A4(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n426_), .A2(new_n422_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n408_), .A2(new_n427_), .A3(new_n410_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n427_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n430_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n429_), .A2(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n377_), .A2(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n416_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n436_));
  INV_X1    g235(.A(G120gat), .ZN(new_n437_));
  INV_X1    g236(.A(new_n274_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n273_), .B1(new_n272_), .B2(new_n265_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n437_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n409_), .A2(new_n440_), .A3(new_n275_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G225gat), .A2(G233gat), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n436_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n436_), .A2(KEYINPUT4), .A3(new_n441_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n442_), .B(KEYINPUT93), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n445_), .B1(new_n436_), .B2(KEYINPUT4), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n443_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n447_));
  XOR2_X1   g246(.A(G1gat), .B(G29gat), .Z(new_n448_));
  XNOR2_X1  g247(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G57gat), .B(G85gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n447_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n452_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n443_), .B(new_n454_), .C1(new_n444_), .C2(new_n446_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n288_), .A2(new_n435_), .A3(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT99), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n453_), .A2(new_n429_), .A3(new_n433_), .A4(new_n455_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n460_), .B1(new_n377_), .B2(new_n461_), .ZN(new_n462_));
  AND4_X1   g261(.A1(new_n453_), .A2(new_n429_), .A3(new_n455_), .A4(new_n433_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n463_), .A2(KEYINPUT99), .A3(new_n369_), .A4(new_n376_), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n363_), .A2(KEYINPUT32), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n465_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n363_), .A2(KEYINPUT32), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n366_), .A2(new_n467_), .A3(new_n367_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n469_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n361_), .B1(new_n342_), .B2(new_n348_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n436_), .A2(new_n441_), .A3(new_n445_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n442_), .B1(new_n436_), .B2(KEYINPUT4), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n452_), .B(new_n472_), .C1(new_n444_), .C2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n471_), .A2(new_n474_), .A3(new_n375_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n455_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n475_), .B1(KEYINPUT33), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT96), .ZN(new_n478_));
  XOR2_X1   g277(.A(KEYINPUT95), .B(KEYINPUT33), .Z(new_n479_));
  AND3_X1   g278(.A1(new_n455_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n478_), .B1(new_n455_), .B2(new_n479_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n470_), .B1(new_n477_), .B2(new_n482_), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n462_), .B(new_n464_), .C1(new_n483_), .C2(new_n434_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n288_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n459_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G15gat), .B(G22gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G1gat), .A2(G8gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT14), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(G1gat), .ZN(new_n491_));
  INV_X1    g290(.A(G8gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n488_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n490_), .A2(new_n494_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n487_), .A2(new_n488_), .A3(new_n493_), .A4(new_n489_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(G36gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(G29gat), .ZN(new_n499_));
  INV_X1    g298(.A(G29gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(G36gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(G50gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(G43gat), .ZN(new_n504_));
  INV_X1    g303(.A(G43gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(G50gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n502_), .A2(new_n507_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n499_), .A2(new_n501_), .A3(new_n504_), .A4(new_n506_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n497_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n510_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G229gat), .A2(G233gat), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n497_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT15), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT67), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n508_), .A2(new_n520_), .A3(new_n509_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n520_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n519_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n509_), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n499_), .A2(new_n501_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT67), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n508_), .A2(new_n520_), .A3(new_n509_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n526_), .A2(KEYINPUT15), .A3(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n518_), .B1(new_n523_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n513_), .A2(new_n515_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n517_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G169gat), .B(G197gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT72), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G113gat), .B(G141gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n533_), .B(new_n534_), .Z(new_n535_));
  NAND2_X1  g334(.A1(new_n531_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n535_), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n537_), .B(new_n517_), .C1(new_n529_), .C2(new_n530_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT73), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n536_), .A2(KEYINPUT73), .A3(new_n538_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n486_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT13), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G120gat), .B(G148gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(new_n293_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT5), .B(G176gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n550_), .A2(KEYINPUT65), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G230gat), .A2(G233gat), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G99gat), .A2(G106gat), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT6), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  OR2_X1    g357(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n559_));
  INV_X1    g358(.A(G106gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n559_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G85gat), .A2(G92gat), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n563_), .A2(KEYINPUT9), .ZN(new_n564_));
  OR2_X1    g363(.A1(G85gat), .A2(G92gat), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n565_), .A2(KEYINPUT9), .A3(new_n563_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n558_), .A2(new_n562_), .A3(new_n564_), .A4(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT7), .ZN(new_n568_));
  INV_X1    g367(.A(G99gat), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(new_n569_), .A3(new_n560_), .ZN(new_n570_));
  OAI21_X1  g369(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n570_), .A2(new_n556_), .A3(new_n557_), .A4(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT8), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n565_), .A2(new_n563_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n573_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n567_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G57gat), .B(G64gat), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT11), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT11), .ZN(new_n580_));
  INV_X1    g379(.A(G57gat), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n581_), .A2(G64gat), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n352_), .A2(G57gat), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n580_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G71gat), .B(G78gat), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n579_), .A2(new_n584_), .A3(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n578_), .A2(new_n585_), .A3(KEYINPUT11), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n577_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n587_), .A2(new_n588_), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n591_), .B(new_n567_), .C1(new_n576_), .C2(new_n575_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n590_), .A2(KEYINPUT12), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT12), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n577_), .A2(new_n594_), .A3(new_n589_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n553_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT64), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  AOI211_X1 g397(.A(KEYINPUT64), .B(new_n553_), .C1(new_n593_), .C2(new_n595_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n590_), .A2(new_n592_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(new_n553_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n551_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(KEYINPUT12), .B1(new_n577_), .B2(new_n589_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n572_), .A2(new_n574_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT8), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n591_), .B1(new_n608_), .B2(new_n567_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n604_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n595_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n552_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT64), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n596_), .A2(new_n597_), .ZN(new_n614_));
  AND4_X1   g413(.A1(new_n602_), .A2(new_n613_), .A3(new_n614_), .A4(new_n551_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n545_), .B1(new_n603_), .B2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n613_), .A2(new_n602_), .A3(new_n614_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n551_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n600_), .A2(new_n602_), .A3(new_n551_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(new_n620_), .A3(KEYINPUT13), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n616_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n591_), .B(new_n497_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(G231gat), .A2(G233gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT69), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n623_), .B(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT71), .B(KEYINPUT16), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G127gat), .B(G155gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G183gat), .B(G211gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT17), .ZN(new_n632_));
  OR3_X1    g431(.A1(new_n631_), .A2(KEYINPUT70), .A3(new_n632_), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n626_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n631_), .A2(new_n632_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n626_), .A2(new_n633_), .A3(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(G232gat), .A2(G233gat), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT66), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT34), .ZN(new_n641_));
  AOI22_X1  g440(.A1(new_n523_), .A2(new_n528_), .B1(new_n608_), .B2(new_n567_), .ZN(new_n642_));
  OAI22_X1  g441(.A1(new_n577_), .A2(new_n511_), .B1(KEYINPUT35), .B2(new_n641_), .ZN(new_n643_));
  OAI211_X1 g442(.A(KEYINPUT35), .B(new_n641_), .C1(new_n642_), .C2(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n641_), .A2(KEYINPUT35), .ZN(new_n645_));
  INV_X1    g444(.A(new_n577_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n646_), .B2(new_n510_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n523_), .A2(new_n528_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(new_n577_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n641_), .A2(KEYINPUT35), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n647_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT68), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n644_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(G190gat), .B(G218gat), .ZN(new_n654_));
  XNOR2_X1  g453(.A(G134gat), .B(G162gat), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n656_), .A2(KEYINPUT36), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n653_), .A2(new_n658_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n644_), .A2(new_n651_), .A3(new_n652_), .A4(new_n657_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n656_), .A2(KEYINPUT36), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n662_), .B1(new_n644_), .B2(new_n651_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT37), .B1(new_n661_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT37), .ZN(new_n666_));
  AOI211_X1 g465(.A(new_n666_), .B(new_n663_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n637_), .B1(new_n665_), .B2(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n622_), .A2(new_n668_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n544_), .A2(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n670_), .A2(new_n491_), .A3(new_n456_), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n671_), .A2(KEYINPUT100), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(KEYINPUT100), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT38), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n672_), .A2(KEYINPUT38), .A3(new_n673_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n663_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n486_), .A2(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(KEYINPUT101), .B1(new_n622_), .B2(new_n543_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT101), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n536_), .A2(KEYINPUT73), .A3(new_n538_), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT73), .B1(new_n536_), .B2(new_n538_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n616_), .A2(new_n682_), .A3(new_n621_), .A4(new_n685_), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n681_), .A2(new_n637_), .A3(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n680_), .A2(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(G1gat), .B1(new_n688_), .B2(new_n457_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n676_), .A2(new_n677_), .A3(new_n689_), .ZN(G1324gat));
  NAND3_X1  g489(.A1(new_n670_), .A2(new_n492_), .A3(new_n377_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n680_), .A2(new_n377_), .A3(new_n687_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(G8gat), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n693_), .A2(KEYINPUT39), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n693_), .A2(KEYINPUT39), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n691_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT40), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n696_), .B(new_n697_), .ZN(G1325gat));
  OAI21_X1  g497(.A(G15gat), .B1(new_n688_), .B2(new_n485_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT41), .Z(new_n700_));
  INV_X1    g499(.A(G15gat), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n670_), .A2(new_n701_), .A3(new_n288_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(G1326gat));
  INV_X1    g502(.A(new_n434_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n704_), .A2(G22gat), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT102), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n670_), .A2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n680_), .A2(new_n434_), .A3(new_n687_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(G22gat), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n709_), .A2(KEYINPUT42), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(KEYINPUT42), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT103), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n712_), .B(new_n713_), .ZN(G1327gat));
  NOR2_X1   g513(.A1(new_n678_), .A2(new_n637_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT106), .ZN(new_n716_));
  INV_X1    g515(.A(new_n622_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n544_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(new_n500_), .A3(new_n456_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n665_), .A2(new_n667_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(KEYINPUT43), .B1(new_n486_), .B2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n462_), .A2(new_n464_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n455_), .A2(new_n479_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT96), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n471_), .A2(new_n474_), .A3(new_n375_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n476_), .A2(KEYINPUT33), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n455_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n727_), .A2(new_n728_), .A3(new_n729_), .A4(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n456_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n434_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n485_), .B1(new_n725_), .B2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n458_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(new_n736_), .A3(new_n722_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n637_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n681_), .A2(new_n738_), .A3(new_n686_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT104), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n681_), .A2(KEYINPUT104), .A3(new_n738_), .A4(new_n686_), .ZN(new_n742_));
  AOI22_X1  g541(.A1(new_n724_), .A2(new_n737_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT44), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n741_), .A2(new_n742_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n736_), .B1(new_n735_), .B2(new_n722_), .ZN(new_n746_));
  AOI211_X1 g545(.A(KEYINPUT43), .B(new_n723_), .C1(new_n734_), .C2(new_n458_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n745_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT44), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n744_), .A2(new_n750_), .A3(new_n456_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT105), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n751_), .A2(new_n752_), .A3(G29gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n751_), .B2(G29gat), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n721_), .B1(new_n753_), .B2(new_n754_), .ZN(G1328gat));
  NAND2_X1  g554(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT108), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT46), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n377_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n498_), .B1(new_n761_), .B2(new_n744_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n544_), .A2(new_n498_), .A3(new_n377_), .A4(new_n718_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n763_), .B(new_n764_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n756_), .B(new_n759_), .C1(new_n762_), .C2(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n377_), .B1(new_n743_), .B2(KEYINPUT44), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n748_), .A2(new_n749_), .ZN(new_n768_));
  OAI21_X1  g567(.A(G36gat), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n764_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n763_), .B(new_n770_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n769_), .A2(new_n757_), .A3(new_n758_), .A4(new_n771_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n766_), .A2(new_n772_), .ZN(G1329gat));
  OAI21_X1  g572(.A(new_n505_), .B1(new_n719_), .B2(new_n485_), .ZN(new_n774_));
  OAI211_X1 g573(.A(G43gat), .B(new_n288_), .C1(new_n743_), .C2(KEYINPUT44), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(new_n768_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g576(.A(G50gat), .B1(new_n720_), .B2(new_n434_), .ZN(new_n778_));
  AOI211_X1 g577(.A(new_n503_), .B(new_n704_), .C1(new_n748_), .C2(new_n749_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(new_n744_), .ZN(G1331gat));
  NOR3_X1   g579(.A1(new_n717_), .A2(new_n685_), .A3(new_n738_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n680_), .A2(new_n781_), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n782_), .A2(new_n581_), .A3(new_n457_), .ZN(new_n783_));
  NOR4_X1   g582(.A1(new_n486_), .A2(new_n685_), .A3(new_n717_), .A4(new_n668_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  OR2_X1    g584(.A1(new_n785_), .A2(KEYINPUT109), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(KEYINPUT109), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(new_n456_), .A3(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n783_), .B1(new_n788_), .B2(new_n581_), .ZN(G1332gat));
  OAI21_X1  g588(.A(G64gat), .B1(new_n782_), .B2(new_n760_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT48), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n784_), .A2(new_n352_), .A3(new_n377_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(G1333gat));
  OAI21_X1  g592(.A(G71gat), .B1(new_n782_), .B2(new_n485_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT49), .ZN(new_n795_));
  OR2_X1    g594(.A1(new_n485_), .A2(G71gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n795_), .B1(new_n785_), .B2(new_n796_), .ZN(G1334gat));
  OR3_X1    g596(.A1(new_n785_), .A2(G78gat), .A3(new_n704_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n680_), .A2(new_n434_), .A3(new_n781_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(G78gat), .ZN(new_n800_));
  OR2_X1    g599(.A1(new_n800_), .A2(KEYINPUT110), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(KEYINPUT110), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n801_), .A2(KEYINPUT50), .A3(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT50), .B1(new_n801_), .B2(new_n802_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n798_), .B1(new_n803_), .B2(new_n804_), .ZN(G1335gat));
  NOR2_X1   g604(.A1(new_n717_), .A2(new_n685_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n735_), .A2(new_n716_), .A3(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(G85gat), .B1(new_n807_), .B2(new_n456_), .ZN(new_n808_));
  NOR3_X1   g607(.A1(new_n717_), .A2(new_n685_), .A3(new_n637_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n810_), .B1(new_n724_), .B2(new_n737_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n456_), .A2(G85gat), .ZN(new_n812_));
  XOR2_X1   g611(.A(new_n812_), .B(KEYINPUT111), .Z(new_n813_));
  AOI21_X1  g612(.A(new_n808_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  XOR2_X1   g613(.A(new_n814_), .B(KEYINPUT112), .Z(G1336gat));
  OAI21_X1  g614(.A(new_n809_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n816_));
  OAI21_X1  g615(.A(G92gat), .B1(new_n816_), .B2(new_n760_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n807_), .A2(new_n349_), .A3(new_n377_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(G1337gat));
  NAND4_X1  g618(.A1(new_n807_), .A2(new_n288_), .A3(new_n559_), .A4(new_n561_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n816_), .A2(new_n485_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n820_), .B1(new_n821_), .B2(new_n569_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g622(.A(G106gat), .B1(new_n816_), .B2(new_n704_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n825_));
  OR2_X1    g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n704_), .A2(G106gat), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n735_), .A2(new_n716_), .A3(new_n806_), .A4(new_n828_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(KEYINPUT113), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n830_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n831_));
  AND3_X1   g630(.A1(new_n826_), .A2(new_n827_), .A3(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n827_), .B1(new_n826_), .B2(new_n831_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n832_), .A2(new_n833_), .ZN(G1339gat));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(new_n669_), .B2(new_n543_), .ZN(new_n836_));
  NOR4_X1   g635(.A1(new_n622_), .A2(new_n668_), .A3(KEYINPUT54), .A4(new_n685_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839_));
  INV_X1    g638(.A(new_n513_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n529_), .A2(new_n840_), .A3(new_n515_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n842_));
  INV_X1    g641(.A(new_n514_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n535_), .B1(new_n843_), .B2(new_n516_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n841_), .B1(new_n842_), .B2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(new_n842_), .B2(new_n844_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n538_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n847_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n598_), .A2(new_n599_), .A3(KEYINPUT55), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n593_), .A2(new_n553_), .A3(new_n595_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT116), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n593_), .A2(new_n852_), .A3(new_n553_), .A4(new_n595_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n596_), .A2(KEYINPUT55), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n549_), .B1(new_n849_), .B2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT56), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT55), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n613_), .A2(new_n860_), .A3(new_n614_), .ZN(new_n861_));
  AOI22_X1  g660(.A1(new_n851_), .A2(new_n853_), .B1(KEYINPUT55), .B2(new_n596_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n863_), .A2(KEYINPUT56), .A3(new_n549_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n859_), .A2(new_n864_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n613_), .A2(new_n602_), .A3(new_n614_), .A4(new_n550_), .ZN(new_n866_));
  AND4_X1   g665(.A1(KEYINPUT115), .A2(new_n866_), .A3(new_n542_), .A4(new_n541_), .ZN(new_n867_));
  AOI21_X1  g666(.A(KEYINPUT115), .B1(new_n685_), .B2(new_n866_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n848_), .B1(new_n865_), .B2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n839_), .B1(new_n870_), .B2(new_n679_), .ZN(new_n871_));
  AOI21_X1  g670(.A(KEYINPUT56), .B1(new_n863_), .B2(new_n549_), .ZN(new_n872_));
  AOI211_X1 g671(.A(new_n858_), .B(new_n550_), .C1(new_n861_), .C2(new_n862_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT115), .ZN(new_n875_));
  INV_X1    g674(.A(new_n866_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(new_n543_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n685_), .A2(KEYINPUT115), .A3(new_n866_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n603_), .A2(new_n615_), .ZN(new_n880_));
  OAI22_X1  g679(.A1(new_n874_), .A2(new_n879_), .B1(new_n880_), .B2(new_n847_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n881_), .A2(KEYINPUT57), .A3(new_n678_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n847_), .A2(new_n876_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT58), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n865_), .A2(KEYINPUT58), .A3(new_n883_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n886_), .A2(new_n887_), .A3(new_n722_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n871_), .A2(new_n882_), .A3(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n838_), .B1(new_n889_), .B2(new_n738_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n434_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n485_), .A2(new_n457_), .A3(new_n377_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n893_), .A2(KEYINPUT59), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n895_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n894_), .A2(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n543_), .A2(new_n273_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT118), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n891_), .A2(new_n685_), .A3(new_n892_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(G113gat), .ZN(new_n901_));
  OAI211_X1 g700(.A(KEYINPUT118), .B(new_n273_), .C1(new_n893_), .C2(new_n543_), .ZN(new_n902_));
  AOI22_X1  g701(.A1(new_n897_), .A2(new_n898_), .B1(new_n901_), .B2(new_n902_), .ZN(G1340gat));
  INV_X1    g702(.A(new_n893_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT60), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n905_), .B1(new_n717_), .B2(G120gat), .ZN(new_n906_));
  OAI211_X1 g705(.A(new_n904_), .B(new_n906_), .C1(new_n905_), .C2(G120gat), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n894_), .A2(new_n896_), .A3(new_n717_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(new_n437_), .ZN(G1341gat));
  NAND3_X1  g708(.A1(new_n904_), .A2(new_n263_), .A3(new_n637_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n894_), .A2(new_n896_), .A3(new_n738_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n911_), .B2(new_n263_), .ZN(G1342gat));
  NAND3_X1  g711(.A1(new_n904_), .A2(new_n261_), .A3(new_n679_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n894_), .A2(new_n896_), .A3(new_n723_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n914_), .B2(new_n261_), .ZN(G1343gat));
  NAND2_X1  g714(.A1(new_n889_), .A2(new_n738_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n838_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  NOR4_X1   g717(.A1(new_n288_), .A2(new_n457_), .A3(new_n377_), .A4(new_n704_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n685_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n622_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g724(.A1(new_n920_), .A2(new_n738_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(KEYINPUT61), .B(G155gat), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(KEYINPUT119), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n926_), .B(new_n928_), .ZN(G1346gat));
  OAI21_X1  g728(.A(G162gat), .B1(new_n920_), .B2(new_n723_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n679_), .A2(new_n382_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n930_), .B1(new_n920_), .B2(new_n931_), .ZN(G1347gat));
  INV_X1    g731(.A(KEYINPUT62), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n485_), .A2(new_n456_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n934_), .A2(new_n377_), .A3(new_n685_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(KEYINPUT120), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n918_), .A2(new_n704_), .A3(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT121), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n937_), .A2(new_n938_), .A3(G169gat), .ZN(new_n939_));
  INV_X1    g738(.A(new_n939_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n938_), .B1(new_n937_), .B2(G169gat), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n933_), .B1(new_n940_), .B2(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n937_), .A2(G169gat), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(KEYINPUT121), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n944_), .A2(KEYINPUT62), .A3(new_n939_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n935_), .A2(new_n233_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n891_), .A2(new_n946_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n942_), .A2(new_n945_), .A3(new_n947_), .ZN(G1348gat));
  NAND3_X1  g747(.A1(new_n891_), .A2(new_n934_), .A3(new_n377_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n949_), .A2(new_n717_), .ZN(new_n950_));
  INV_X1    g749(.A(G176gat), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n950_), .B(new_n951_), .ZN(G1349gat));
  INV_X1    g751(.A(new_n949_), .ZN(new_n953_));
  AOI21_X1  g752(.A(G183gat), .B1(new_n953_), .B2(new_n637_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n321_), .A2(new_n322_), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n949_), .A2(new_n738_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n954_), .B1(new_n955_), .B2(new_n956_), .ZN(G1350gat));
  OAI21_X1  g756(.A(G190gat), .B1(new_n949_), .B2(new_n723_), .ZN(new_n958_));
  NAND3_X1  g757(.A1(new_n679_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n958_), .B1(new_n949_), .B2(new_n959_), .ZN(G1351gat));
  INV_X1    g759(.A(KEYINPUT123), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n485_), .A2(new_n463_), .ZN(new_n962_));
  OR2_X1    g761(.A1(new_n962_), .A2(KEYINPUT122), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n962_), .A2(KEYINPUT122), .ZN(new_n964_));
  NAND3_X1  g763(.A1(new_n963_), .A2(new_n377_), .A3(new_n964_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n965_), .B1(new_n916_), .B2(new_n917_), .ZN(new_n966_));
  INV_X1    g765(.A(new_n966_), .ZN(new_n967_));
  NOR2_X1   g766(.A1(new_n967_), .A2(new_n543_), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n961_), .B1(new_n968_), .B2(G197gat), .ZN(new_n969_));
  OAI211_X1 g768(.A(KEYINPUT123), .B(new_n311_), .C1(new_n967_), .C2(new_n543_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n968_), .A2(G197gat), .ZN(new_n971_));
  AND3_X1   g770(.A1(new_n969_), .A2(new_n970_), .A3(new_n971_), .ZN(G1352gat));
  NAND2_X1  g771(.A1(new_n966_), .A2(new_n622_), .ZN(new_n973_));
  OR3_X1    g772(.A1(new_n973_), .A2(KEYINPUT124), .A3(new_n296_), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n973_), .A2(G204gat), .ZN(new_n975_));
  OAI21_X1  g774(.A(KEYINPUT124), .B1(new_n973_), .B2(new_n296_), .ZN(new_n976_));
  NAND3_X1  g775(.A1(new_n974_), .A2(new_n975_), .A3(new_n976_), .ZN(G1353gat));
  AOI21_X1  g776(.A(new_n738_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n966_), .A2(new_n978_), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n979_), .A2(KEYINPUT125), .ZN(new_n980_));
  INV_X1    g779(.A(KEYINPUT125), .ZN(new_n981_));
  NAND3_X1  g780(.A1(new_n966_), .A2(new_n981_), .A3(new_n978_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n980_), .A2(new_n982_), .ZN(new_n983_));
  NOR2_X1   g782(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n984_));
  XNOR2_X1  g783(.A(new_n983_), .B(new_n984_), .ZN(G1354gat));
  INV_X1    g784(.A(KEYINPUT126), .ZN(new_n986_));
  AOI21_X1  g785(.A(new_n986_), .B1(new_n966_), .B2(new_n679_), .ZN(new_n987_));
  NOR4_X1   g786(.A1(new_n890_), .A2(KEYINPUT126), .A3(new_n678_), .A4(new_n965_), .ZN(new_n988_));
  NOR3_X1   g787(.A1(new_n987_), .A2(new_n988_), .A3(G218gat), .ZN(new_n989_));
  NAND2_X1  g788(.A1(new_n722_), .A2(G218gat), .ZN(new_n990_));
  NOR2_X1   g789(.A1(new_n967_), .A2(new_n990_), .ZN(new_n991_));
  OAI21_X1  g790(.A(KEYINPUT127), .B1(new_n989_), .B2(new_n991_), .ZN(new_n992_));
  INV_X1    g791(.A(KEYINPUT127), .ZN(new_n993_));
  INV_X1    g792(.A(G218gat), .ZN(new_n994_));
  NOR3_X1   g793(.A1(new_n890_), .A2(new_n678_), .A3(new_n965_), .ZN(new_n995_));
  OAI21_X1  g794(.A(new_n994_), .B1(new_n995_), .B2(new_n986_), .ZN(new_n996_));
  OAI221_X1 g795(.A(new_n993_), .B1(new_n967_), .B2(new_n990_), .C1(new_n996_), .C2(new_n988_), .ZN(new_n997_));
  NAND2_X1  g796(.A1(new_n992_), .A2(new_n997_), .ZN(G1355gat));
endmodule


