//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 0 0 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n879_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_, new_n932_, new_n933_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n963_, new_n964_,
    new_n965_;
  INV_X1    g000(.A(KEYINPUT95), .ZN(new_n202_));
  INV_X1    g001(.A(G197gat), .ZN(new_n203_));
  INV_X1    g002(.A(G204gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G197gat), .A2(G204gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT21), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n205_), .A2(KEYINPUT21), .A3(new_n206_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G211gat), .B(G218gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n210_), .A2(new_n211_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G169gat), .ZN(new_n216_));
  INV_X1    g015(.A(G176gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT24), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  NOR3_X1   g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  XOR2_X1   g020(.A(KEYINPUT25), .B(G183gat), .Z(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT26), .B(G190gat), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n221_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n220_), .A2(new_n219_), .ZN(new_n226_));
  INV_X1    g025(.A(G183gat), .ZN(new_n227_));
  INV_X1    g026(.A(G190gat), .ZN(new_n228_));
  NOR3_X1   g027(.A1(new_n227_), .A2(new_n228_), .A3(KEYINPUT23), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT23), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n225_), .A2(new_n226_), .A3(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT90), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n232_), .A2(KEYINPUT79), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT79), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n231_), .A2(new_n237_), .A3(KEYINPUT23), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(new_n230_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT89), .ZN(new_n241_));
  NOR2_X1   g040(.A1(G183gat), .A2(G190gat), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n240_), .A2(new_n241_), .A3(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n229_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT89), .B1(new_n245_), .B2(new_n242_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT22), .B(G169gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(new_n217_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n218_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n235_), .B1(new_n247_), .B2(new_n252_), .ZN(new_n253_));
  AOI211_X1 g052(.A(KEYINPUT90), .B(new_n251_), .C1(new_n244_), .C2(new_n246_), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n215_), .B(new_n234_), .C1(new_n253_), .C2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G226gat), .A2(G233gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT19), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT20), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT78), .ZN(new_n260_));
  NOR2_X1   g059(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  AND2_X1   g061(.A1(KEYINPUT77), .A2(G190gat), .ZN(new_n263_));
  NOR2_X1   g062(.A1(KEYINPUT77), .A2(G190gat), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT26), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n222_), .B1(new_n262_), .B2(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n260_), .B1(new_n266_), .B2(new_n221_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n245_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n221_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT77), .B(G190gat), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n261_), .B1(new_n270_), .B2(KEYINPUT26), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n269_), .B(KEYINPUT78), .C1(new_n271_), .C2(new_n222_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n267_), .A2(new_n268_), .A3(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n233_), .B1(new_n270_), .B2(G183gat), .ZN(new_n274_));
  INV_X1    g073(.A(new_n249_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT80), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT80), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n249_), .A2(new_n277_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n274_), .A2(new_n276_), .A3(new_n250_), .A4(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n273_), .A2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n259_), .B1(new_n280_), .B2(new_n214_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n255_), .A2(new_n258_), .A3(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n273_), .A2(new_n279_), .A3(new_n215_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT20), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n234_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n284_), .B1(new_n285_), .B2(new_n214_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n282_), .B1(new_n286_), .B2(new_n258_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G8gat), .B(G36gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT18), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G64gat), .B(G92gat), .ZN(new_n290_));
  XOR2_X1   g089(.A(new_n289_), .B(new_n290_), .Z(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n287_), .A2(new_n292_), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n291_), .B(new_n282_), .C1(new_n286_), .C2(new_n258_), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT27), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(KEYINPUT27), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n285_), .A2(new_n214_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n284_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(new_n258_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n247_), .A2(new_n252_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n300_), .A2(new_n215_), .A3(new_n234_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n281_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(new_n257_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n291_), .B1(new_n299_), .B2(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n296_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G225gat), .A2(G233gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G113gat), .B(G120gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(G134gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(G127gat), .ZN(new_n310_));
  INV_X1    g109(.A(G127gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(G134gat), .ZN(new_n312_));
  AND3_X1   g111(.A1(new_n310_), .A2(new_n312_), .A3(KEYINPUT84), .ZN(new_n313_));
  AOI21_X1  g112(.A(KEYINPUT84), .B1(new_n310_), .B2(new_n312_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n308_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT84), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n311_), .A2(G134gat), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n309_), .A2(G127gat), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n316_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n310_), .A2(new_n312_), .A3(KEYINPUT84), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(new_n320_), .A3(new_n307_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n315_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT86), .ZN(new_n323_));
  INV_X1    g122(.A(G155gat), .ZN(new_n324_));
  INV_X1    g123(.A(G162gat), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n323_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT86), .B1(G155gat), .B2(G162gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n326_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT3), .ZN(new_n330_));
  INV_X1    g129(.A(G141gat), .ZN(new_n331_));
  INV_X1    g130(.A(G148gat), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .A4(KEYINPUT87), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT87), .ZN(new_n334_));
  OAI22_X1  g133(.A1(new_n334_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G141gat), .A2(G148gat), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT2), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n333_), .A2(new_n335_), .A3(new_n338_), .A4(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n329_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n328_), .A2(KEYINPUT1), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT1), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n343_), .A2(G155gat), .A3(G162gat), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n326_), .A2(new_n342_), .A3(new_n344_), .A4(new_n327_), .ZN(new_n345_));
  XOR2_X1   g144(.A(G141gat), .B(G148gat), .Z(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n341_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n322_), .A2(new_n348_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n315_), .A2(new_n341_), .A3(new_n321_), .A4(new_n347_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(new_n350_), .A3(KEYINPUT4), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT4), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n322_), .A2(new_n348_), .A3(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n306_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G1gat), .B(G29gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G57gat), .B(G85gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n306_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n361_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n362_));
  OR3_X1    g161(.A1(new_n354_), .A2(new_n360_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT94), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n360_), .B1(new_n354_), .B2(new_n362_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n363_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  OAI211_X1 g165(.A(KEYINPUT94), .B(new_n360_), .C1(new_n354_), .C2(new_n362_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(G106gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n348_), .A2(KEYINPUT29), .ZN(new_n370_));
  INV_X1    g169(.A(G78gat), .ZN(new_n371_));
  AND2_X1   g170(.A1(G228gat), .A2(G233gat), .ZN(new_n372_));
  AOI22_X1  g171(.A1(new_n212_), .A2(new_n213_), .B1(KEYINPUT88), .B2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n370_), .A2(new_n371_), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n371_), .B1(new_n370_), .B2(new_n373_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n369_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n370_), .A2(new_n373_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(G78gat), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(G106gat), .A3(new_n374_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G22gat), .B(G50gat), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n377_), .A2(new_n380_), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n382_), .B1(new_n377_), .B2(new_n380_), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT28), .B1(new_n348_), .B2(KEYINPUT29), .ZN(new_n386_));
  OR3_X1    g185(.A1(new_n348_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n372_), .A2(KEYINPUT88), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n386_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n389_), .B1(new_n387_), .B2(new_n386_), .ZN(new_n391_));
  OAI22_X1  g190(.A1(new_n384_), .A2(new_n385_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n385_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n390_), .A2(new_n391_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n393_), .A2(new_n394_), .A3(new_n383_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n368_), .A2(new_n392_), .A3(new_n395_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n295_), .A2(new_n305_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT93), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n293_), .A2(new_n294_), .ZN(new_n399_));
  OAI211_X1 g198(.A(KEYINPUT33), .B(new_n360_), .C1(new_n354_), .C2(new_n362_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n351_), .A2(new_n306_), .A3(new_n353_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n349_), .A2(new_n350_), .A3(new_n361_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(new_n359_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n400_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT92), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT33), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n365_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n406_), .B1(new_n365_), .B2(new_n407_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n405_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n398_), .B1(new_n399_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n291_), .A2(KEYINPUT32), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n413_), .B1(new_n299_), .B2(new_n303_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n368_), .A2(new_n414_), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n282_), .B(new_n413_), .C1(new_n286_), .C2(new_n258_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n365_), .A2(new_n407_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT92), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n404_), .B1(new_n419_), .B2(new_n408_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n420_), .A2(KEYINPUT93), .A3(new_n294_), .A4(new_n293_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n412_), .A2(new_n417_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n392_), .A2(new_n395_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n397_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT30), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n280_), .B(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G15gat), .B(G43gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT81), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(G99gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G227gat), .A2(G233gat), .ZN(new_n430_));
  INV_X1    g229(.A(G71gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n429_), .B(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT83), .B1(new_n426_), .B2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n280_), .B(KEYINPUT30), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT83), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n437_), .A3(new_n433_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n435_), .A2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT82), .B1(new_n436_), .B2(new_n433_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT82), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n426_), .A2(new_n434_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n439_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT85), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT85), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n439_), .A2(new_n443_), .A3(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n322_), .B(KEYINPUT31), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n445_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  OR3_X1    g248(.A1(new_n444_), .A2(KEYINPUT85), .A3(new_n448_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n202_), .B1(new_n424_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n423_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n419_), .A2(new_n408_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n455_), .A2(new_n293_), .A3(new_n294_), .A4(new_n405_), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n456_), .A2(new_n398_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n454_), .B1(new_n457_), .B2(new_n421_), .ZN(new_n458_));
  OAI211_X1 g257(.A(KEYINPUT95), .B(new_n451_), .C1(new_n458_), .C2(new_n397_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n295_), .ZN(new_n460_));
  OR2_X1    g259(.A1(new_n296_), .A2(new_n304_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n462_), .A2(new_n454_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n452_), .A2(new_n463_), .A3(new_n368_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n453_), .A2(new_n459_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT72), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G99gat), .A2(G106gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT6), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT6), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n469_), .A2(G99gat), .A3(G106gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  OR2_X1    g270(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(new_n369_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(G85gat), .ZN(new_n475_));
  INV_X1    g274(.A(G92gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G85gat), .A2(G92gat), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(KEYINPUT9), .A3(new_n478_), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n478_), .A2(KEYINPUT9), .ZN(new_n480_));
  AND4_X1   g279(.A1(new_n471_), .A2(new_n474_), .A3(new_n479_), .A4(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT8), .ZN(new_n482_));
  INV_X1    g281(.A(G99gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n483_), .A2(new_n369_), .A3(KEYINPUT64), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT7), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT7), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n486_), .A2(new_n483_), .A3(new_n369_), .A4(KEYINPUT64), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n485_), .A2(new_n471_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n477_), .A2(new_n478_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n481_), .B1(new_n482_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT64), .ZN(new_n493_));
  NOR3_X1   g292(.A1(new_n493_), .A2(G99gat), .A3(G106gat), .ZN(new_n494_));
  AOI22_X1  g293(.A1(new_n494_), .A2(new_n486_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n489_), .B1(new_n495_), .B2(new_n485_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT8), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n492_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G29gat), .B(G36gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G43gat), .B(G50gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT15), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n498_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G232gat), .A2(G233gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT34), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT35), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT69), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n505_), .A2(KEYINPUT35), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n503_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT65), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n471_), .A2(new_n474_), .A3(new_n479_), .A4(new_n480_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n511_), .B1(new_n496_), .B2(KEYINPUT8), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n491_), .A2(new_n482_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n510_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n492_), .A2(KEYINPUT65), .A3(new_n497_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(new_n501_), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT71), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n514_), .A2(new_n515_), .A3(KEYINPUT71), .A4(new_n501_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n509_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n512_), .A2(new_n513_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT15), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n501_), .B(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(KEYINPUT70), .B1(new_n522_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT70), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n498_), .A2(new_n502_), .A3(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(new_n527_), .A3(new_n508_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n528_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n521_), .B1(new_n529_), .B2(new_n507_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G190gat), .B(G218gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G134gat), .B(G162gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n533_), .A2(KEYINPUT36), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n466_), .B1(new_n530_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n518_), .A2(new_n519_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n528_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n507_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n520_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n541_), .A2(KEYINPUT72), .A3(new_n534_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n536_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n533_), .A2(KEYINPUT36), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n530_), .A2(new_n535_), .A3(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n465_), .A2(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(G120gat), .B(G148gat), .Z(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G176gat), .B(G204gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G57gat), .B(G64gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT11), .ZN(new_n554_));
  XOR2_X1   g353(.A(G71gat), .B(G78gat), .Z(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n554_), .A2(new_n555_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n553_), .A2(KEYINPUT11), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n556_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n514_), .A2(new_n515_), .A3(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n498_), .A2(KEYINPUT12), .A3(new_n559_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n512_), .A2(new_n513_), .A3(new_n510_), .ZN(new_n564_));
  AOI21_X1  g363(.A(KEYINPUT65), .B1(new_n492_), .B2(new_n497_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n559_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT12), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G230gat), .A2(G233gat), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n563_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT66), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n514_), .A2(new_n515_), .A3(new_n571_), .A4(new_n560_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n569_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n566_), .A2(KEYINPUT66), .A3(new_n561_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n552_), .B1(new_n570_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n570_), .A2(new_n576_), .A3(new_n552_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n578_), .A2(KEYINPUT68), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT68), .ZN(new_n581_));
  INV_X1    g380(.A(new_n579_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n581_), .B1(new_n582_), .B2(new_n577_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT13), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n580_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n584_), .B1(new_n580_), .B2(new_n583_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G15gat), .B(G22gat), .ZN(new_n588_));
  INV_X1    g387(.A(G1gat), .ZN(new_n589_));
  INV_X1    g388(.A(G8gat), .ZN(new_n590_));
  OAI21_X1  g389(.A(KEYINPUT14), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n588_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G1gat), .B(G8gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n501_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n595_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(KEYINPUT75), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT75), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n594_), .A2(new_n595_), .A3(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G229gat), .A2(G233gat), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n502_), .A2(new_n594_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n605_), .A2(new_n602_), .A3(new_n596_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G113gat), .B(G141gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT76), .ZN(new_n609_));
  XOR2_X1   g408(.A(G169gat), .B(G197gat), .Z(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n607_), .B(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(G127gat), .B(G155gat), .Z(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT16), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G183gat), .B(G211gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n594_), .B(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(new_n559_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n616_), .B1(new_n619_), .B2(KEYINPUT17), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n620_), .B1(KEYINPUT17), .B2(new_n616_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n619_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(KEYINPUT74), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n621_), .B(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n587_), .A2(new_n612_), .A3(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT96), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n547_), .A2(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(G1gat), .B1(new_n627_), .B2(new_n368_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT38), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n465_), .A2(new_n612_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(KEYINPUT73), .A2(KEYINPUT37), .ZN(new_n631_));
  AOI21_X1  g430(.A(KEYINPUT72), .B1(new_n541_), .B2(new_n534_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n507_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n633_));
  NOR4_X1   g432(.A1(new_n633_), .A2(new_n466_), .A3(new_n535_), .A4(new_n520_), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n631_), .B(new_n545_), .C1(new_n632_), .C2(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(KEYINPUT73), .A2(KEYINPUT37), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n636_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n543_), .A2(new_n631_), .A3(new_n545_), .A4(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n624_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n630_), .A2(new_n642_), .A3(new_n587_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n368_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(new_n589_), .A3(new_n644_), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n645_), .A2(KEYINPUT97), .A3(new_n629_), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT97), .B1(new_n645_), .B2(new_n629_), .ZN(new_n647_));
  OAI221_X1 g446(.A(new_n628_), .B1(new_n629_), .B2(new_n645_), .C1(new_n646_), .C2(new_n647_), .ZN(G1324gat));
  XNOR2_X1  g447(.A(KEYINPUT98), .B(KEYINPUT40), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n547_), .A2(new_n462_), .A3(new_n626_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(G8gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT39), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n643_), .A2(new_n590_), .A3(new_n462_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n649_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n651_), .A2(KEYINPUT39), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT39), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n656_), .B1(new_n650_), .B2(G8gat), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n653_), .B(new_n649_), .C1(new_n655_), .C2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n654_), .A2(new_n659_), .ZN(G1325gat));
  OAI21_X1  g459(.A(G15gat), .B1(new_n627_), .B2(new_n451_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT41), .Z(new_n662_));
  INV_X1    g461(.A(G15gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n643_), .A2(new_n663_), .A3(new_n452_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(G1326gat));
  OAI21_X1  g464(.A(G22gat), .B1(new_n627_), .B2(new_n423_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT42), .ZN(new_n667_));
  INV_X1    g466(.A(G22gat), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n643_), .A2(new_n668_), .A3(new_n454_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(G1327gat));
  INV_X1    g469(.A(new_n587_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n546_), .A2(new_n624_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n671_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n630_), .A2(new_n674_), .ZN(new_n675_));
  OR3_X1    g474(.A1(new_n675_), .A2(G29gat), .A3(new_n368_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n587_), .A2(new_n612_), .A3(new_n641_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT99), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n465_), .A2(new_n679_), .A3(new_n640_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n465_), .B2(new_n640_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n678_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI211_X1 g483(.A(KEYINPUT44), .B(new_n678_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n684_), .A2(new_n644_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT100), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n686_), .A2(new_n687_), .A3(G29gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n686_), .B2(G29gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n676_), .B1(new_n688_), .B2(new_n689_), .ZN(G1328gat));
  INV_X1    g489(.A(KEYINPUT46), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT102), .B1(new_n691_), .B2(KEYINPUT101), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n684_), .A2(new_n462_), .A3(new_n685_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(G36gat), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n691_), .A2(KEYINPUT102), .ZN(new_n696_));
  INV_X1    g495(.A(new_n462_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n697_), .A2(G36gat), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n465_), .A2(new_n612_), .A3(new_n674_), .A4(new_n698_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n699_), .A2(KEYINPUT45), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(KEYINPUT45), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n696_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n693_), .B1(new_n695_), .B2(new_n703_), .ZN(new_n704_));
  AOI211_X1 g503(.A(new_n692_), .B(new_n702_), .C1(new_n694_), .C2(G36gat), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1329gat));
  NAND4_X1  g505(.A1(new_n684_), .A2(G43gat), .A3(new_n452_), .A4(new_n685_), .ZN(new_n707_));
  INV_X1    g506(.A(G43gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n708_), .B1(new_n675_), .B2(new_n451_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g510(.A1(new_n675_), .A2(G50gat), .A3(new_n423_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n684_), .A2(new_n454_), .A3(new_n685_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT103), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(G50gat), .B1(new_n713_), .B2(new_n714_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(G1331gat));
  INV_X1    g516(.A(new_n612_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n671_), .A2(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n719_), .A2(new_n641_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n547_), .A2(G57gat), .A3(new_n644_), .A4(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT104), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n721_), .A2(new_n722_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n719_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n465_), .A2(new_n725_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n726_), .A2(new_n640_), .A3(new_n641_), .ZN(new_n727_));
  AOI21_X1  g526(.A(G57gat), .B1(new_n727_), .B2(new_n644_), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n723_), .A2(new_n724_), .A3(new_n728_), .ZN(G1332gat));
  NAND2_X1  g528(.A1(new_n547_), .A2(new_n720_), .ZN(new_n730_));
  OAI21_X1  g529(.A(G64gat), .B1(new_n730_), .B2(new_n697_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT48), .ZN(new_n732_));
  INV_X1    g531(.A(new_n727_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n697_), .A2(G64gat), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT105), .Z(new_n735_));
  OAI21_X1  g534(.A(new_n732_), .B1(new_n733_), .B2(new_n735_), .ZN(G1333gat));
  NAND3_X1  g535(.A1(new_n727_), .A2(new_n431_), .A3(new_n452_), .ZN(new_n737_));
  OAI21_X1  g536(.A(G71gat), .B1(new_n730_), .B2(new_n451_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(KEYINPUT49), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(KEYINPUT49), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n737_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT106), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  OAI211_X1 g542(.A(KEYINPUT106), .B(new_n737_), .C1(new_n739_), .C2(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1334gat));
  OAI21_X1  g544(.A(G78gat), .B1(new_n730_), .B2(new_n423_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT50), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n727_), .A2(new_n371_), .A3(new_n454_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1335gat));
  NOR2_X1   g548(.A1(new_n726_), .A2(new_n673_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n750_), .A2(new_n475_), .A3(new_n644_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n680_), .A2(new_n681_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n719_), .A2(new_n624_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(new_n644_), .A3(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n755_), .B2(new_n475_), .ZN(G1336gat));
  NAND3_X1  g555(.A1(new_n752_), .A2(new_n462_), .A3(new_n753_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(G92gat), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n750_), .A2(new_n476_), .A3(new_n462_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT107), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n758_), .A2(new_n759_), .A3(KEYINPUT107), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1337gat));
  AND4_X1   g563(.A1(new_n452_), .A2(new_n750_), .A3(new_n472_), .A4(new_n473_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n752_), .A2(new_n452_), .A3(new_n753_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(G99gat), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n767_), .A2(KEYINPUT108), .A3(KEYINPUT51), .ZN(new_n768_));
  NOR2_X1   g567(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n769_));
  AND2_X1   g568(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n767_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n768_), .A2(new_n771_), .ZN(G1338gat));
  NAND3_X1  g571(.A1(new_n750_), .A2(new_n369_), .A3(new_n454_), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n753_), .B(new_n454_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n774_), .A2(new_n775_), .A3(G106gat), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n774_), .B2(G106gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT53), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n773_), .B(new_n780_), .C1(new_n776_), .C2(new_n777_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1339gat));
  NAND3_X1  g581(.A1(new_n452_), .A2(new_n463_), .A3(new_n644_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n783_), .A2(KEYINPUT59), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n587_), .A2(new_n639_), .A3(new_n637_), .A4(new_n624_), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT54), .B1(new_n785_), .B2(new_n612_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n642_), .A2(new_n787_), .A3(new_n718_), .A4(new_n587_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n612_), .A2(new_n579_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n552_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n560_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n561_), .B(new_n562_), .C1(new_n794_), .C2(KEYINPUT12), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n793_), .B1(new_n795_), .B2(new_n573_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n795_), .A2(new_n573_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n795_), .A2(new_n793_), .A3(new_n573_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n792_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT56), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(KEYINPUT56), .B(new_n792_), .C1(new_n798_), .C2(new_n799_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n791_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n607_), .A2(new_n611_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n601_), .A2(new_n602_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n611_), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n807_), .A2(KEYINPUT109), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n605_), .A2(new_n603_), .A3(new_n596_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n809_), .B1(new_n807_), .B2(KEYINPUT109), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n805_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n580_), .A2(new_n583_), .A3(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n546_), .B1(new_n804_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT110), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n814_), .A2(KEYINPUT57), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n813_), .A2(new_n816_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n546_), .B(new_n815_), .C1(new_n804_), .C2(new_n812_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n803_), .A2(KEYINPUT111), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n569_), .B1(new_n563_), .B2(new_n568_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n570_), .B1(new_n821_), .B2(new_n793_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n799_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT111), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n824_), .A2(new_n825_), .A3(KEYINPUT56), .A4(new_n792_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n820_), .A2(new_n826_), .A3(new_n802_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n811_), .A2(new_n579_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT58), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n827_), .A2(KEYINPUT58), .A3(new_n828_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n640_), .A3(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n624_), .B1(new_n819_), .B2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n784_), .B1(new_n790_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n832_), .A2(new_n640_), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT58), .B1(new_n827_), .B2(new_n828_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT112), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT112), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n831_), .A2(new_n839_), .A3(new_n640_), .A4(new_n832_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n838_), .A2(new_n840_), .A3(new_n819_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n641_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n783_), .B1(new_n842_), .B2(new_n789_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n612_), .B(new_n835_), .C1(new_n843_), .C2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(G113gat), .ZN(new_n846_));
  INV_X1    g645(.A(G113gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n843_), .A2(new_n847_), .A3(new_n612_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n846_), .A2(KEYINPUT113), .A3(new_n848_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1340gat));
  OAI211_X1 g652(.A(new_n671_), .B(new_n835_), .C1(new_n843_), .C2(new_n844_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(G120gat), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n587_), .A2(KEYINPUT60), .ZN(new_n856_));
  MUX2_X1   g655(.A(new_n856_), .B(KEYINPUT60), .S(G120gat), .Z(new_n857_));
  NAND2_X1  g656(.A1(new_n843_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n855_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n855_), .A2(KEYINPUT114), .A3(new_n858_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1341gat));
  OAI21_X1  g662(.A(new_n835_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n864_));
  OAI21_X1  g663(.A(G127gat), .B1(new_n864_), .B2(new_n641_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n843_), .A2(new_n311_), .A3(new_n624_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(G1342gat));
  INV_X1    g666(.A(new_n640_), .ZN(new_n868_));
  OAI21_X1  g667(.A(G134gat), .B1(new_n864_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n546_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n843_), .A2(new_n309_), .A3(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(G1343gat));
  NAND2_X1  g671(.A1(new_n842_), .A2(new_n789_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n451_), .A2(new_n697_), .A3(new_n454_), .A4(new_n644_), .ZN(new_n874_));
  XOR2_X1   g673(.A(new_n874_), .B(KEYINPUT115), .Z(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n718_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(new_n331_), .ZN(G1344gat));
  NOR2_X1   g677(.A1(new_n876_), .A2(new_n587_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(new_n332_), .ZN(G1345gat));
  OR3_X1    g679(.A1(new_n876_), .A2(KEYINPUT116), .A3(new_n641_), .ZN(new_n881_));
  OAI21_X1  g680(.A(KEYINPUT116), .B1(new_n876_), .B2(new_n641_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT61), .B(G155gat), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n881_), .A2(new_n882_), .A3(new_n884_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1346gat));
  OAI21_X1  g687(.A(G162gat), .B1(new_n876_), .B2(new_n868_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n870_), .A2(new_n325_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n876_), .B2(new_n890_), .ZN(G1347gat));
  INV_X1    g690(.A(KEYINPUT121), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT117), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n644_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n452_), .A2(new_n894_), .A3(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n462_), .A2(new_n368_), .ZN(new_n897_));
  OAI21_X1  g696(.A(KEYINPUT117), .B1(new_n897_), .B2(new_n451_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n718_), .B1(new_n896_), .B2(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n454_), .B1(new_n899_), .B2(KEYINPUT118), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n894_), .B1(new_n452_), .B2(new_n895_), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n897_), .A2(new_n451_), .A3(KEYINPUT117), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n612_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT118), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n900_), .A2(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n834_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n789_), .B2(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n893_), .B1(new_n908_), .B2(new_n216_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n790_), .A2(new_n834_), .ZN(new_n910_));
  OAI211_X1 g709(.A(KEYINPUT119), .B(G169gat), .C1(new_n910_), .C2(new_n906_), .ZN(new_n911_));
  AND3_X1   g710(.A1(new_n909_), .A2(KEYINPUT62), .A3(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n907_), .A2(new_n789_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n901_), .A2(new_n902_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n914_), .A2(new_n454_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n913_), .A2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n612_), .A2(new_n248_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(KEYINPUT120), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT62), .ZN(new_n921_));
  OAI211_X1 g720(.A(new_n893_), .B(new_n921_), .C1(new_n908_), .C2(new_n216_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n920_), .A2(new_n922_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n892_), .B1(new_n912_), .B2(new_n923_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n909_), .A2(KEYINPUT62), .A3(new_n911_), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n925_), .A2(KEYINPUT121), .A3(new_n922_), .A4(new_n920_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n926_), .ZN(G1348gat));
  AOI21_X1  g726(.A(G176gat), .B1(new_n917_), .B2(new_n671_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n454_), .B1(new_n842_), .B2(new_n789_), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n914_), .A2(new_n217_), .A3(new_n587_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n928_), .B1(new_n929_), .B2(new_n930_), .ZN(G1349gat));
  NOR3_X1   g730(.A1(new_n916_), .A2(new_n223_), .A3(new_n641_), .ZN(new_n932_));
  OAI211_X1 g731(.A(new_n929_), .B(new_n624_), .C1(new_n902_), .C2(new_n901_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n932_), .B1(new_n227_), .B2(new_n933_), .ZN(G1350gat));
  NAND3_X1  g733(.A1(new_n917_), .A2(new_n224_), .A3(new_n870_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n917_), .A2(new_n640_), .ZN(new_n936_));
  AND3_X1   g735(.A1(new_n936_), .A2(KEYINPUT122), .A3(G190gat), .ZN(new_n937_));
  AOI21_X1  g736(.A(KEYINPUT122), .B1(new_n936_), .B2(G190gat), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n935_), .B1(new_n937_), .B2(new_n938_), .ZN(G1351gat));
  NOR3_X1   g738(.A1(new_n452_), .A2(new_n897_), .A3(new_n423_), .ZN(new_n940_));
  AND2_X1   g739(.A1(new_n873_), .A2(new_n940_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(new_n612_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n942_), .A2(new_n203_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n943_), .A2(new_n944_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n942_), .A2(KEYINPUT124), .A3(new_n203_), .ZN(new_n946_));
  OAI21_X1  g745(.A(KEYINPUT123), .B1(new_n942_), .B2(new_n203_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT123), .ZN(new_n948_));
  NAND4_X1  g747(.A1(new_n941_), .A2(new_n948_), .A3(G197gat), .A4(new_n612_), .ZN(new_n949_));
  AOI22_X1  g748(.A1(new_n945_), .A2(new_n946_), .B1(new_n947_), .B2(new_n949_), .ZN(G1352gat));
  NAND2_X1  g749(.A1(new_n941_), .A2(new_n671_), .ZN(new_n951_));
  INV_X1    g750(.A(KEYINPUT125), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n951_), .B1(new_n952_), .B2(G204gat), .ZN(new_n953_));
  XNOR2_X1  g752(.A(KEYINPUT125), .B(G204gat), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n953_), .B1(new_n951_), .B2(new_n954_), .ZN(G1353gat));
  AND3_X1   g754(.A1(new_n873_), .A2(new_n624_), .A3(new_n940_), .ZN(new_n956_));
  XOR2_X1   g755(.A(KEYINPUT63), .B(G211gat), .Z(new_n957_));
  AOI21_X1  g756(.A(KEYINPUT126), .B1(new_n956_), .B2(new_n957_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n956_), .A2(new_n957_), .ZN(new_n959_));
  OR2_X1    g758(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n959_), .B1(new_n960_), .B2(new_n956_), .ZN(new_n961_));
  AOI21_X1  g760(.A(new_n958_), .B1(new_n961_), .B2(KEYINPUT126), .ZN(G1354gat));
  AOI21_X1  g761(.A(G218gat), .B1(new_n941_), .B2(new_n870_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n640_), .A2(G218gat), .ZN(new_n964_));
  XNOR2_X1  g763(.A(new_n964_), .B(KEYINPUT127), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n963_), .B1(new_n941_), .B2(new_n965_), .ZN(G1355gat));
endmodule


