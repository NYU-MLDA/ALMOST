//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 0 1 0 0 1 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202_));
  INV_X1    g001(.A(G183gat), .ZN(new_n203_));
  INV_X1    g002(.A(G190gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT23), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n206_), .A2(G183gat), .A3(G190gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT80), .ZN(new_n208_));
  AND2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n207_), .A2(new_n208_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n205_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT26), .B(G190gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT25), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n203_), .A2(KEYINPUT78), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT78), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(G183gat), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n213_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n212_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(G169gat), .ZN(new_n220_));
  INV_X1    g019(.A(G176gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(new_n221_), .A3(KEYINPUT79), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT79), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n223_), .B1(G169gat), .B2(G176gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n222_), .A2(new_n224_), .A3(KEYINPUT24), .A4(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n222_), .A2(new_n224_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT24), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n211_), .A2(new_n219_), .A3(new_n226_), .A4(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n205_), .A2(new_n207_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n214_), .A2(new_n216_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n231_), .B1(new_n232_), .B2(G190gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT22), .B(G169gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(new_n221_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n225_), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n230_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT30), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT81), .ZN(new_n239_));
  INV_X1    g038(.A(G227gat), .ZN(new_n240_));
  INV_X1    g039(.A(G233gat), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n239_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n239_), .A2(new_n242_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n202_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n245_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n202_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n247_), .A2(new_n243_), .A3(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT82), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G127gat), .B(G134gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G113gat), .B(G120gat), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n252_), .A2(new_n253_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n251_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n252_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n253_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n252_), .A2(new_n253_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(KEYINPUT82), .A3(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n256_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT31), .ZN(new_n263_));
  XOR2_X1   g062(.A(G71gat), .B(G99gat), .Z(new_n264_));
  XOR2_X1   g063(.A(new_n263_), .B(new_n264_), .Z(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n250_), .A2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n246_), .A2(new_n249_), .A3(new_n265_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  AND3_X1   g068(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n270_));
  INV_X1    g069(.A(G141gat), .ZN(new_n271_));
  INV_X1    g070(.A(G148gat), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(new_n272_), .A3(KEYINPUT3), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT3), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n274_), .B1(G141gat), .B2(G148gat), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n270_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT2), .ZN(new_n277_));
  AND3_X1   g076(.A1(KEYINPUT83), .A2(G141gat), .A3(G148gat), .ZN(new_n278_));
  AOI21_X1  g077(.A(KEYINPUT83), .B1(G141gat), .B2(G148gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n277_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n276_), .A2(new_n280_), .ZN(new_n281_));
  AND2_X1   g080(.A1(G155gat), .A2(G162gat), .ZN(new_n282_));
  NOR2_X1   g081(.A1(G155gat), .A2(G162gat), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n281_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n271_), .A2(new_n272_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n286_), .B(new_n287_), .C1(new_n278_), .C2(new_n279_), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n282_), .A2(new_n283_), .A3(KEYINPUT1), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n285_), .A2(KEYINPUT84), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT84), .ZN(new_n292_));
  INV_X1    g091(.A(new_n284_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n293_), .B1(new_n276_), .B2(new_n280_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n288_), .A2(new_n289_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n292_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n291_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n298_), .A2(KEYINPUT29), .ZN(new_n299_));
  INV_X1    g098(.A(G218gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(G211gat), .ZN(new_n301_));
  INV_X1    g100(.A(G211gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(G218gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(G204gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(G197gat), .ZN(new_n306_));
  INV_X1    g105(.A(G197gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(G204gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n304_), .B1(KEYINPUT21), .B2(new_n309_), .ZN(new_n310_));
  OR3_X1    g109(.A1(new_n307_), .A2(KEYINPUT87), .A3(G204gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n306_), .A2(KEYINPUT87), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT21), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n311_), .A2(new_n312_), .A3(new_n313_), .A4(new_n308_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n311_), .A2(new_n312_), .A3(new_n308_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n313_), .B1(new_n301_), .B2(new_n303_), .ZN(new_n316_));
  AOI22_X1  g115(.A1(new_n310_), .A2(new_n314_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G228gat), .A2(G233gat), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n318_), .B(KEYINPUT86), .Z(new_n319_));
  NOR2_X1   g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT29), .B1(new_n294_), .B2(new_n295_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n291_), .A2(new_n296_), .A3(KEYINPUT29), .ZN(new_n323_));
  INV_X1    g122(.A(new_n317_), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n319_), .ZN(new_n326_));
  OAI211_X1 g125(.A(G78gat), .B(new_n322_), .C1(new_n325_), .C2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(G78gat), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n326_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n322_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n328_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n327_), .A2(G106gat), .A3(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT85), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(G106gat), .B1(new_n327_), .B2(new_n331_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n299_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n327_), .A2(new_n331_), .ZN(new_n337_));
  INV_X1    g136(.A(G106gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n299_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n339_), .A2(new_n333_), .A3(new_n340_), .A4(new_n332_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G22gat), .B(G50gat), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n342_), .B(KEYINPUT28), .Z(new_n343_));
  AND3_X1   g142(.A1(new_n336_), .A2(new_n341_), .A3(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n343_), .B1(new_n336_), .B2(new_n341_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G226gat), .A2(G233gat), .ZN(new_n347_));
  XOR2_X1   g146(.A(new_n347_), .B(KEYINPUT88), .Z(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT19), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n230_), .A2(new_n317_), .A3(new_n236_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(KEYINPUT89), .A3(KEYINPUT20), .ZN(new_n352_));
  INV_X1    g151(.A(new_n212_), .ZN(new_n353_));
  XOR2_X1   g152(.A(KEYINPUT25), .B(G183gat), .Z(new_n354_));
  OAI21_X1  g153(.A(new_n226_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n220_), .A2(new_n221_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n231_), .B1(KEYINPUT24), .B2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT90), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT90), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n231_), .B(new_n359_), .C1(KEYINPUT24), .C2(new_n356_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n355_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n235_), .A2(new_n225_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n203_), .A2(new_n204_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n362_), .B1(new_n211_), .B2(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n324_), .B1(new_n361_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n352_), .A2(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(KEYINPUT89), .B1(new_n351_), .B2(KEYINPUT20), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n350_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT20), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n361_), .A2(new_n364_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n369_), .B1(new_n370_), .B2(new_n317_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n237_), .A2(new_n324_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(new_n349_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n368_), .A2(new_n373_), .ZN(new_n374_));
  XOR2_X1   g173(.A(KEYINPUT91), .B(KEYINPUT18), .Z(new_n375_));
  XNOR2_X1  g174(.A(G64gat), .B(G92gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G8gat), .B(G36gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT92), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n377_), .B(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n374_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT93), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n368_), .A2(new_n380_), .A3(new_n373_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT98), .B(KEYINPUT27), .ZN(new_n386_));
  INV_X1    g185(.A(new_n374_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n387_), .A2(KEYINPUT93), .A3(new_n380_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n385_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n371_), .A2(new_n372_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  OR2_X1    g190(.A1(new_n366_), .A2(new_n367_), .ZN(new_n392_));
  MUX2_X1   g191(.A(new_n391_), .B(new_n392_), .S(new_n349_), .Z(new_n393_));
  OAI211_X1 g192(.A(KEYINPUT27), .B(new_n384_), .C1(new_n393_), .C2(new_n380_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n389_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n262_), .A2(new_n291_), .A3(new_n296_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n285_), .B(new_n290_), .C1(new_n254_), .C2(new_n255_), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n396_), .A2(new_n397_), .A3(KEYINPUT4), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT4), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n262_), .A2(new_n291_), .A3(new_n296_), .A4(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G225gat), .A2(G233gat), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT94), .B1(new_n398_), .B2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n396_), .A2(new_n397_), .A3(KEYINPUT4), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT94), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n405_), .A2(new_n406_), .A3(new_n402_), .A4(new_n400_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n396_), .A2(new_n397_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n408_), .A2(new_n402_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n404_), .A2(new_n407_), .A3(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G1gat), .B(G29gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(KEYINPUT0), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(G57gat), .ZN(new_n414_));
  OR2_X1    g213(.A1(new_n412_), .A2(KEYINPUT0), .ZN(new_n415_));
  INV_X1    g214(.A(G57gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n412_), .A2(KEYINPUT0), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n414_), .A2(new_n418_), .A3(G85gat), .ZN(new_n419_));
  AOI21_X1  g218(.A(G85gat), .B1(new_n414_), .B2(new_n418_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(KEYINPUT96), .B1(new_n411_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n421_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n404_), .A2(new_n423_), .A3(new_n410_), .A4(new_n407_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n404_), .A2(new_n410_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n426_), .A2(KEYINPUT96), .A3(new_n423_), .A4(new_n407_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NOR4_X1   g228(.A1(new_n269_), .A2(new_n346_), .A3(new_n395_), .A4(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT33), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n424_), .A2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n421_), .B1(new_n408_), .B2(new_n401_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT95), .ZN(new_n434_));
  OR2_X1    g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n400_), .A2(new_n401_), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n433_), .A2(new_n434_), .B1(new_n436_), .B2(new_n405_), .ZN(new_n437_));
  AOI22_X1  g236(.A1(new_n424_), .A2(new_n431_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n368_), .A2(new_n380_), .A3(new_n373_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n380_), .B1(new_n368_), .B2(new_n373_), .ZN(new_n440_));
  NOR3_X1   g239(.A1(new_n439_), .A2(new_n440_), .A3(KEYINPUT93), .ZN(new_n441_));
  NOR3_X1   g240(.A1(new_n374_), .A2(new_n383_), .A3(new_n381_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n432_), .B(new_n438_), .C1(new_n441_), .C2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n390_), .A2(new_n350_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n380_), .A2(KEYINPUT32), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n444_), .B(new_n445_), .C1(new_n392_), .C2(new_n350_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n446_), .B1(new_n387_), .B2(new_n445_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n425_), .A2(new_n427_), .A3(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n443_), .A2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n449_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT97), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n336_), .A2(new_n341_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n343_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n336_), .A2(new_n341_), .A3(new_n343_), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n455_), .A2(new_n456_), .B1(new_n443_), .B2(new_n448_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT97), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n389_), .A2(new_n394_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n459_), .A2(new_n456_), .A3(new_n455_), .A4(new_n428_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n452_), .A2(new_n458_), .A3(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n430_), .B1(new_n461_), .B2(new_n269_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT74), .B(G1gat), .ZN(new_n463_));
  INV_X1    g262(.A(G8gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT14), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G15gat), .B(G22gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  XOR2_X1   g266(.A(new_n467_), .B(G1gat), .Z(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(G8gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n467_), .B(G1gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n464_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G231gat), .A2(G233gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(G71gat), .B(G78gat), .Z(new_n475_));
  XNOR2_X1  g274(.A(G57gat), .B(G64gat), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n475_), .B1(KEYINPUT11), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(KEYINPUT11), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n474_), .B(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(KEYINPUT75), .B(KEYINPUT16), .Z(new_n482_));
  XNOR2_X1  g281(.A(G127gat), .B(G155gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(G183gat), .B(G211gat), .Z(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n487_), .A2(KEYINPUT17), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n487_), .A2(KEYINPUT17), .ZN(new_n489_));
  OR3_X1    g288(.A1(new_n481_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n481_), .A2(new_n488_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT37), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G190gat), .B(G218gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G134gat), .B(G162gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G29gat), .B(G36gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G43gat), .B(G50gat), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n497_), .B(new_n498_), .Z(new_n499_));
  XOR2_X1   g298(.A(new_n499_), .B(KEYINPUT15), .Z(new_n500_));
  INV_X1    g299(.A(KEYINPUT70), .ZN(new_n501_));
  NOR2_X1   g300(.A1(G85gat), .A2(G92gat), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G85gat), .A2(G92gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n505_), .A2(KEYINPUT8), .ZN(new_n506_));
  NOR2_X1   g305(.A1(G99gat), .A2(G106gat), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT7), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n507_), .B1(KEYINPUT67), .B2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT67), .B(KEYINPUT7), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n509_), .B1(new_n510_), .B2(new_n507_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G99gat), .A2(G106gat), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT6), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n506_), .B1(new_n511_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT68), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n514_), .B1(new_n511_), .B2(new_n516_), .ZN(new_n517_));
  OAI211_X1 g316(.A(KEYINPUT68), .B(new_n509_), .C1(new_n510_), .C2(new_n507_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n505_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT8), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n515_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT69), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(KEYINPUT10), .B(G99gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT64), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n514_), .B1(new_n526_), .B2(new_n338_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n504_), .A2(KEYINPUT65), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n502_), .B1(new_n528_), .B2(KEYINPUT9), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n529_), .B1(KEYINPUT9), .B2(new_n528_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT66), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n527_), .A2(new_n531_), .ZN(new_n532_));
  OAI211_X1 g331(.A(KEYINPUT69), .B(new_n515_), .C1(new_n519_), .C2(new_n520_), .ZN(new_n533_));
  AND4_X1   g332(.A1(new_n501_), .A2(new_n523_), .A3(new_n532_), .A4(new_n533_), .ZN(new_n534_));
  AOI22_X1  g333(.A1(new_n521_), .A2(new_n522_), .B1(new_n531_), .B2(new_n527_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n501_), .B1(new_n535_), .B2(new_n533_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n500_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n521_), .A2(new_n532_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n499_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G232gat), .A2(G233gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT34), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT35), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT73), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT35), .ZN(new_n547_));
  INV_X1    g346(.A(new_n543_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n546_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n541_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n537_), .A2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n552_), .A2(new_n545_), .A3(new_n544_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n544_), .A2(new_n545_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n537_), .A2(new_n554_), .A3(new_n551_), .ZN(new_n555_));
  AOI211_X1 g354(.A(KEYINPUT36), .B(new_n496_), .C1(new_n553_), .C2(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n496_), .B(KEYINPUT36), .Z(new_n557_));
  NAND3_X1  g356(.A1(new_n553_), .A2(new_n555_), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n493_), .B1(new_n556_), .B2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n553_), .A2(new_n555_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n496_), .A2(KEYINPUT36), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n563_), .A2(KEYINPUT37), .A3(new_n558_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n560_), .A2(new_n564_), .ZN(new_n565_));
  NOR3_X1   g364(.A1(new_n462_), .A2(new_n492_), .A3(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G120gat), .B(G148gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(new_n305_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT5), .B(G176gat), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n568_), .B(new_n569_), .Z(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n479_), .A2(KEYINPUT12), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n523_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT70), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n535_), .A2(new_n501_), .A3(new_n533_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n572_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(KEYINPUT12), .B1(new_n538_), .B2(new_n479_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n539_), .A2(new_n480_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G230gat), .A2(G233gat), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NOR3_X1   g379(.A1(new_n576_), .A2(new_n577_), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n538_), .A2(new_n479_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n579_), .B1(new_n578_), .B2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n571_), .B1(new_n581_), .B2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n572_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n585_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n580_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n577_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n586_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n583_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n589_), .A2(new_n590_), .A3(new_n570_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n584_), .A2(KEYINPUT71), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT71), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n593_), .B(new_n571_), .C1(new_n581_), .C2(new_n583_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(KEYINPUT72), .B(KEYINPUT13), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n592_), .A2(new_n594_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT13), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n599_), .A2(KEYINPUT72), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n600_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n598_), .A2(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n469_), .A2(new_n471_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(new_n500_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n472_), .A2(new_n540_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(G229gat), .A2(G233gat), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n604_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT76), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n603_), .A2(new_n499_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(new_n605_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n606_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n608_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  AOI211_X1 g411(.A(KEYINPUT76), .B(new_n606_), .C1(new_n609_), .C2(new_n605_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n607_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G169gat), .B(G197gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(G141gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT77), .B(G113gat), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n616_), .B(new_n617_), .Z(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n614_), .A2(new_n619_), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n607_), .B(new_n618_), .C1(new_n612_), .C2(new_n613_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n602_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n566_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT99), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT99), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n566_), .A2(new_n627_), .A3(new_n624_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n429_), .A2(new_n463_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n631_), .A2(KEYINPUT38), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(KEYINPUT38), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n556_), .A2(new_n559_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n462_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n492_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n624_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n635_), .A2(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(G1gat), .B1(new_n639_), .B2(new_n428_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n632_), .A2(new_n633_), .A3(new_n640_), .ZN(G1324gat));
  NAND4_X1  g440(.A1(new_n626_), .A2(new_n464_), .A3(new_n395_), .A4(new_n628_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n635_), .A2(new_n638_), .A3(new_n395_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT39), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(new_n644_), .A3(G8gat), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n644_), .B1(new_n643_), .B2(G8gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n642_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT100), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT100), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n642_), .B(new_n650_), .C1(new_n647_), .C2(new_n646_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n649_), .A2(KEYINPUT40), .A3(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(KEYINPUT40), .B1(new_n649_), .B2(new_n651_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1325gat));
  OAI21_X1  g453(.A(G15gat), .B1(new_n639_), .B2(new_n269_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT41), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n625_), .A2(G15gat), .A3(new_n269_), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1326gat));
  NAND2_X1  g457(.A1(new_n455_), .A2(new_n456_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G22gat), .B1(new_n639_), .B2(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT42), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n659_), .A2(G22gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n661_), .B1(new_n625_), .B2(new_n662_), .ZN(G1327gat));
  INV_X1    g462(.A(new_n634_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n462_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n624_), .A2(new_n492_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(G29gat), .B1(new_n669_), .B2(new_n429_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n565_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n460_), .B1(new_n457_), .B2(KEYINPUT97), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n659_), .A2(new_n449_), .A3(KEYINPUT97), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n269_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n269_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n675_), .A2(new_n659_), .A3(new_n459_), .A4(new_n428_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n671_), .B1(new_n674_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT101), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT43), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n680_));
  OAI211_X1 g479(.A(KEYINPUT101), .B(new_n680_), .C1(new_n462_), .C2(new_n671_), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n679_), .A2(new_n681_), .A3(KEYINPUT44), .A4(new_n667_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n682_), .A2(G29gat), .A3(new_n429_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n679_), .A2(new_n667_), .A3(new_n681_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n670_), .B1(new_n683_), .B2(new_n686_), .ZN(G1328gat));
  INV_X1    g486(.A(KEYINPUT46), .ZN(new_n688_));
  XOR2_X1   g487(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n459_), .A2(G36gat), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n690_), .B1(new_n668_), .B2(new_n692_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n665_), .A2(new_n667_), .A3(new_n691_), .A4(new_n689_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n686_), .A2(new_n395_), .A3(new_n682_), .ZN(new_n696_));
  AOI211_X1 g495(.A(KEYINPUT103), .B(new_n695_), .C1(new_n696_), .C2(G36gat), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT103), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n684_), .A2(new_n685_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n682_), .A2(new_n395_), .ZN(new_n700_));
  OAI21_X1  g499(.A(G36gat), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n695_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n698_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n688_), .B1(new_n697_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(G36gat), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n682_), .A2(new_n395_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n706_), .B2(new_n686_), .ZN(new_n707_));
  OAI21_X1  g506(.A(KEYINPUT103), .B1(new_n707_), .B2(new_n695_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n701_), .A2(new_n698_), .A3(new_n702_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(KEYINPUT46), .A3(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n704_), .A2(new_n710_), .ZN(G1329gat));
  NAND3_X1  g510(.A1(new_n682_), .A2(G43gat), .A3(new_n675_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n668_), .A2(new_n269_), .ZN(new_n713_));
  OAI22_X1  g512(.A1(new_n699_), .A2(new_n712_), .B1(G43gat), .B2(new_n713_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g514(.A1(new_n682_), .A2(G50gat), .A3(new_n346_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n668_), .A2(new_n659_), .ZN(new_n717_));
  OAI22_X1  g516(.A1(new_n699_), .A2(new_n716_), .B1(G50gat), .B2(new_n717_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT104), .ZN(G1331gat));
  NOR2_X1   g518(.A1(new_n492_), .A2(new_n622_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n635_), .A2(new_n602_), .A3(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(G57gat), .B1(new_n721_), .B2(new_n428_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n566_), .A2(new_n623_), .A3(new_n602_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT105), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n429_), .A2(new_n416_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n722_), .B1(new_n724_), .B2(new_n725_), .ZN(G1332gat));
  OAI21_X1  g525(.A(G64gat), .B1(new_n721_), .B2(new_n459_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT48), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n459_), .A2(G64gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n724_), .B2(new_n729_), .ZN(G1333gat));
  OAI21_X1  g529(.A(G71gat), .B1(new_n721_), .B2(new_n269_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT49), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n269_), .A2(G71gat), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT106), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n732_), .B1(new_n724_), .B2(new_n734_), .ZN(G1334gat));
  OAI21_X1  g534(.A(G78gat), .B1(new_n721_), .B2(new_n659_), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n736_), .A2(KEYINPUT50), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n736_), .A2(KEYINPUT50), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n346_), .A2(new_n328_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT107), .ZN(new_n741_));
  OAI22_X1  g540(.A1(new_n738_), .A2(new_n739_), .B1(new_n724_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  OAI221_X1 g543(.A(KEYINPUT108), .B1(new_n724_), .B2(new_n741_), .C1(new_n738_), .C2(new_n739_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1335gat));
  OR2_X1    g545(.A1(new_n598_), .A2(new_n601_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n747_), .A2(new_n622_), .A3(new_n636_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n679_), .A2(new_n681_), .A3(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(G85gat), .B1(new_n749_), .B2(new_n428_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n665_), .A2(new_n748_), .ZN(new_n751_));
  INV_X1    g550(.A(G85gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(new_n752_), .A3(new_n429_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n750_), .A2(new_n753_), .ZN(G1336gat));
  OAI21_X1  g553(.A(G92gat), .B1(new_n749_), .B2(new_n459_), .ZN(new_n755_));
  INV_X1    g554(.A(G92gat), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n751_), .A2(new_n756_), .A3(new_n395_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1337gat));
  OAI21_X1  g557(.A(G99gat), .B1(new_n749_), .B2(new_n269_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n751_), .A2(new_n526_), .A3(new_n675_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g561(.A1(new_n679_), .A2(new_n681_), .A3(new_n346_), .A4(new_n748_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(G106gat), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT109), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n766_), .A2(KEYINPUT52), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n763_), .A2(KEYINPUT109), .A3(G106gat), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n766_), .A2(KEYINPUT52), .A3(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n751_), .A2(new_n338_), .A3(new_n346_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n767_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT53), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n767_), .A2(new_n773_), .A3(new_n769_), .A4(new_n770_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(G1339gat));
  NAND2_X1  g574(.A1(new_n610_), .A2(new_n606_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n604_), .A2(new_n605_), .A3(new_n611_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(new_n619_), .A3(new_n777_), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n591_), .A2(new_n621_), .A3(new_n778_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n586_), .A2(new_n587_), .A3(KEYINPUT55), .A4(new_n588_), .ZN(new_n780_));
  XOR2_X1   g579(.A(KEYINPUT111), .B(KEYINPUT55), .Z(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n581_), .B2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n586_), .A2(new_n578_), .A3(new_n588_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n579_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  OAI211_X1 g584(.A(KEYINPUT56), .B(new_n571_), .C1(new_n782_), .C2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n783_), .A2(new_n784_), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n788_), .B(new_n780_), .C1(new_n581_), .C2(new_n781_), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT56), .B1(new_n789_), .B2(new_n571_), .ZN(new_n790_));
  OAI211_X1 g589(.A(KEYINPUT58), .B(new_n779_), .C1(new_n787_), .C2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n565_), .ZN(new_n792_));
  XOR2_X1   g591(.A(KEYINPUT114), .B(KEYINPUT58), .Z(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n571_), .B1(new_n782_), .B2(new_n785_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT56), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n786_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n794_), .B1(new_n798_), .B2(new_n779_), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT115), .B1(new_n792_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n801_));
  XNOR2_X1  g600(.A(KEYINPUT112), .B(KEYINPUT57), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n621_), .A2(new_n778_), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n592_), .A2(new_n804_), .A3(new_n594_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n622_), .A2(new_n591_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n805_), .B1(new_n798_), .B2(new_n807_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n801_), .B(new_n803_), .C1(new_n808_), .C2(new_n634_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n779_), .B1(new_n787_), .B2(new_n790_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n793_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n565_), .A4(new_n791_), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n800_), .A2(new_n809_), .A3(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n803_), .B1(new_n808_), .B2(new_n634_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n808_), .A2(new_n634_), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n815_), .A2(KEYINPUT113), .B1(new_n816_), .B2(KEYINPUT57), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n636_), .B1(new_n814_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT110), .ZN(new_n820_));
  INV_X1    g619(.A(new_n720_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n820_), .B1(new_n602_), .B2(new_n821_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n720_), .B(KEYINPUT110), .C1(new_n598_), .C2(new_n601_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n819_), .B1(new_n824_), .B2(new_n671_), .ZN(new_n825_));
  AOI211_X1 g624(.A(KEYINPUT54), .B(new_n565_), .C1(new_n822_), .C2(new_n823_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT116), .B1(new_n818_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n824_), .A2(new_n671_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT54), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n824_), .A2(new_n819_), .A3(new_n671_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n815_), .A2(KEYINPUT113), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n816_), .A2(KEYINPUT57), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n800_), .A2(new_n809_), .A3(new_n813_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n492_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT116), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n832_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  NOR4_X1   g638(.A1(new_n269_), .A2(new_n346_), .A3(new_n395_), .A4(new_n428_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n828_), .A2(new_n839_), .A3(new_n622_), .A4(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(G113gat), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(KEYINPUT117), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n841_), .A2(new_n845_), .A3(new_n842_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT59), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n840_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n834_), .A2(new_n815_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n792_), .A2(new_n799_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n492_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n848_), .B1(new_n832_), .B2(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n828_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(KEYINPUT59), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n623_), .A2(new_n842_), .ZN(new_n855_));
  AOI22_X1  g654(.A1(new_n844_), .A2(new_n846_), .B1(new_n854_), .B2(new_n855_), .ZN(G1340gat));
  AND2_X1   g655(.A1(new_n828_), .A2(new_n839_), .ZN(new_n857_));
  INV_X1    g656(.A(G120gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n747_), .B2(KEYINPUT60), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n858_), .A2(KEYINPUT60), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n857_), .A2(new_n840_), .A3(new_n859_), .A4(new_n860_), .ZN(new_n861_));
  AOI211_X1 g660(.A(new_n747_), .B(new_n852_), .C1(new_n853_), .C2(KEYINPUT59), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n862_), .B2(new_n858_), .ZN(G1341gat));
  INV_X1    g662(.A(G127gat), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n857_), .A2(new_n864_), .A3(new_n636_), .A4(new_n840_), .ZN(new_n865_));
  AOI211_X1 g664(.A(new_n492_), .B(new_n852_), .C1(new_n853_), .C2(KEYINPUT59), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(new_n864_), .ZN(G1342gat));
  INV_X1    g666(.A(G134gat), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n857_), .A2(new_n868_), .A3(new_n634_), .A4(new_n840_), .ZN(new_n869_));
  AOI211_X1 g668(.A(new_n671_), .B(new_n852_), .C1(new_n853_), .C2(KEYINPUT59), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n870_), .B2(new_n868_), .ZN(G1343gat));
  XNOR2_X1  g670(.A(KEYINPUT119), .B(G141gat), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(KEYINPUT120), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n269_), .A2(new_n346_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n875_), .A2(new_n395_), .A3(new_n428_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(KEYINPUT118), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n857_), .A2(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n874_), .B1(new_n878_), .B2(new_n623_), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n857_), .A2(new_n622_), .A3(new_n877_), .A4(new_n873_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1344gat));
  OAI21_X1  g680(.A(G148gat), .B1(new_n878_), .B2(new_n747_), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n857_), .A2(new_n272_), .A3(new_n602_), .A4(new_n877_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1345gat));
  NAND4_X1  g683(.A1(new_n828_), .A2(new_n839_), .A3(new_n636_), .A4(new_n877_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT61), .B(G155gat), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(KEYINPUT121), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n885_), .B(new_n887_), .ZN(G1346gat));
  OAI21_X1  g687(.A(G162gat), .B1(new_n878_), .B2(new_n671_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n664_), .A2(G162gat), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n857_), .A2(new_n877_), .A3(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n891_), .ZN(G1347gat));
  NAND2_X1  g691(.A1(new_n832_), .A2(new_n851_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n675_), .A2(new_n395_), .A3(new_n428_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(KEYINPUT122), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n895_), .A2(new_n346_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n893_), .A2(new_n622_), .A3(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT123), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n220_), .B1(new_n898_), .B2(KEYINPUT62), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n898_), .A2(KEYINPUT62), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n893_), .A2(new_n896_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n623_), .ZN(new_n903_));
  AOI22_X1  g702(.A1(new_n900_), .A2(new_n901_), .B1(new_n903_), .B2(new_n234_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n904_), .B1(new_n900_), .B2(new_n901_), .ZN(G1348gat));
  OAI21_X1  g704(.A(new_n221_), .B1(new_n902_), .B2(new_n747_), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n895_), .A2(new_n221_), .A3(new_n747_), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n828_), .A2(new_n839_), .A3(new_n659_), .A4(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT124), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n906_), .A2(new_n908_), .A3(KEYINPUT124), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1349gat));
  INV_X1    g712(.A(new_n354_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n902_), .A2(new_n914_), .A3(new_n492_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n895_), .A2(new_n492_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n857_), .A2(new_n659_), .A3(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n232_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n915_), .B1(new_n917_), .B2(new_n918_), .ZN(G1350gat));
  OAI21_X1  g718(.A(G190gat), .B1(new_n902_), .B2(new_n671_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n634_), .A2(new_n212_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n902_), .B2(new_n921_), .ZN(G1351gat));
  NOR3_X1   g721(.A1(new_n875_), .A2(new_n459_), .A3(new_n429_), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n828_), .A2(new_n839_), .A3(new_n622_), .A4(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n924_), .A2(new_n925_), .A3(new_n307_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n924_), .B2(new_n307_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n924_), .A2(new_n307_), .ZN(new_n928_));
  NOR3_X1   g727(.A1(new_n926_), .A2(new_n927_), .A3(new_n928_), .ZN(G1352gat));
  NAND4_X1  g728(.A1(new_n828_), .A2(new_n839_), .A3(new_n602_), .A4(new_n923_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(G204gat), .ZN(G1353gat));
  NAND4_X1  g730(.A1(new_n828_), .A2(new_n839_), .A3(new_n636_), .A4(new_n923_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n933_));
  AND2_X1   g732(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n932_), .A2(new_n933_), .A3(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n932_), .A2(new_n933_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT126), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n932_), .A2(KEYINPUT126), .A3(new_n933_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n935_), .B1(new_n938_), .B2(new_n939_), .ZN(G1354gat));
  NAND4_X1  g739(.A1(new_n857_), .A2(new_n300_), .A3(new_n634_), .A4(new_n923_), .ZN(new_n941_));
  AND3_X1   g740(.A1(new_n857_), .A2(new_n565_), .A3(new_n923_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n941_), .B1(new_n942_), .B2(new_n300_), .ZN(G1355gat));
endmodule


