//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 1 0 0 0 1 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n820_,
    new_n821_, new_n822_, new_n824_, new_n825_, new_n827_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n845_, new_n846_, new_n848_, new_n849_, new_n851_, new_n852_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G211gat), .B(G218gat), .ZN(new_n207_));
  INV_X1    g006(.A(G197gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G204gat), .ZN(new_n209_));
  INV_X1    g008(.A(G204gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G197gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n207_), .B1(new_n212_), .B2(KEYINPUT21), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT92), .ZN(new_n214_));
  AND3_X1   g013(.A1(new_n209_), .A2(new_n211_), .A3(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT21), .B1(new_n209_), .B2(new_n214_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT93), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT21), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n210_), .A2(G197gat), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n218_), .B1(new_n219_), .B2(KEYINPUT92), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT93), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n209_), .A2(new_n211_), .A3(new_n214_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n213_), .B1(new_n217_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n212_), .ZN(new_n225_));
  NOR3_X1   g024(.A1(new_n225_), .A2(new_n207_), .A3(new_n218_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT94), .B1(new_n224_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n213_), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n221_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n228_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT94), .ZN(new_n232_));
  INV_X1    g031(.A(new_n226_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n235_));
  XOR2_X1   g034(.A(KEYINPUT84), .B(G190gat), .Z(new_n236_));
  AOI21_X1  g035(.A(new_n235_), .B1(new_n236_), .B2(KEYINPUT26), .ZN(new_n237_));
  XOR2_X1   g036(.A(KEYINPUT25), .B(G183gat), .Z(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT23), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT85), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT23), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n244_), .A2(G183gat), .A3(G190gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n240_), .A2(KEYINPUT85), .A3(KEYINPUT23), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n243_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  NOR3_X1   g046(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G169gat), .A2(G176gat), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n248_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n247_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT87), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n245_), .A2(new_n254_), .ZN(new_n255_));
  AOI22_X1  g054(.A1(new_n245_), .A2(new_n254_), .B1(KEYINPUT23), .B2(new_n240_), .ZN(new_n256_));
  INV_X1    g055(.A(G183gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT84), .B(G190gat), .ZN(new_n258_));
  AOI22_X1  g057(.A1(new_n255_), .A2(new_n256_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(G169gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT22), .B1(new_n260_), .B2(KEYINPUT86), .ZN(new_n261_));
  INV_X1    g060(.A(G176gat), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT22), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(G169gat), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n261_), .B(new_n262_), .C1(KEYINPUT86), .C2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(new_n251_), .ZN(new_n266_));
  OAI22_X1  g065(.A1(new_n239_), .A2(new_n253_), .B1(new_n259_), .B2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n227_), .A2(new_n234_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT97), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT97), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n227_), .A2(new_n234_), .A3(new_n270_), .A4(new_n267_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n255_), .A2(new_n256_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT26), .B(G190gat), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n273_), .B(new_n252_), .C1(new_n238_), .C2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT96), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n260_), .A2(KEYINPUT22), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n264_), .A2(new_n278_), .A3(new_n262_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n251_), .ZN(new_n280_));
  INV_X1    g079(.A(G190gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n257_), .A2(new_n281_), .ZN(new_n282_));
  AOI211_X1 g081(.A(new_n277_), .B(new_n280_), .C1(new_n247_), .C2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n247_), .A2(new_n282_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n280_), .ZN(new_n285_));
  AOI21_X1  g084(.A(KEYINPUT96), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n276_), .B1(new_n283_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n231_), .A2(new_n233_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G226gat), .A2(G233gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT20), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n289_), .A2(new_n293_), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n272_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT20), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n296_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n267_), .ZN(new_n298_));
  NOR3_X1   g097(.A1(new_n224_), .A2(KEYINPUT94), .A3(new_n226_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n232_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n298_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n292_), .B1(new_n297_), .B2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n206_), .B1(new_n295_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n297_), .A2(new_n301_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n292_), .ZN(new_n305_));
  AOI22_X1  g104(.A1(new_n272_), .A2(new_n294_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(new_n205_), .ZN(new_n307_));
  AOI21_X1  g106(.A(KEYINPUT27), .B1(new_n303_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT27), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n309_), .B1(new_n306_), .B2(new_n205_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n297_), .A2(new_n301_), .A3(new_n292_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n284_), .A2(new_n285_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n276_), .A2(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n224_), .A2(new_n226_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(KEYINPUT98), .B(KEYINPUT20), .Z(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n318_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n311_), .B1(new_n319_), .B2(new_n292_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(new_n206_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n310_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT100), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT100), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n310_), .A2(new_n324_), .A3(new_n321_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n308_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G225gat), .A2(G233gat), .ZN(new_n327_));
  NOR2_X1   g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G155gat), .A2(G162gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NOR3_X1   g130(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT89), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT2), .ZN(new_n334_));
  INV_X1    g133(.A(G141gat), .ZN(new_n335_));
  INV_X1    g134(.A(G148gat), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n334_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n331_), .B1(new_n333_), .B2(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(G141gat), .A2(G148gat), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n335_), .A2(new_n336_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n328_), .B1(KEYINPUT1), .B2(new_n330_), .ZN(new_n344_));
  OR2_X1    g143(.A1(new_n330_), .A2(KEYINPUT1), .ZN(new_n345_));
  AOI211_X1 g144(.A(new_n342_), .B(new_n343_), .C1(new_n344_), .C2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n341_), .A2(new_n346_), .ZN(new_n347_));
  XOR2_X1   g146(.A(G127gat), .B(G134gat), .Z(new_n348_));
  XOR2_X1   g147(.A(G113gat), .B(G120gat), .Z(new_n349_));
  XOR2_X1   g148(.A(new_n348_), .B(new_n349_), .Z(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n347_), .A2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n350_), .B1(new_n341_), .B2(new_n346_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n352_), .A2(KEYINPUT4), .A3(new_n353_), .ZN(new_n354_));
  OR2_X1    g153(.A1(new_n353_), .A2(KEYINPUT4), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n327_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n352_), .A2(new_n353_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n327_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G1gat), .B(G29gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(G85gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT0), .B(G57gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  OR3_X1    g163(.A1(new_n356_), .A2(new_n359_), .A3(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n364_), .B1(new_n356_), .B2(new_n359_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n288_), .B1(new_n347_), .B2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n369_), .A2(G228gat), .A3(G233gat), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT91), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n371_), .B1(new_n347_), .B2(new_n368_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G228gat), .A2(G233gat), .ZN(new_n373_));
  OAI211_X1 g172(.A(KEYINPUT91), .B(KEYINPUT29), .C1(new_n341_), .C2(new_n346_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n372_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n227_), .A2(new_n234_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n370_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  XOR2_X1   g176(.A(G22gat), .B(G50gat), .Z(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n378_), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n370_), .B(new_n380_), .C1(new_n375_), .C2(new_n376_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n347_), .A2(new_n368_), .ZN(new_n383_));
  XOR2_X1   g182(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G78gat), .B(G106gat), .ZN(new_n386_));
  INV_X1    g185(.A(new_n384_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n347_), .A2(new_n368_), .A3(new_n387_), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n385_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n386_), .B1(new_n385_), .B2(new_n388_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n382_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n379_), .A2(new_n391_), .A3(new_n381_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n367_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n320_), .A2(KEYINPUT99), .A3(KEYINPUT32), .A4(new_n205_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n397_));
  INV_X1    g196(.A(new_n318_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n272_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n305_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n397_), .B1(new_n400_), .B2(new_n311_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT99), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n402_), .B1(new_n306_), .B2(new_n397_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n396_), .B(new_n367_), .C1(new_n401_), .C2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n357_), .A2(new_n358_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n363_), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n354_), .A2(new_n355_), .A3(new_n327_), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT33), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n366_), .ZN(new_n409_));
  OAI211_X1 g208(.A(KEYINPUT33), .B(new_n364_), .C1(new_n356_), .C2(new_n359_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n409_), .A2(new_n303_), .A3(new_n307_), .A4(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n404_), .A2(new_n411_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n393_), .A2(new_n394_), .ZN(new_n413_));
  AOI22_X1  g212(.A1(new_n326_), .A2(new_n395_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G71gat), .B(G99gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(G43gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G227gat), .A2(G233gat), .ZN(new_n417_));
  INV_X1    g216(.A(G15gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n416_), .B(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT30), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n267_), .B(new_n421_), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n422_), .A2(KEYINPUT88), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(KEYINPUT88), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n420_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n424_), .A2(new_n420_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n350_), .B(KEYINPUT31), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  OR3_X1    g227(.A1(new_n425_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n428_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n303_), .A2(new_n307_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n309_), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n310_), .A2(new_n324_), .A3(new_n321_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n324_), .B1(new_n310_), .B2(new_n321_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n413_), .B(new_n433_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n367_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n431_), .A2(new_n437_), .ZN(new_n438_));
  OAI22_X1  g237(.A1(new_n414_), .A2(new_n431_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT78), .B(G15gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(G22gat), .ZN(new_n441_));
  INV_X1    g240(.A(G1gat), .ZN(new_n442_));
  INV_X1    g241(.A(G8gat), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT14), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n441_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT79), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  XOR2_X1   g246(.A(G1gat), .B(G8gat), .Z(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n445_), .B(KEYINPUT79), .ZN(new_n450_));
  INV_X1    g249(.A(new_n448_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n449_), .A2(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(G29gat), .B(G36gat), .Z(new_n454_));
  XOR2_X1   g253(.A(G43gat), .B(G50gat), .Z(new_n455_));
  XOR2_X1   g254(.A(new_n454_), .B(new_n455_), .Z(new_n456_));
  XOR2_X1   g255(.A(new_n456_), .B(KEYINPUT15), .Z(new_n457_));
  NAND2_X1  g256(.A1(new_n453_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT83), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G229gat), .A2(G233gat), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n453_), .A2(new_n456_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n460_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT82), .ZN(new_n465_));
  INV_X1    g264(.A(new_n456_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n466_), .B1(new_n449_), .B2(new_n452_), .ZN(new_n467_));
  OR3_X1    g266(.A1(new_n462_), .A2(new_n465_), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n461_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n465_), .B1(new_n462_), .B2(new_n467_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n468_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G113gat), .B(G141gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G169gat), .B(G197gat), .ZN(new_n473_));
  XOR2_X1   g272(.A(new_n472_), .B(new_n473_), .Z(new_n474_));
  AND3_X1   g273(.A1(new_n464_), .A2(new_n471_), .A3(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n474_), .B1(new_n464_), .B2(new_n471_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n439_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT101), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G230gat), .A2(G233gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT64), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT8), .ZN(new_n485_));
  NOR2_X1   g284(.A1(G99gat), .A2(G106gat), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT7), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(KEYINPUT66), .B(KEYINPUT6), .Z(new_n489_));
  NAND2_X1  g288(.A1(G99gat), .A2(G106gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT66), .B(KEYINPUT6), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n492_), .A2(G99gat), .A3(G106gat), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n488_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G85gat), .B(G92gat), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n485_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n495_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n492_), .B(new_n490_), .ZN(new_n498_));
  OAI211_X1 g297(.A(KEYINPUT8), .B(new_n497_), .C1(new_n498_), .C2(new_n488_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n495_), .A2(KEYINPUT65), .ZN(new_n500_));
  INV_X1    g299(.A(G106gat), .ZN(new_n501_));
  XOR2_X1   g300(.A(KEYINPUT10), .B(G99gat), .Z(new_n502_));
  AOI22_X1  g301(.A1(new_n500_), .A2(KEYINPUT9), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n491_), .A2(new_n493_), .ZN(new_n504_));
  INV_X1    g303(.A(G85gat), .ZN(new_n505_));
  INV_X1    g304(.A(G92gat), .ZN(new_n506_));
  AOI21_X1  g305(.A(KEYINPUT9), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n507_), .B1(new_n495_), .B2(KEYINPUT65), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n503_), .A2(new_n504_), .A3(new_n508_), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n496_), .A2(new_n499_), .A3(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G57gat), .B(G64gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT11), .ZN(new_n512_));
  XOR2_X1   g311(.A(G71gat), .B(G78gat), .Z(new_n513_));
  OR2_X1    g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n511_), .A2(KEYINPUT11), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n512_), .A2(new_n513_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n514_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n510_), .A2(new_n517_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n496_), .A2(new_n499_), .A3(new_n509_), .A4(new_n517_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n484_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT67), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n496_), .A2(new_n499_), .A3(new_n509_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT68), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT12), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n517_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT68), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n496_), .A2(new_n499_), .A3(new_n528_), .A4(new_n509_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n524_), .A2(new_n527_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT69), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n519_), .A2(new_n483_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT70), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT70), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n519_), .A2(new_n535_), .A3(new_n483_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n525_), .B1(new_n510_), .B2(new_n517_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n524_), .A2(new_n527_), .A3(KEYINPUT69), .A4(new_n529_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n532_), .A2(new_n537_), .A3(new_n538_), .A4(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n522_), .A2(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(G120gat), .B(G148gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G176gat), .B(G204gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n541_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n546_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n522_), .A2(new_n540_), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n550_), .B1(KEYINPUT72), .B2(KEYINPUT13), .ZN(new_n551_));
  XOR2_X1   g350(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n552_));
  OAI21_X1  g351(.A(new_n551_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n523_), .A2(new_n456_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT75), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n457_), .A2(new_n524_), .A3(new_n529_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G232gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT74), .B(KEYINPUT35), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n555_), .A2(new_n556_), .A3(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n560_), .A2(new_n561_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n564_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n555_), .A2(new_n556_), .A3(new_n566_), .A4(new_n562_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G190gat), .B(G218gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT76), .ZN(new_n570_));
  XOR2_X1   g369(.A(G134gat), .B(G162gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n572_), .B(KEYINPUT36), .Z(new_n573_));
  NAND2_X1  g372(.A1(new_n568_), .A2(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n572_), .A2(KEYINPUT36), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n565_), .A2(new_n575_), .A3(new_n567_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n574_), .A2(KEYINPUT37), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n576_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n573_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n579_), .B1(new_n568_), .B2(KEYINPUT77), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT77), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n565_), .A2(new_n581_), .A3(new_n567_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n578_), .B1(new_n580_), .B2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n577_), .B1(new_n583_), .B2(KEYINPUT37), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n453_), .B(KEYINPUT80), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G231gat), .A2(G233gat), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n586_), .B(KEYINPUT81), .Z(new_n587_));
  XOR2_X1   g386(.A(new_n517_), .B(new_n587_), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n585_), .B(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G127gat), .B(G155gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT16), .ZN(new_n591_));
  XOR2_X1   g390(.A(G183gat), .B(G211gat), .Z(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT17), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n589_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT17), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n589_), .B1(new_n596_), .B2(new_n593_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n584_), .A2(new_n599_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n481_), .A2(new_n553_), .A3(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n367_), .B(KEYINPUT102), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(new_n442_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT38), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n583_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n439_), .A2(new_n606_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n607_), .A2(new_n478_), .A3(new_n553_), .A4(new_n598_), .ZN(new_n608_));
  OAI21_X1  g407(.A(G1gat), .B1(new_n608_), .B2(new_n437_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n603_), .A2(new_n604_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n605_), .A2(new_n609_), .A3(new_n610_), .ZN(G1324gat));
  OAI21_X1  g410(.A(G8gat), .B1(new_n608_), .B2(new_n326_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT39), .ZN(new_n613_));
  INV_X1    g412(.A(new_n326_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n601_), .A2(new_n443_), .A3(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g416(.A(new_n431_), .ZN(new_n618_));
  OAI21_X1  g417(.A(G15gat), .B1(new_n608_), .B2(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n619_), .B(KEYINPUT41), .Z(new_n620_));
  NAND3_X1  g419(.A1(new_n601_), .A2(new_n418_), .A3(new_n431_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(G1326gat));
  OAI21_X1  g421(.A(G22gat), .B1(new_n608_), .B2(new_n413_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT103), .Z(new_n624_));
  OR2_X1    g423(.A1(new_n624_), .A2(KEYINPUT42), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(KEYINPUT42), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n413_), .A2(G22gat), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT104), .Z(new_n628_));
  NAND2_X1  g427(.A1(new_n601_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n625_), .A2(new_n626_), .A3(new_n629_), .ZN(G1327gat));
  NAND2_X1  g429(.A1(new_n412_), .A2(new_n413_), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n395_), .B(new_n433_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n431_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n436_), .A2(new_n367_), .A3(new_n618_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n584_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT43), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT43), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n584_), .B(new_n637_), .C1(new_n633_), .C2(new_n634_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n636_), .A2(KEYINPUT106), .A3(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n553_), .A2(new_n478_), .A3(new_n599_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT105), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n553_), .A2(KEYINPUT105), .A3(new_n478_), .A4(new_n599_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n642_), .A2(KEYINPUT106), .A3(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n639_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT44), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT44), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n639_), .A2(new_n644_), .A3(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n649_), .A2(KEYINPUT107), .A3(new_n602_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(G29gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(KEYINPUT107), .B1(new_n649_), .B2(new_n602_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n553_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n599_), .A2(new_n583_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n481_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT108), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n481_), .A2(KEYINPUT108), .A3(new_n655_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n437_), .A2(G29gat), .ZN(new_n661_));
  OAI22_X1  g460(.A1(new_n651_), .A2(new_n652_), .B1(new_n660_), .B2(new_n661_), .ZN(G1328gat));
  NOR2_X1   g461(.A1(new_n326_), .A2(G36gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n658_), .A2(new_n659_), .A3(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n665_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n658_), .A2(new_n659_), .A3(new_n667_), .A4(new_n663_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT109), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n649_), .A2(new_n669_), .A3(new_n614_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(G36gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n669_), .B1(new_n649_), .B2(new_n614_), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n666_), .B(new_n668_), .C1(new_n671_), .C2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT46), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n649_), .A2(new_n614_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT109), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n677_), .A2(G36gat), .A3(new_n670_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n678_), .A2(KEYINPUT46), .A3(new_n666_), .A4(new_n668_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n675_), .A2(new_n679_), .ZN(G1329gat));
  INV_X1    g479(.A(new_n649_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G43gat), .B1(new_n681_), .B2(new_n618_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n618_), .A2(G43gat), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n658_), .A2(new_n659_), .A3(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT47), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n685_), .B(new_n686_), .ZN(G1330gat));
  INV_X1    g486(.A(new_n413_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n658_), .A2(new_n688_), .A3(new_n659_), .ZN(new_n689_));
  INV_X1    g488(.A(G50gat), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n413_), .A2(new_n690_), .ZN(new_n691_));
  AOI22_X1  g490(.A1(new_n689_), .A2(new_n690_), .B1(new_n649_), .B2(new_n691_), .ZN(G1331gat));
  NOR3_X1   g491(.A1(new_n553_), .A2(new_n599_), .A3(new_n478_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n607_), .A2(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G57gat), .B1(new_n694_), .B2(new_n437_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n439_), .A2(new_n477_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(new_n653_), .A3(new_n600_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n602_), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n698_), .A2(G57gat), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n695_), .B1(new_n697_), .B2(new_n699_), .ZN(G1332gat));
  OAI21_X1  g499(.A(G64gat), .B1(new_n694_), .B2(new_n326_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT48), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n326_), .A2(G64gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n697_), .B2(new_n703_), .ZN(G1333gat));
  OAI21_X1  g503(.A(G71gat), .B1(new_n694_), .B2(new_n618_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT49), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n618_), .A2(G71gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n706_), .B1(new_n697_), .B2(new_n707_), .ZN(G1334gat));
  OAI21_X1  g507(.A(G78gat), .B1(new_n694_), .B2(new_n413_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT50), .ZN(new_n710_));
  OR3_X1    g509(.A1(new_n697_), .A2(G78gat), .A3(new_n413_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT111), .Z(G1335gat));
  NAND4_X1  g512(.A1(new_n696_), .A2(new_n653_), .A3(new_n599_), .A4(new_n583_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n715_), .A2(new_n505_), .A3(new_n602_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT113), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n636_), .A2(KEYINPUT112), .A3(new_n638_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n553_), .A2(new_n478_), .A3(new_n598_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT112), .B1(new_n636_), .B2(new_n638_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n636_), .A2(new_n638_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT112), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n725_), .A2(KEYINPUT113), .A3(new_n719_), .A4(new_n718_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n722_), .A2(new_n367_), .A3(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n716_), .B1(new_n727_), .B2(new_n505_), .ZN(G1336gat));
  NAND3_X1  g527(.A1(new_n715_), .A2(new_n506_), .A3(new_n614_), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n722_), .A2(new_n614_), .A3(new_n726_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n730_), .B2(new_n506_), .ZN(G1337gat));
  NAND3_X1  g530(.A1(new_n715_), .A2(new_n431_), .A3(new_n502_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n722_), .A2(new_n431_), .A3(new_n726_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT114), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n733_), .A2(new_n734_), .A3(G99gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n733_), .B2(G99gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n732_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT51), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n738_), .A2(KEYINPUT115), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(new_n740_));
  OAI221_X1 g539(.A(new_n732_), .B1(KEYINPUT115), .B2(new_n738_), .C1(new_n735_), .C2(new_n736_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1338gat));
  AND2_X1   g541(.A1(new_n719_), .A2(new_n688_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n501_), .B1(new_n723_), .B2(new_n743_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT52), .Z(new_n745_));
  NAND3_X1  g544(.A1(new_n715_), .A2(new_n501_), .A3(new_n688_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n747_), .B(new_n748_), .ZN(G1339gat));
  NAND3_X1  g548(.A1(new_n600_), .A2(new_n477_), .A3(new_n553_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT54), .Z(new_n751_));
  NAND3_X1  g550(.A1(new_n464_), .A2(new_n471_), .A3(new_n474_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n460_), .A2(new_n469_), .A3(new_n463_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n468_), .A2(new_n461_), .A3(new_n470_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n474_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n753_), .A2(new_n754_), .A3(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n550_), .A2(new_n752_), .A3(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n549_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT119), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT55), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(new_n540_), .B2(new_n760_), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n532_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n762_), .A2(KEYINPUT119), .A3(KEYINPUT55), .A4(new_n537_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT117), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n540_), .A2(new_n764_), .A3(new_n760_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n540_), .B2(new_n760_), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n761_), .B(new_n763_), .C1(new_n765_), .C2(new_n766_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n532_), .A2(new_n538_), .A3(new_n539_), .A4(new_n519_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n484_), .B1(new_n768_), .B2(KEYINPUT118), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n769_), .B1(KEYINPUT118), .B2(new_n768_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n546_), .B1(new_n767_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT56), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  OAI211_X1 g572(.A(KEYINPUT56), .B(new_n546_), .C1(new_n767_), .C2(new_n770_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n758_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n757_), .B1(new_n775_), .B2(KEYINPUT120), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT120), .ZN(new_n777_));
  AOI211_X1 g576(.A(new_n777_), .B(new_n758_), .C1(new_n773_), .C2(new_n774_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n606_), .B1(new_n776_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT57), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  OAI211_X1 g580(.A(KEYINPUT57), .B(new_n606_), .C1(new_n776_), .C2(new_n778_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n752_), .A2(new_n756_), .A3(new_n549_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n584_), .B1(new_n784_), .B2(KEYINPUT58), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT121), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(KEYINPUT58), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT121), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n788_), .B(new_n584_), .C1(new_n784_), .C2(KEYINPUT58), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n786_), .A2(new_n787_), .A3(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n781_), .A2(new_n782_), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n751_), .B1(new_n791_), .B2(new_n599_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n436_), .A2(new_n698_), .A3(new_n618_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  OAI22_X1  g593(.A1(new_n792_), .A2(new_n794_), .B1(KEYINPUT122), .B2(KEYINPUT59), .ZN(new_n795_));
  XNOR2_X1  g594(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n789_), .A2(new_n787_), .ZN(new_n797_));
  AOI22_X1  g596(.A1(new_n797_), .A2(new_n786_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n598_), .B1(new_n798_), .B2(new_n782_), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n793_), .B(new_n796_), .C1(new_n799_), .C2(new_n751_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n795_), .A2(new_n800_), .A3(new_n478_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(G113gat), .ZN(new_n802_));
  OR4_X1    g601(.A1(G113gat), .A2(new_n792_), .A3(new_n477_), .A4(new_n794_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(G1340gat));
  NAND3_X1  g603(.A1(new_n795_), .A2(new_n800_), .A3(new_n653_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(G120gat), .ZN(new_n806_));
  INV_X1    g605(.A(new_n792_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n553_), .A2(KEYINPUT60), .ZN(new_n808_));
  MUX2_X1   g607(.A(new_n808_), .B(KEYINPUT60), .S(G120gat), .Z(new_n809_));
  NAND3_X1  g608(.A1(new_n807_), .A2(new_n793_), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n806_), .A2(new_n810_), .ZN(G1341gat));
  NAND4_X1  g610(.A1(new_n795_), .A2(new_n800_), .A3(G127gat), .A4(new_n598_), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n792_), .A2(new_n599_), .A3(new_n794_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT123), .B1(new_n813_), .B2(G127gat), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n598_), .B(new_n793_), .C1(new_n799_), .C2(new_n751_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT123), .ZN(new_n816_));
  INV_X1    g615(.A(G127gat), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n815_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n812_), .A2(new_n814_), .A3(new_n818_), .ZN(G1342gat));
  NAND3_X1  g618(.A1(new_n795_), .A2(new_n800_), .A3(new_n584_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(G134gat), .ZN(new_n821_));
  OR4_X1    g620(.A1(G134gat), .A2(new_n792_), .A3(new_n606_), .A4(new_n794_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(G1343gat));
  NOR4_X1   g622(.A1(new_n614_), .A2(new_n698_), .A3(new_n413_), .A4(new_n431_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n807_), .A2(new_n478_), .A3(new_n824_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g625(.A1(new_n807_), .A2(new_n653_), .A3(new_n824_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g627(.A1(new_n807_), .A2(new_n598_), .A3(new_n824_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(KEYINPUT61), .B(G155gat), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n829_), .B(new_n830_), .ZN(G1346gat));
  AND3_X1   g630(.A1(new_n807_), .A2(new_n584_), .A3(new_n824_), .ZN(new_n832_));
  INV_X1    g631(.A(G162gat), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n807_), .A2(new_n824_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n583_), .A2(new_n833_), .ZN(new_n835_));
  OAI22_X1  g634(.A1(new_n832_), .A2(new_n833_), .B1(new_n834_), .B2(new_n835_), .ZN(G1347gat));
  NOR4_X1   g635(.A1(new_n326_), .A2(new_n618_), .A3(new_n602_), .A4(new_n688_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n792_), .A2(new_n477_), .A3(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT62), .ZN(new_n840_));
  OR3_X1    g639(.A1(new_n839_), .A2(new_n840_), .A3(new_n260_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n839_), .B2(new_n260_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n839_), .A2(new_n264_), .A3(new_n278_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n841_), .A2(new_n842_), .A3(new_n843_), .ZN(G1348gat));
  NOR2_X1   g643(.A1(new_n792_), .A2(new_n838_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n653_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(G176gat), .ZN(G1349gat));
  AOI21_X1  g646(.A(G183gat), .B1(new_n845_), .B2(new_n598_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n792_), .A2(new_n599_), .A3(new_n838_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n848_), .B1(new_n238_), .B2(new_n849_), .ZN(G1350gat));
  NAND3_X1  g649(.A1(new_n845_), .A2(new_n274_), .A3(new_n583_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n845_), .A2(new_n584_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n852_), .B2(new_n281_), .ZN(G1351gat));
  NAND3_X1  g652(.A1(new_n614_), .A2(new_n395_), .A3(new_n618_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n792_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n478_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g656(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n858_), .B1(new_n855_), .B2(new_n653_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n860_));
  XOR2_X1   g659(.A(new_n860_), .B(KEYINPUT125), .Z(new_n861_));
  NOR2_X1   g660(.A1(new_n859_), .A2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n861_), .ZN(new_n863_));
  AOI211_X1 g662(.A(new_n858_), .B(new_n863_), .C1(new_n855_), .C2(new_n653_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n862_), .A2(new_n864_), .ZN(G1353gat));
  INV_X1    g664(.A(KEYINPUT63), .ZN(new_n866_));
  INV_X1    g665(.A(G211gat), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n598_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(KEYINPUT126), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT127), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n870_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n866_), .A2(new_n867_), .A3(KEYINPUT127), .ZN(new_n872_));
  AOI22_X1  g671(.A1(new_n855_), .A2(new_n869_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n855_), .A2(new_n869_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n873_), .B1(new_n874_), .B2(new_n872_), .ZN(G1354gat));
  INV_X1    g674(.A(G218gat), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n855_), .A2(new_n876_), .A3(new_n583_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n855_), .A2(new_n584_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n878_), .B2(new_n876_), .ZN(G1355gat));
endmodule


