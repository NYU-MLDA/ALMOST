//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 1 1 0 1 0 0 1 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 1 1 1 1 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n817_, new_n818_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n946_, new_n947_,
    new_n948_, new_n950_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n960_, new_n961_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n979_, new_n980_, new_n981_, new_n983_, new_n984_,
    new_n985_, new_n987_, new_n988_, new_n990_, new_n991_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n999_, new_n1000_,
    new_n1001_;
  NAND2_X1  g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT86), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT86), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G141gat), .A3(G148gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT2), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n203_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n209_));
  AND2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT3), .ZN(new_n211_));
  INV_X1    g010(.A(G141gat), .ZN(new_n212_));
  INV_X1    g011(.A(G148gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT89), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT89), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n216_), .A2(new_n211_), .A3(new_n212_), .A4(new_n213_), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n207_), .A2(new_n210_), .A3(new_n215_), .A4(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT90), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT87), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT87), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(G155gat), .A3(G162gat), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n220_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n225_));
  AND3_X1   g024(.A1(new_n218_), .A2(new_n219_), .A3(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n219_), .B1(new_n218_), .B2(new_n225_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n203_), .B(new_n205_), .C1(G141gat), .C2(G148gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n222_), .A2(new_n224_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n220_), .B1(new_n230_), .B2(KEYINPUT1), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT1), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n222_), .A2(new_n224_), .ZN(new_n233_));
  AOI22_X1  g032(.A1(new_n231_), .A2(KEYINPUT88), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT88), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n232_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n235_), .B1(new_n236_), .B2(new_n220_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n229_), .B1(new_n234_), .B2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT91), .B1(new_n228_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n218_), .A2(new_n225_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT90), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n218_), .A2(new_n219_), .A3(new_n225_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT91), .ZN(new_n244_));
  INV_X1    g043(.A(new_n220_), .ZN(new_n245_));
  OAI211_X1 g044(.A(KEYINPUT88), .B(new_n245_), .C1(new_n233_), .C2(new_n232_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n233_), .A2(new_n232_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n246_), .A2(new_n237_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n229_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n243_), .A2(new_n244_), .A3(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G127gat), .B(G134gat), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n253_), .A2(KEYINPUT84), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(KEYINPUT84), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G113gat), .B(G120gat), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n254_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n256_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n239_), .A2(new_n251_), .A3(new_n252_), .A4(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G225gat), .A2(G233gat), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n243_), .A2(new_n259_), .A3(new_n250_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT95), .ZN(new_n266_));
  AOI22_X1  g065(.A1(new_n241_), .A2(new_n242_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT95), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(new_n268_), .A3(new_n259_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n266_), .A2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n239_), .A2(new_n251_), .A3(new_n260_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n270_), .A2(KEYINPUT4), .A3(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n264_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n270_), .A2(new_n271_), .A3(new_n262_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G1gat), .B(G29gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(G85gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT0), .B(G57gat), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n276_), .B(new_n277_), .Z(new_n278_));
  NAND3_X1  g077(.A1(new_n273_), .A2(new_n274_), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT96), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n280_), .A2(KEYINPUT33), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G8gat), .B(G36gat), .Z(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT18), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G64gat), .B(G92gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G226gat), .A2(G233gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT19), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NOR3_X1   g089(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT24), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n292_), .B1(G169gat), .B2(G176gat), .ZN(new_n293_));
  NOR2_X1   g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n291_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(G190gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT26), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT26), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(G190gat), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT25), .ZN(new_n301_));
  INV_X1    g100(.A(G183gat), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n298_), .B(new_n300_), .C1(new_n303_), .C2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n296_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT83), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G183gat), .A2(G190gat), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n307_), .B1(new_n308_), .B2(KEYINPUT23), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(KEYINPUT23), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT23), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n311_), .A2(G183gat), .A3(G190gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n309_), .B1(new_n313_), .B2(new_n307_), .ZN(new_n314_));
  OR2_X1    g113(.A1(KEYINPUT82), .A2(G176gat), .ZN(new_n315_));
  INV_X1    g114(.A(G169gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT22), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT22), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(G169gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(KEYINPUT82), .A2(G176gat), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n315_), .A2(new_n317_), .A3(new_n319_), .A4(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  AOI22_X1  g122(.A1(new_n310_), .A2(new_n312_), .B1(new_n302_), .B2(new_n297_), .ZN(new_n324_));
  OAI22_X1  g123(.A1(new_n306_), .A2(new_n314_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT21), .ZN(new_n326_));
  AND2_X1   g125(.A1(G197gat), .A2(G204gat), .ZN(new_n327_));
  NOR2_X1   g126(.A1(G197gat), .A2(G204gat), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n326_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(G197gat), .ZN(new_n330_));
  INV_X1    g129(.A(G204gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G197gat), .A2(G204gat), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(KEYINPUT21), .A3(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G211gat), .B(G218gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n329_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(G218gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(G211gat), .ZN(new_n338_));
  INV_X1    g137(.A(G211gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(G218gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n341_), .A2(KEYINPUT21), .A3(new_n332_), .A4(new_n333_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n336_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n325_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT94), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT94), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n325_), .A2(new_n346_), .A3(new_n343_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT20), .ZN(new_n349_));
  AND2_X1   g148(.A1(new_n321_), .A2(new_n322_), .ZN(new_n350_));
  AOI21_X1  g149(.A(KEYINPUT83), .B1(new_n310_), .B2(new_n312_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT81), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(new_n302_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(KEYINPUT81), .A2(G183gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  OAI22_X1  g154(.A1(new_n351_), .A2(new_n309_), .B1(G190gat), .B2(new_n355_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n310_), .A2(new_n312_), .ZN(new_n357_));
  INV_X1    g156(.A(G176gat), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n292_), .A2(new_n316_), .A3(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n322_), .A2(KEYINPUT24), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n359_), .B1(new_n360_), .B2(new_n294_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n357_), .A2(new_n361_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n298_), .A2(new_n300_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n301_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n363_), .B1(new_n364_), .B2(new_n304_), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n350_), .A2(new_n356_), .B1(new_n362_), .B2(new_n365_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n336_), .A2(new_n342_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n349_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n290_), .B1(new_n348_), .B2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT20), .B1(new_n366_), .B2(new_n367_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n290_), .B1(new_n325_), .B2(new_n343_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n287_), .B1(new_n369_), .B2(new_n372_), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n370_), .A2(new_n371_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n356_), .A2(new_n350_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n362_), .A2(new_n365_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(new_n367_), .A3(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT20), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n378_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n286_), .B(new_n374_), .C1(new_n379_), .C2(new_n290_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n373_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n270_), .A2(new_n271_), .A3(new_n263_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n278_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n272_), .A2(new_n262_), .A3(new_n261_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n381_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n281_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n273_), .A2(new_n274_), .A3(new_n278_), .A4(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n282_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n286_), .A2(KEYINPUT32), .ZN(new_n390_));
  NOR3_X1   g189(.A1(new_n369_), .A2(new_n390_), .A3(new_n372_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n325_), .A2(new_n346_), .A3(new_n343_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n346_), .B1(new_n325_), .B2(new_n343_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n368_), .B(new_n290_), .C1(new_n392_), .C2(new_n393_), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n336_), .A2(KEYINPUT92), .A3(new_n342_), .ZN(new_n395_));
  AOI21_X1  g194(.A(KEYINPUT92), .B1(new_n336_), .B2(new_n342_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n325_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n289_), .B1(new_n370_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n394_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n390_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT97), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n399_), .A2(KEYINPUT97), .A3(new_n390_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n391_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n273_), .A2(new_n274_), .A3(new_n278_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n278_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n404_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n389_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n239_), .A2(KEYINPUT29), .A3(new_n251_), .ZN(new_n409_));
  AND2_X1   g208(.A1(G228gat), .A2(G233gat), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n367_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT29), .ZN(new_n413_));
  OAI22_X1  g212(.A1(new_n267_), .A2(new_n413_), .B1(new_n396_), .B2(new_n395_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(new_n410_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n412_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G78gat), .B(G106gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(KEYINPUT29), .B1(new_n239_), .B2(new_n251_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G22gat), .B(G50gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT28), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n419_), .B(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT93), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n409_), .A2(new_n411_), .B1(new_n414_), .B2(new_n410_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n417_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n418_), .A2(new_n423_), .A3(new_n424_), .A4(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT93), .B1(new_n425_), .B2(new_n426_), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n430_), .A2(new_n423_), .B1(new_n418_), .B2(new_n427_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n408_), .A2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT98), .B1(new_n405_), .B2(new_n406_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n273_), .A2(new_n274_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n383_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT98), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n437_), .A3(new_n279_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n434_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n399_), .A2(new_n287_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n440_), .A2(new_n380_), .A3(KEYINPUT27), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT99), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT27), .ZN(new_n443_));
  INV_X1    g242(.A(new_n380_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n368_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(new_n289_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n286_), .B1(new_n446_), .B2(new_n374_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n443_), .B1(new_n444_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT99), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n440_), .A2(new_n380_), .A3(new_n449_), .A4(KEYINPUT27), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n442_), .A2(new_n448_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n430_), .A2(new_n423_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n418_), .A2(new_n427_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n451_), .B1(new_n454_), .B2(new_n428_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n439_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n433_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G227gat), .A2(G233gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(G15gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT30), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n366_), .B(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(new_n260_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G71gat), .B(G99gat), .ZN(new_n463_));
  INV_X1    g262(.A(G43gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT31), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n462_), .B(new_n466_), .ZN(new_n467_));
  XOR2_X1   g266(.A(new_n467_), .B(KEYINPUT85), .Z(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT100), .ZN(new_n470_));
  AND3_X1   g269(.A1(new_n442_), .A2(new_n448_), .A3(new_n450_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n432_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n454_), .A2(new_n428_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT100), .B1(new_n473_), .B2(new_n451_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n467_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n476_), .B1(new_n434_), .B2(new_n438_), .ZN(new_n477_));
  AOI22_X1  g276(.A1(new_n457_), .A2(new_n469_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n478_));
  XOR2_X1   g277(.A(G29gat), .B(G36gat), .Z(new_n479_));
  XOR2_X1   g278(.A(G43gat), .B(G50gat), .Z(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(G1gat), .ZN(new_n483_));
  INV_X1    g282(.A(G8gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT14), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT74), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT74), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n487_), .B(KEYINPUT14), .C1(new_n483_), .C2(new_n484_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G15gat), .B(G22gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n486_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT75), .ZN(new_n491_));
  XOR2_X1   g290(.A(G1gat), .B(G8gat), .Z(new_n492_));
  INV_X1    g291(.A(KEYINPUT75), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n486_), .A2(new_n493_), .A3(new_n488_), .A4(new_n489_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n491_), .A2(new_n492_), .A3(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n492_), .B1(new_n491_), .B2(new_n494_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n482_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n497_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n499_), .A2(new_n481_), .A3(new_n495_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n498_), .A2(new_n500_), .A3(KEYINPUT79), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G229gat), .A2(G233gat), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT79), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n504_), .B(new_n482_), .C1(new_n496_), .C2(new_n497_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n501_), .A2(new_n503_), .A3(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n481_), .B(KEYINPUT15), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n507_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n508_), .A2(new_n502_), .A3(new_n500_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n506_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G113gat), .B(G141gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G169gat), .B(G197gat), .ZN(new_n512_));
  XOR2_X1   g311(.A(new_n511_), .B(new_n512_), .Z(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n510_), .A2(KEYINPUT80), .A3(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(KEYINPUT80), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n506_), .A2(new_n516_), .A3(new_n509_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT70), .ZN(new_n520_));
  XOR2_X1   g319(.A(KEYINPUT10), .B(G99gat), .Z(new_n521_));
  INV_X1    g320(.A(G106gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(G85gat), .ZN(new_n524_));
  INV_X1    g323(.A(G92gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G85gat), .A2(G92gat), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n526_), .A2(KEYINPUT9), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(G99gat), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT6), .B1(new_n529_), .B2(new_n522_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT6), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n531_), .A2(G99gat), .A3(G106gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n527_), .A2(KEYINPUT9), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n523_), .A2(new_n528_), .A3(new_n533_), .A4(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT8), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NOR3_X1   g337(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT65), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT7), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n541_), .A2(new_n529_), .A3(new_n522_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT65), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n542_), .A2(new_n543_), .A3(new_n537_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n540_), .A2(new_n544_), .A3(new_n533_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT64), .ZN(new_n546_));
  INV_X1    g345(.A(new_n527_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(G85gat), .A2(G92gat), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n546_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n526_), .A2(KEYINPUT64), .A3(new_n527_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n536_), .B1(new_n545_), .B2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n549_), .A2(new_n550_), .A3(new_n536_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n542_), .A2(new_n537_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n554_), .B1(new_n556_), .B2(new_n533_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n535_), .B1(new_n553_), .B2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G57gat), .B(G64gat), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(KEYINPUT11), .ZN(new_n560_));
  XOR2_X1   g359(.A(G71gat), .B(G78gat), .Z(new_n561_));
  OR2_X1    g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n559_), .A2(KEYINPUT11), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n560_), .A2(new_n561_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n562_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n558_), .A2(new_n566_), .A3(KEYINPUT12), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n565_), .B(new_n535_), .C1(new_n553_), .C2(new_n557_), .ZN(new_n568_));
  AOI22_X1  g367(.A1(new_n555_), .A2(KEYINPUT65), .B1(new_n530_), .B2(new_n532_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n551_), .B1(new_n569_), .B2(new_n544_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n555_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n571_));
  OAI22_X1  g370(.A1(new_n570_), .A2(new_n536_), .B1(new_n571_), .B2(new_n554_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n565_), .B1(new_n572_), .B2(new_n535_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT68), .B(KEYINPUT12), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n567_), .B(new_n568_), .C1(new_n573_), .C2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G230gat), .A2(G233gat), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(KEYINPUT69), .B1(new_n575_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n568_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n558_), .A2(new_n566_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n574_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n579_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT69), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n582_), .A2(new_n583_), .A3(new_n576_), .A4(new_n567_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n578_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT66), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n558_), .A2(new_n566_), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(new_n568_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n586_), .B1(new_n558_), .B2(new_n566_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n577_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(KEYINPUT67), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT67), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n592_), .B(new_n577_), .C1(new_n588_), .C2(new_n589_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G120gat), .B(G148gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT5), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G176gat), .B(G204gat), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n596_), .B(new_n597_), .Z(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n585_), .A2(new_n594_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n599_), .B1(new_n585_), .B2(new_n594_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n520_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n591_), .A2(new_n593_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n578_), .A2(new_n584_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n598_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(KEYINPUT70), .A3(new_n600_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n603_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT13), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n603_), .A2(KEYINPUT13), .A3(new_n607_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n507_), .A2(new_n558_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n572_), .A2(new_n535_), .A3(new_n481_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G232gat), .A2(G233gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT34), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(KEYINPUT35), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n617_), .A2(KEYINPUT35), .ZN(new_n620_));
  OR3_X1    g419(.A1(new_n615_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT71), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n622_), .B1(new_n615_), .B2(new_n619_), .ZN(new_n623_));
  AOI211_X1 g422(.A(KEYINPUT71), .B(new_n618_), .C1(new_n613_), .C2(new_n614_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n621_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT73), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n623_), .A2(new_n624_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(KEYINPUT73), .A3(new_n621_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G190gat), .B(G218gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT72), .ZN(new_n631_));
  XOR2_X1   g430(.A(G134gat), .B(G162gat), .Z(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT36), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n627_), .A2(new_n629_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT36), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n633_), .A2(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n625_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(KEYINPUT37), .B1(new_n635_), .B2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(G231gat), .A2(G233gat), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n566_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n566_), .A2(new_n641_), .ZN(new_n644_));
  OAI22_X1  g443(.A1(new_n643_), .A2(new_n644_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n565_), .A2(G231gat), .A3(G233gat), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n646_), .A2(new_n495_), .A3(new_n642_), .A4(new_n499_), .ZN(new_n647_));
  XOR2_X1   g446(.A(G127gat), .B(G155gat), .Z(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT16), .ZN(new_n649_));
  XNOR2_X1  g448(.A(G183gat), .B(G211gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT17), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n651_), .A2(new_n652_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n645_), .A2(new_n647_), .A3(new_n653_), .A4(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT77), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n645_), .A2(new_n647_), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n658_), .A2(KEYINPUT76), .A3(new_n654_), .ZN(new_n659_));
  AOI21_X1  g458(.A(KEYINPUT76), .B1(new_n658_), .B2(new_n654_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(KEYINPUT78), .B1(new_n657_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT77), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n656_), .B(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT78), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n664_), .B(new_n665_), .C1(new_n660_), .C2(new_n659_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n662_), .A2(new_n666_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n625_), .A2(new_n634_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT37), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n668_), .A2(new_n638_), .A3(new_n669_), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n640_), .A2(new_n667_), .A3(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NOR4_X1   g471(.A1(new_n478_), .A2(new_n519_), .A3(new_n612_), .A4(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n439_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(new_n674_), .A3(new_n483_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT38), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(KEYINPUT102), .B2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(KEYINPUT102), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n677_), .B(new_n678_), .Z(new_n679_));
  NAND2_X1  g478(.A1(new_n635_), .A2(new_n639_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n478_), .A2(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n657_), .A2(new_n661_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n612_), .A2(new_n684_), .A3(new_n519_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n682_), .A2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT101), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n687_), .A2(new_n674_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n679_), .B1(new_n483_), .B2(new_n688_), .ZN(G1324gat));
  NAND3_X1  g488(.A1(new_n682_), .A2(new_n451_), .A3(new_n685_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(G8gat), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(KEYINPUT39), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT103), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n691_), .A2(new_n694_), .A3(KEYINPUT39), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n696_), .B1(new_n691_), .B2(KEYINPUT39), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT39), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n690_), .A2(KEYINPUT104), .A3(new_n698_), .A4(G8gat), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n693_), .A2(new_n695_), .A3(new_n697_), .A4(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n673_), .A2(new_n484_), .A3(new_n451_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT40), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n700_), .A2(KEYINPUT40), .A3(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1325gat));
  INV_X1    g505(.A(G15gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n707_), .B1(new_n687_), .B2(new_n468_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT41), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n673_), .A2(new_n707_), .A3(new_n468_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1326gat));
  INV_X1    g510(.A(G22gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n712_), .B1(new_n687_), .B2(new_n473_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT42), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n713_), .B(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n673_), .A2(new_n712_), .A3(new_n473_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1327gat));
  INV_X1    g516(.A(G29gat), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n640_), .A2(new_n670_), .ZN(new_n719_));
  OAI21_X1  g518(.A(KEYINPUT43), .B1(new_n478_), .B2(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n470_), .B1(new_n432_), .B2(new_n471_), .ZN(new_n721_));
  AND4_X1   g520(.A1(new_n470_), .A2(new_n471_), .A3(new_n428_), .A4(new_n454_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n477_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  AOI22_X1  g522(.A1(new_n432_), .A2(new_n408_), .B1(new_n439_), .B2(new_n455_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n723_), .B1(new_n724_), .B2(new_n468_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n640_), .A2(new_n670_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n725_), .A2(new_n726_), .A3(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n720_), .A2(new_n728_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n610_), .A2(new_n611_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n730_), .A2(new_n518_), .A3(new_n667_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(KEYINPUT44), .B1(new_n729_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n734_));
  AOI211_X1 g533(.A(new_n734_), .B(new_n731_), .C1(new_n720_), .C2(new_n728_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n733_), .A2(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n718_), .B1(new_n736_), .B2(new_n674_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n478_), .A2(new_n519_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n681_), .A2(new_n667_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n612_), .A2(new_n739_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n738_), .A2(new_n740_), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n741_), .A2(new_n718_), .A3(new_n674_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n737_), .A2(new_n742_), .ZN(G1328gat));
  NOR2_X1   g542(.A1(new_n471_), .A2(G36gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n738_), .A2(new_n740_), .A3(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT106), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT106), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n738_), .A2(new_n747_), .A3(new_n740_), .A4(new_n744_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n746_), .A2(KEYINPUT45), .A3(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(KEYINPUT45), .B1(new_n746_), .B2(new_n748_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT105), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(new_n736_), .B2(new_n451_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n471_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n754_), .B1(new_n434_), .B2(new_n438_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n473_), .B1(new_n389_), .B2(new_n407_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n469_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  AOI211_X1 g556(.A(KEYINPUT43), .B(new_n719_), .C1(new_n757_), .C2(new_n723_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n726_), .B1(new_n725_), .B2(new_n727_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n732_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n734_), .ZN(new_n761_));
  OAI211_X1 g560(.A(KEYINPUT44), .B(new_n732_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n761_), .A2(new_n752_), .A3(new_n451_), .A4(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(G36gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n751_), .B1(new_n753_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT46), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  OAI211_X1 g566(.A(KEYINPUT46), .B(new_n751_), .C1(new_n753_), .C2(new_n764_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(G1329gat));
  AOI21_X1  g568(.A(G43gat), .B1(new_n741_), .B2(new_n468_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n476_), .A2(new_n464_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n736_), .B2(new_n771_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n772_), .B(new_n773_), .ZN(G1330gat));
  AOI21_X1  g573(.A(G50gat), .B1(new_n741_), .B2(new_n473_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n473_), .A2(G50gat), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n736_), .B2(new_n776_), .ZN(G1331gat));
  NOR2_X1   g576(.A1(new_n478_), .A2(new_n518_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n730_), .A2(new_n672_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n439_), .B1(new_n780_), .B2(KEYINPUT108), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n781_), .B1(KEYINPUT108), .B2(new_n780_), .ZN(new_n782_));
  INV_X1    g581(.A(G57gat), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT109), .ZN(new_n785_));
  INV_X1    g584(.A(new_n667_), .ZN(new_n786_));
  AND4_X1   g585(.A1(new_n682_), .A2(new_n519_), .A3(new_n612_), .A4(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(G57gat), .A3(new_n674_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n785_), .A2(new_n788_), .ZN(G1332gat));
  INV_X1    g588(.A(G64gat), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n787_), .B2(new_n451_), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT48), .Z(new_n792_));
  NAND2_X1  g591(.A1(new_n451_), .A2(new_n790_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n792_), .B1(new_n780_), .B2(new_n793_), .ZN(G1333gat));
  NAND2_X1  g593(.A1(new_n787_), .A2(new_n468_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(G71gat), .ZN(new_n796_));
  XNOR2_X1  g595(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n796_), .B(new_n797_), .ZN(new_n798_));
  OR2_X1    g597(.A1(new_n469_), .A2(G71gat), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n780_), .B2(new_n799_), .ZN(G1334gat));
  INV_X1    g599(.A(G78gat), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n787_), .B2(new_n473_), .ZN(new_n802_));
  XOR2_X1   g601(.A(new_n802_), .B(KEYINPUT50), .Z(new_n803_));
  NAND2_X1  g602(.A1(new_n473_), .A2(new_n801_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT111), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n803_), .B1(new_n780_), .B2(new_n805_), .ZN(G1335gat));
  NAND3_X1  g605(.A1(new_n612_), .A2(new_n519_), .A3(new_n667_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT112), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n807_), .B(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n729_), .ZN(new_n810_));
  OAI21_X1  g609(.A(G85gat), .B1(new_n810_), .B2(new_n439_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n730_), .A2(new_n739_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n778_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n814_), .A2(new_n524_), .A3(new_n674_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n811_), .A2(new_n815_), .ZN(G1336gat));
  OAI21_X1  g615(.A(G92gat), .B1(new_n810_), .B2(new_n471_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n814_), .A2(new_n525_), .A3(new_n451_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(G1337gat));
  OAI21_X1  g618(.A(G99gat), .B1(new_n810_), .B2(new_n469_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n814_), .A2(new_n467_), .A3(new_n521_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n820_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g623(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n809_), .A2(new_n473_), .A3(new_n729_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n826_), .B1(new_n827_), .B2(G106gat), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n827_), .A2(new_n826_), .A3(G106gat), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n814_), .A2(new_n522_), .A3(new_n473_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n825_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n830_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n832_), .B(new_n825_), .C1(new_n834_), .C2(new_n828_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n833_), .A2(new_n836_), .ZN(G1339gat));
  INV_X1    g636(.A(KEYINPUT59), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n503_), .B1(new_n501_), .B2(new_n505_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n502_), .B1(new_n508_), .B2(new_n500_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n514_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n506_), .A2(new_n513_), .A3(new_n509_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n600_), .A2(KEYINPUT115), .A3(new_n518_), .ZN(new_n845_));
  AOI21_X1  g644(.A(KEYINPUT115), .B1(new_n600_), .B2(new_n518_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n582_), .A2(KEYINPUT55), .A3(new_n576_), .A4(new_n567_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n575_), .A2(new_n577_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n578_), .A2(new_n584_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n598_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT56), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n853_), .A2(KEYINPUT56), .A3(new_n598_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n608_), .A2(new_n844_), .B1(new_n847_), .B2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n839_), .B1(new_n859_), .B2(new_n681_), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n601_), .A2(new_n520_), .A3(new_n602_), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT70), .B1(new_n606_), .B2(new_n600_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n844_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n846_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n600_), .A2(KEYINPUT115), .A3(new_n518_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n858_), .A2(new_n864_), .A3(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n863_), .A2(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(KEYINPUT57), .A3(new_n680_), .ZN(new_n868_));
  AOI21_X1  g667(.A(KEYINPUT117), .B1(new_n860_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870_));
  AOI21_X1  g669(.A(KEYINPUT56), .B1(new_n853_), .B2(new_n598_), .ZN(new_n871_));
  AOI211_X1 g670(.A(new_n855_), .B(new_n599_), .C1(new_n850_), .C2(new_n852_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n871_), .A2(new_n872_), .A3(KEYINPUT118), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n854_), .A2(KEYINPUT118), .A3(new_n855_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n600_), .A2(new_n844_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n870_), .B1(new_n873_), .B2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT118), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n856_), .A2(new_n878_), .A3(new_n857_), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n879_), .A2(KEYINPUT58), .A3(new_n874_), .A4(new_n875_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n877_), .A2(new_n727_), .A3(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(KEYINPUT57), .B1(new_n867_), .B2(new_n680_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT117), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n881_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n684_), .B1(new_n869_), .B2(new_n884_), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n671_), .A2(new_n610_), .A3(new_n519_), .A4(new_n611_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n886_), .B(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n885_), .A2(new_n889_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n475_), .A2(new_n674_), .A3(new_n467_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  AND2_X1   g691(.A1(new_n892_), .A2(KEYINPUT119), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n892_), .A2(KEYINPUT119), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n838_), .B1(new_n890_), .B2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n838_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n860_), .A2(new_n868_), .A3(new_n881_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n667_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n888_), .B1(new_n899_), .B2(KEYINPUT120), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n898_), .A2(new_n901_), .A3(new_n667_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n897_), .B1(new_n900_), .B2(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(KEYINPUT121), .B1(new_n896_), .B2(new_n903_), .ZN(new_n904_));
  AOI211_X1 g703(.A(new_n839_), .B(new_n681_), .C1(new_n863_), .C2(new_n866_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n883_), .B1(new_n882_), .B2(new_n905_), .ZN(new_n906_));
  AND3_X1   g705(.A1(new_n877_), .A2(new_n727_), .A3(new_n880_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n907_), .B1(new_n860_), .B2(KEYINPUT117), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n888_), .B1(new_n909_), .B2(new_n684_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n895_), .ZN(new_n911_));
  OAI21_X1  g710(.A(KEYINPUT59), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n899_), .A2(KEYINPUT120), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n913_), .A2(new_n889_), .A3(new_n902_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n897_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n912_), .A2(new_n916_), .A3(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(G113gat), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n519_), .A2(new_n919_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n904_), .A2(new_n918_), .A3(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n910_), .A2(new_n911_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n919_), .B1(new_n923_), .B2(new_n519_), .ZN(new_n924_));
  AND2_X1   g723(.A1(new_n921_), .A2(new_n924_), .ZN(G1340gat));
  INV_X1    g724(.A(G120gat), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n926_), .B1(new_n730_), .B2(KEYINPUT60), .ZN(new_n927_));
  OAI211_X1 g726(.A(new_n922_), .B(new_n927_), .C1(KEYINPUT60), .C2(new_n926_), .ZN(new_n928_));
  NOR3_X1   g727(.A1(new_n896_), .A2(new_n903_), .A3(new_n730_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n929_), .B2(new_n926_), .ZN(G1341gat));
  INV_X1    g729(.A(G127gat), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n684_), .A2(new_n931_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n904_), .A2(new_n918_), .A3(new_n932_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n931_), .B1(new_n923_), .B2(new_n667_), .ZN(new_n934_));
  AND2_X1   g733(.A1(new_n933_), .A2(new_n934_), .ZN(G1342gat));
  XOR2_X1   g734(.A(KEYINPUT123), .B(G134gat), .Z(new_n936_));
  NOR2_X1   g735(.A1(new_n719_), .A2(new_n936_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n904_), .A2(new_n918_), .A3(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n683_), .B1(new_n906_), .B2(new_n908_), .ZN(new_n939_));
  OAI211_X1 g738(.A(new_n895_), .B(new_n681_), .C1(new_n939_), .C2(new_n888_), .ZN(new_n940_));
  INV_X1    g739(.A(G134gat), .ZN(new_n941_));
  AND3_X1   g740(.A1(new_n940_), .A2(KEYINPUT122), .A3(new_n941_), .ZN(new_n942_));
  AOI21_X1  g741(.A(KEYINPUT122), .B1(new_n940_), .B2(new_n941_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n942_), .A2(new_n943_), .ZN(new_n944_));
  AND2_X1   g743(.A1(new_n938_), .A2(new_n944_), .ZN(G1343gat));
  NOR2_X1   g744(.A1(new_n439_), .A2(new_n754_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n890_), .A2(new_n469_), .A3(new_n946_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n947_), .A2(new_n519_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(new_n212_), .ZN(G1344gat));
  NOR2_X1   g748(.A1(new_n947_), .A2(new_n730_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(new_n213_), .ZN(G1345gat));
  OAI21_X1  g750(.A(KEYINPUT124), .B1(new_n947_), .B2(new_n667_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n468_), .B1(new_n885_), .B2(new_n889_), .ZN(new_n953_));
  INV_X1    g752(.A(KEYINPUT124), .ZN(new_n954_));
  NAND4_X1  g753(.A1(new_n953_), .A2(new_n954_), .A3(new_n786_), .A4(new_n946_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(KEYINPUT61), .B(G155gat), .ZN(new_n956_));
  AND3_X1   g755(.A1(new_n952_), .A2(new_n955_), .A3(new_n956_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n956_), .B1(new_n952_), .B2(new_n955_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n957_), .A2(new_n958_), .ZN(G1346gat));
  OAI21_X1  g758(.A(G162gat), .B1(new_n947_), .B2(new_n719_), .ZN(new_n960_));
  OR2_X1    g759(.A1(new_n680_), .A2(G162gat), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n960_), .B1(new_n947_), .B2(new_n961_), .ZN(G1347gat));
  NOR3_X1   g761(.A1(new_n674_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n963_));
  INV_X1    g762(.A(new_n963_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n964_), .A2(new_n473_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n914_), .A2(new_n965_), .ZN(new_n966_));
  OAI21_X1  g765(.A(G169gat), .B1(new_n966_), .B2(new_n519_), .ZN(new_n967_));
  INV_X1    g766(.A(KEYINPUT62), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n967_), .A2(new_n968_), .ZN(new_n969_));
  INV_X1    g768(.A(new_n966_), .ZN(new_n970_));
  NAND4_X1  g769(.A1(new_n970_), .A2(new_n317_), .A3(new_n319_), .A4(new_n518_), .ZN(new_n971_));
  OAI211_X1 g770(.A(KEYINPUT62), .B(G169gat), .C1(new_n966_), .C2(new_n519_), .ZN(new_n972_));
  NAND3_X1  g771(.A1(new_n969_), .A2(new_n971_), .A3(new_n972_), .ZN(G1348gat));
  NAND2_X1  g772(.A1(new_n970_), .A2(new_n612_), .ZN(new_n974_));
  AND2_X1   g773(.A1(new_n315_), .A2(new_n320_), .ZN(new_n975_));
  NOR2_X1   g774(.A1(new_n910_), .A2(new_n473_), .ZN(new_n976_));
  NOR3_X1   g775(.A1(new_n964_), .A2(new_n730_), .A3(new_n358_), .ZN(new_n977_));
  AOI22_X1  g776(.A1(new_n974_), .A2(new_n975_), .B1(new_n976_), .B2(new_n977_), .ZN(G1349gat));
  NAND3_X1  g777(.A1(new_n976_), .A2(new_n786_), .A3(new_n963_), .ZN(new_n979_));
  INV_X1    g778(.A(new_n355_), .ZN(new_n980_));
  NOR3_X1   g779(.A1(new_n684_), .A2(new_n304_), .A3(new_n303_), .ZN(new_n981_));
  AOI22_X1  g780(.A1(new_n979_), .A2(new_n980_), .B1(new_n970_), .B2(new_n981_), .ZN(G1350gat));
  OAI21_X1  g781(.A(G190gat), .B1(new_n966_), .B2(new_n719_), .ZN(new_n983_));
  NAND2_X1  g782(.A1(new_n681_), .A2(new_n363_), .ZN(new_n984_));
  XNOR2_X1  g783(.A(new_n984_), .B(KEYINPUT125), .ZN(new_n985_));
  OAI21_X1  g784(.A(new_n983_), .B1(new_n966_), .B2(new_n985_), .ZN(G1351gat));
  NAND4_X1  g785(.A1(new_n953_), .A2(new_n439_), .A3(new_n473_), .A4(new_n451_), .ZN(new_n987_));
  NOR2_X1   g786(.A1(new_n987_), .A2(new_n519_), .ZN(new_n988_));
  XNOR2_X1  g787(.A(new_n988_), .B(new_n330_), .ZN(G1352gat));
  NOR2_X1   g788(.A1(new_n987_), .A2(new_n730_), .ZN(new_n990_));
  OR2_X1    g789(.A1(new_n331_), .A2(KEYINPUT126), .ZN(new_n991_));
  XNOR2_X1  g790(.A(new_n990_), .B(new_n991_), .ZN(G1353gat));
  INV_X1    g791(.A(new_n987_), .ZN(new_n993_));
  XOR2_X1   g792(.A(KEYINPUT63), .B(G211gat), .Z(new_n994_));
  NAND3_X1  g793(.A1(new_n993_), .A2(new_n683_), .A3(new_n994_), .ZN(new_n995_));
  NOR2_X1   g794(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n996_));
  OAI21_X1  g795(.A(new_n996_), .B1(new_n987_), .B2(new_n684_), .ZN(new_n997_));
  AND2_X1   g796(.A1(new_n995_), .A2(new_n997_), .ZN(G1354gat));
  XOR2_X1   g797(.A(KEYINPUT127), .B(G218gat), .Z(new_n999_));
  NOR3_X1   g798(.A1(new_n987_), .A2(new_n719_), .A3(new_n999_), .ZN(new_n1000_));
  NAND2_X1  g799(.A1(new_n993_), .A2(new_n681_), .ZN(new_n1001_));
  AOI21_X1  g800(.A(new_n1000_), .B1(new_n1001_), .B2(new_n999_), .ZN(G1355gat));
endmodule


