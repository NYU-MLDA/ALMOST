//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n932_, new_n933_, new_n935_, new_n936_, new_n937_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_;
  NAND2_X1  g000(.A1(KEYINPUT75), .A2(KEYINPUT37), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT75), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT37), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT36), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G232gat), .A2(G233gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT34), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT74), .B1(new_n208_), .B2(KEYINPUT35), .ZN(new_n209_));
  OR2_X1    g008(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n210_));
  INV_X1    g009(.A(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G85gat), .ZN(new_n214_));
  INV_X1    g013(.A(G92gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G85gat), .A2(G92gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(KEYINPUT9), .A3(new_n217_), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n217_), .A2(KEYINPUT9), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n213_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G99gat), .A2(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT6), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT6), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(G99gat), .A3(G106gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n224_), .A3(KEYINPUT65), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n223_), .B1(G99gat), .B2(G106gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n221_), .A2(KEYINPUT6), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n226_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n220_), .B1(new_n225_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n222_), .A2(new_n224_), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT7), .ZN(new_n233_));
  INV_X1    g032(.A(G99gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(new_n234_), .A3(new_n211_), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n231_), .A2(new_n232_), .A3(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n237_));
  AND2_X1   g036(.A1(G85gat), .A2(G92gat), .ZN(new_n238_));
  NOR2_X1   g037(.A1(G85gat), .A2(G92gat), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n237_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n216_), .A2(KEYINPUT66), .A3(new_n217_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT8), .B1(new_n236_), .B2(new_n242_), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n235_), .A2(new_n232_), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n222_), .A2(new_n224_), .A3(KEYINPUT65), .ZN(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT65), .B1(new_n222_), .B2(new_n224_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n244_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT8), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n240_), .A2(new_n241_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n247_), .A2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n230_), .B1(new_n243_), .B2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G29gat), .B(G36gat), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(G43gat), .B(G50gat), .Z(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G43gat), .B(G50gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n253_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n209_), .B1(new_n252_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT71), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT15), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n259_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n256_), .A2(KEYINPUT15), .A3(new_n258_), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n229_), .A2(new_n225_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n266_), .A2(new_n213_), .A3(new_n218_), .A4(new_n219_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n249_), .B1(new_n266_), .B2(new_n244_), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n240_), .A2(new_n241_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n231_), .A2(new_n232_), .A3(new_n235_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n248_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n267_), .B1(new_n268_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n265_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n260_), .A2(new_n261_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n261_), .B1(new_n260_), .B2(new_n273_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT35), .ZN(new_n277_));
  INV_X1    g076(.A(new_n208_), .ZN(new_n278_));
  OAI22_X1  g077(.A1(new_n275_), .A2(new_n276_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n276_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n278_), .A2(new_n277_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n280_), .A2(new_n281_), .A3(new_n274_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G190gat), .B(G218gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT72), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G134gat), .B(G162gat), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n284_), .B(new_n285_), .Z(new_n286_));
  NAND3_X1  g085(.A1(new_n279_), .A2(new_n282_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n279_), .A2(new_n282_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n286_), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n206_), .A2(new_n287_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n289_), .A2(new_n206_), .A3(new_n290_), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n202_), .B(new_n205_), .C1(new_n291_), .C2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n289_), .A2(new_n290_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n287_), .A2(new_n206_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n289_), .A2(new_n206_), .A3(new_n290_), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n296_), .A2(new_n203_), .A3(new_n204_), .A4(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n293_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT77), .ZN(new_n300_));
  INV_X1    g099(.A(G1gat), .ZN(new_n301_));
  INV_X1    g100(.A(G8gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT14), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT76), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT76), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n305_), .B(KEYINPUT14), .C1(new_n301_), .C2(new_n302_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G15gat), .B(G22gat), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n304_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(G1gat), .B(G8gat), .Z(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n304_), .A2(new_n309_), .A3(new_n306_), .A4(new_n307_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(G231gat), .A3(G233gat), .ZN(new_n314_));
  INV_X1    g113(.A(G231gat), .ZN(new_n315_));
  INV_X1    g114(.A(G233gat), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n311_), .B(new_n312_), .C1(new_n315_), .C2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G57gat), .B(G64gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G71gat), .B(G78gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n318_), .A2(new_n319_), .A3(KEYINPUT11), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(KEYINPUT11), .ZN(new_n321_));
  INV_X1    g120(.A(new_n319_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n318_), .A2(KEYINPUT11), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n320_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n314_), .A2(new_n317_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n326_), .B1(new_n314_), .B2(new_n317_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n300_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n329_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n331_), .A2(KEYINPUT77), .A3(new_n327_), .ZN(new_n332_));
  XOR2_X1   g131(.A(G127gat), .B(G155gat), .Z(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT16), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G183gat), .B(G211gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT17), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n330_), .A2(new_n332_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT78), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n340_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n331_), .A2(KEYINPUT78), .A3(new_n327_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n336_), .B(KEYINPUT17), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n339_), .A2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT12), .B1(new_n252_), .B2(new_n325_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT12), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n272_), .A2(new_n347_), .A3(new_n326_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n267_), .B(new_n325_), .C1(new_n268_), .C2(new_n271_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G230gat), .A2(G233gat), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n351_), .B(KEYINPUT64), .Z(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n350_), .A2(KEYINPUT68), .A3(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n350_), .A2(new_n353_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT68), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n349_), .A2(new_n354_), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n272_), .A2(new_n326_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n359_), .A2(KEYINPUT67), .A3(new_n350_), .ZN(new_n360_));
  OR3_X1    g159(.A1(new_n252_), .A2(KEYINPUT67), .A3(new_n325_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n361_), .A3(new_n352_), .ZN(new_n362_));
  XOR2_X1   g161(.A(KEYINPUT69), .B(KEYINPUT5), .Z(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT70), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G120gat), .B(G148gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G176gat), .B(G204gat), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n366_), .B(new_n367_), .Z(new_n368_));
  AND3_X1   g167(.A1(new_n358_), .A2(new_n362_), .A3(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n368_), .B1(new_n358_), .B2(new_n362_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT13), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT13), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n373_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n299_), .A2(new_n345_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n313_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G229gat), .A2(G233gat), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n311_), .A2(new_n259_), .A3(new_n312_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n380_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n311_), .A2(new_n259_), .A3(new_n312_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n259_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n383_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G113gat), .B(G141gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT80), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G169gat), .B(G197gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n382_), .A2(new_n386_), .A3(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT81), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n390_), .B1(new_n382_), .B2(new_n386_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  AOI211_X1 g194(.A(new_n392_), .B(new_n390_), .C1(new_n382_), .C2(new_n386_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G113gat), .B(G120gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT87), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G127gat), .B(G134gat), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT87), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n398_), .B(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(new_n400_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT88), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n402_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n399_), .A2(KEYINPUT88), .A3(new_n401_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT89), .ZN(new_n410_));
  NOR2_X1   g209(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n411_));
  INV_X1    g210(.A(G169gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G183gat), .A2(G190gat), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT23), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT85), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT82), .B(G183gat), .ZN(new_n418_));
  OR2_X1    g217(.A1(new_n418_), .A2(G190gat), .ZN(new_n419_));
  OR3_X1    g218(.A1(new_n414_), .A2(KEYINPUT85), .A3(KEYINPUT23), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n417_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n413_), .B1(new_n421_), .B2(KEYINPUT86), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT86), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n417_), .A2(new_n419_), .A3(new_n423_), .A4(new_n420_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(G176gat), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n412_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT24), .ZN(new_n428_));
  NOR2_X1   g227(.A1(G169gat), .A2(G176gat), .ZN(new_n429_));
  NOR3_X1   g228(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT84), .ZN(new_n431_));
  INV_X1    g230(.A(new_n416_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n429_), .A2(new_n428_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n430_), .A2(KEYINPUT84), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n418_), .A2(KEYINPUT25), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n437_), .B1(KEYINPUT25), .B2(G183gat), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT26), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT83), .B1(new_n439_), .B2(G190gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(KEYINPUT26), .B(G190gat), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n438_), .B(new_n440_), .C1(KEYINPUT83), .C2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n436_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n425_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G71gat), .B(G99gat), .ZN(new_n445_));
  INV_X1    g244(.A(G43gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT30), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n444_), .A2(new_n449_), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n424_), .A2(new_n422_), .B1(new_n436_), .B2(new_n442_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n448_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G227gat), .A2(G233gat), .ZN(new_n454_));
  INV_X1    g253(.A(G15gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n410_), .B1(new_n453_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT31), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n450_), .A2(new_n452_), .A3(new_n456_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n459_), .B1(new_n458_), .B2(new_n460_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n409_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n458_), .A2(new_n460_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT31), .ZN(new_n466_));
  INV_X1    g265(.A(new_n409_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n466_), .A2(new_n467_), .A3(new_n461_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n464_), .A2(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(G1gat), .B(G29gat), .Z(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT103), .B(KEYINPUT0), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G57gat), .B(G85gat), .ZN(new_n473_));
  XOR2_X1   g272(.A(new_n472_), .B(new_n473_), .Z(new_n474_));
  XOR2_X1   g273(.A(G155gat), .B(G162gat), .Z(new_n475_));
  NOR2_X1   g274(.A1(G141gat), .A2(G148gat), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT3), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G141gat), .A2(G148gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT92), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n478_), .B(new_n479_), .C1(new_n481_), .C2(KEYINPUT2), .ZN(new_n482_));
  AND2_X1   g281(.A1(new_n481_), .A2(KEYINPUT2), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n475_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT93), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  OAI211_X1 g285(.A(KEYINPUT93), .B(new_n475_), .C1(new_n482_), .C2(new_n483_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G155gat), .A2(G162gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(G155gat), .A2(G162gat), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n489_), .B1(new_n490_), .B2(KEYINPUT1), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT90), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  OAI211_X1 g292(.A(KEYINPUT90), .B(new_n489_), .C1(new_n490_), .C2(KEYINPUT1), .ZN(new_n494_));
  OR3_X1    g293(.A1(new_n489_), .A2(KEYINPUT91), .A3(KEYINPUT1), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT91), .B1(new_n489_), .B2(KEYINPUT1), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n493_), .A2(new_n494_), .A3(new_n495_), .A4(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n480_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n498_), .A2(new_n476_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n488_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n409_), .A2(new_n501_), .ZN(new_n502_));
  AOI22_X1  g301(.A1(new_n486_), .A2(new_n487_), .B1(new_n497_), .B2(new_n499_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n402_), .A2(new_n405_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n502_), .A2(KEYINPUT4), .A3(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G225gat), .A2(G233gat), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT4), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n409_), .A2(new_n501_), .A3(new_n509_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n506_), .A2(KEYINPUT102), .A3(new_n508_), .A4(new_n510_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n502_), .A2(new_n505_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n507_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n510_), .A2(new_n508_), .ZN(new_n515_));
  AOI21_X1  g314(.A(KEYINPUT102), .B1(new_n515_), .B2(new_n506_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n474_), .B1(new_n514_), .B2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n506_), .A2(new_n508_), .A3(new_n510_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT102), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n474_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n520_), .A2(new_n521_), .A3(new_n511_), .A4(new_n513_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n517_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G226gat), .A2(G233gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT19), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G211gat), .B(G218gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT94), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G197gat), .B(G204gat), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n529_), .A2(KEYINPUT96), .ZN(new_n530_));
  OAI21_X1  g329(.A(KEYINPUT21), .B1(new_n529_), .B2(KEYINPUT96), .ZN(new_n531_));
  OR3_X1    g330(.A1(new_n528_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n529_), .B(KEYINPUT21), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n528_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT95), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT95), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n528_), .A2(new_n533_), .A3(new_n536_), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n532_), .A2(new_n535_), .A3(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(KEYINPUT22), .B(G169gat), .Z(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT101), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n426_), .ZN(new_n541_));
  OR2_X1    g340(.A1(G183gat), .A2(G190gat), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n427_), .B1(new_n432_), .B2(new_n542_), .ZN(new_n543_));
  NOR3_X1   g342(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT25), .B(G183gat), .ZN(new_n545_));
  AOI211_X1 g344(.A(new_n544_), .B(new_n430_), .C1(new_n441_), .C2(new_n545_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n417_), .A2(new_n420_), .ZN(new_n547_));
  AOI22_X1  g346(.A1(new_n541_), .A2(new_n543_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT20), .B1(new_n538_), .B2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n532_), .A2(new_n535_), .A3(new_n537_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n444_), .A2(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n526_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G8gat), .B(G36gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT18), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G64gat), .B(G92gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT20), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n558_), .B1(new_n538_), .B2(new_n548_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n526_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n444_), .A2(new_n550_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n559_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n552_), .A2(new_n557_), .A3(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT27), .ZN(new_n564_));
  NOR3_X1   g363(.A1(new_n549_), .A2(new_n551_), .A3(new_n526_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n560_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n564_), .B1(new_n556_), .B2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT106), .B(KEYINPUT27), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n557_), .B1(new_n552_), .B2(new_n562_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n569_), .B1(new_n571_), .B2(new_n563_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n568_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT29), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n503_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT28), .ZN(new_n576_));
  XOR2_X1   g375(.A(G22gat), .B(G50gat), .Z(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(G228gat), .ZN(new_n579_));
  OAI221_X1 g378(.A(new_n550_), .B1(new_n579_), .B2(new_n316_), .C1(new_n574_), .C2(new_n503_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT97), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n501_), .A2(new_n581_), .A3(KEYINPUT29), .ZN(new_n582_));
  OAI21_X1  g381(.A(KEYINPUT97), .B1(new_n503_), .B2(new_n574_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(new_n583_), .A3(new_n550_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n579_), .A2(new_n316_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT98), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(KEYINPUT98), .B1(new_n584_), .B2(new_n585_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n580_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G78gat), .B(G106gat), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n578_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n586_), .B(new_n587_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n591_), .B(KEYINPUT99), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n593_), .A2(KEYINPUT100), .A3(new_n594_), .A4(new_n580_), .ZN(new_n595_));
  OAI211_X1 g394(.A(new_n594_), .B(new_n580_), .C1(new_n588_), .C2(new_n589_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT100), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n592_), .A2(new_n595_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n578_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n594_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n590_), .A2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n600_), .B1(new_n602_), .B2(new_n596_), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n524_), .B(new_n573_), .C1(new_n599_), .C2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n514_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n605_), .A2(KEYINPUT33), .A3(new_n521_), .A4(new_n520_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT33), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n522_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n563_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n609_), .A2(new_n570_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n506_), .A2(new_n507_), .A3(new_n510_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT104), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n612_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n521_), .B1(new_n512_), .B2(new_n508_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n613_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n606_), .A2(new_n608_), .A3(new_n610_), .A4(new_n616_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n557_), .A2(KEYINPUT32), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n618_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n559_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n541_), .A2(new_n543_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n546_), .A2(new_n547_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n558_), .B1(new_n623_), .B2(new_n550_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n538_), .A2(new_n451_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n560_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NOR3_X1   g425(.A1(new_n620_), .A2(new_n626_), .A3(new_n618_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT105), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n619_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n567_), .A2(KEYINPUT105), .A3(new_n618_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n523_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n617_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n602_), .A2(new_n596_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(new_n578_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n592_), .A2(new_n595_), .A3(new_n598_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n632_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n469_), .B1(new_n604_), .B2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n634_), .A2(new_n635_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n469_), .A2(new_n524_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n573_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n638_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n397_), .B1(new_n637_), .B2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n378_), .A2(new_n642_), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n524_), .A2(KEYINPUT107), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n524_), .A2(KEYINPUT107), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n643_), .A2(new_n301_), .A3(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(KEYINPUT108), .B(KEYINPUT38), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n291_), .A2(new_n292_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n651_), .A2(new_n345_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n393_), .B(new_n394_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n375_), .A2(new_n653_), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n652_), .B(new_n654_), .C1(new_n637_), .C2(new_n641_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G1gat), .B1(new_n655_), .B2(new_n524_), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n647_), .A2(new_n648_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n657_), .A2(KEYINPUT109), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(KEYINPUT109), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n649_), .B(new_n656_), .C1(new_n658_), .C2(new_n659_), .ZN(G1324gat));
  XNOR2_X1  g459(.A(KEYINPUT110), .B(KEYINPUT111), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT40), .ZN(new_n662_));
  OAI21_X1  g461(.A(G8gat), .B1(new_n655_), .B2(new_n573_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT39), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT39), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n665_), .B(G8gat), .C1(new_n655_), .C2(new_n573_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  NOR4_X1   g466(.A1(new_n378_), .A2(new_n642_), .A3(G8gat), .A4(new_n573_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n662_), .B1(new_n667_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n667_), .A2(new_n669_), .A3(new_n662_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n661_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n672_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n661_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n674_), .A2(new_n670_), .A3(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n673_), .A2(new_n676_), .ZN(G1325gat));
  INV_X1    g476(.A(new_n469_), .ZN(new_n678_));
  OAI21_X1  g477(.A(G15gat), .B1(new_n655_), .B2(new_n678_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT41), .Z(new_n680_));
  NAND3_X1  g479(.A1(new_n643_), .A2(new_n455_), .A3(new_n469_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1326gat));
  XNOR2_X1  g481(.A(new_n638_), .B(KEYINPUT112), .ZN(new_n683_));
  OAI21_X1  g482(.A(G22gat), .B1(new_n655_), .B2(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT42), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n683_), .A2(G22gat), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n643_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(G1327gat));
  NAND2_X1  g487(.A1(new_n604_), .A2(new_n636_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n641_), .B1(new_n689_), .B2(new_n678_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n690_), .A2(new_n375_), .A3(new_n653_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n339_), .A2(new_n344_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n650_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G29gat), .B1(new_n695_), .B2(new_n523_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n299_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT43), .B1(new_n690_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT43), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n699_), .B(new_n299_), .C1(new_n637_), .C2(new_n641_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n654_), .A2(new_n345_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT44), .B1(new_n701_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705_));
  AOI211_X1 g504(.A(new_n705_), .B(new_n702_), .C1(new_n698_), .C2(new_n700_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n704_), .A2(new_n706_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n646_), .A2(G29gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n696_), .B1(new_n707_), .B2(new_n708_), .ZN(G1328gat));
  NOR2_X1   g508(.A1(new_n573_), .A2(G36gat), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  OR3_X1    g510(.A1(new_n694_), .A2(KEYINPUT45), .A3(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(KEYINPUT45), .B1(new_n694_), .B2(new_n711_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n704_), .A2(new_n706_), .A3(new_n573_), .ZN(new_n715_));
  INV_X1    g514(.A(G36gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n714_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT46), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  OAI211_X1 g518(.A(KEYINPUT46), .B(new_n714_), .C1(new_n715_), .C2(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1329gat));
  NOR2_X1   g520(.A1(new_n678_), .A2(new_n446_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n707_), .A2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n446_), .B1(new_n694_), .B2(new_n678_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT47), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT47), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n723_), .A2(new_n727_), .A3(new_n724_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1330gat));
  OR3_X1    g528(.A1(new_n694_), .A2(G50gat), .A3(new_n683_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n707_), .A2(KEYINPUT113), .A3(new_n638_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(G50gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(KEYINPUT113), .B1(new_n707_), .B2(new_n638_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n730_), .B1(new_n732_), .B2(new_n733_), .ZN(G1331gat));
  INV_X1    g533(.A(new_n375_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n690_), .A2(new_n735_), .A3(new_n397_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(new_n652_), .ZN(new_n737_));
  OAI21_X1  g536(.A(G57gat), .B1(new_n737_), .B2(new_n524_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n736_), .A2(new_n697_), .A3(new_n692_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n646_), .ZN(new_n740_));
  OR2_X1    g539(.A1(new_n740_), .A2(G57gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n738_), .B1(new_n739_), .B2(new_n741_), .ZN(G1332gat));
  OAI21_X1  g541(.A(G64gat), .B1(new_n737_), .B2(new_n573_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT48), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n573_), .A2(G64gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n744_), .B1(new_n739_), .B2(new_n745_), .ZN(G1333gat));
  OAI21_X1  g545(.A(G71gat), .B1(new_n737_), .B2(new_n678_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT49), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n678_), .A2(G71gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n739_), .B2(new_n749_), .ZN(G1334gat));
  OAI21_X1  g549(.A(G78gat), .B1(new_n737_), .B2(new_n683_), .ZN(new_n751_));
  XOR2_X1   g550(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n752_));
  XNOR2_X1  g551(.A(new_n751_), .B(new_n752_), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n683_), .A2(G78gat), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n753_), .B1(new_n739_), .B2(new_n754_), .ZN(G1335gat));
  NAND3_X1  g554(.A1(new_n375_), .A2(new_n345_), .A3(new_n653_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n698_), .B2(new_n700_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(G85gat), .B1(new_n758_), .B2(new_n524_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n736_), .A2(new_n693_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(new_n214_), .A3(new_n646_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n759_), .A2(new_n762_), .ZN(G1336gat));
  OAI21_X1  g562(.A(G92gat), .B1(new_n758_), .B2(new_n573_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n761_), .A2(new_n215_), .A3(new_n640_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(G1337gat));
  OAI21_X1  g565(.A(G99gat), .B1(new_n758_), .B2(new_n678_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n469_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n760_), .B2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g569(.A1(new_n761_), .A2(new_n211_), .A3(new_n638_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n757_), .A2(new_n638_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n773_), .B2(G106gat), .ZN(new_n774_));
  AOI211_X1 g573(.A(KEYINPUT52), .B(new_n211_), .C1(new_n757_), .C2(new_n638_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n771_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT53), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n778_), .B(new_n771_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(G1339gat));
  NOR4_X1   g579(.A1(new_n740_), .A2(new_n638_), .A3(new_n640_), .A4(new_n678_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n380_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n390_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT119), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n379_), .A2(new_n383_), .A3(new_n381_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n782_), .A2(KEYINPUT119), .A3(new_n783_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n786_), .A2(new_n787_), .A3(KEYINPUT120), .A4(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n391_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n787_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n259_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n313_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n381_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n390_), .B1(new_n794_), .B2(new_n380_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n791_), .B1(new_n795_), .B2(KEYINPUT119), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT120), .B1(new_n796_), .B2(new_n786_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n790_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT121), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n798_), .B(new_n799_), .C1(new_n370_), .C2(new_n369_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT120), .ZN(new_n801_));
  INV_X1    g600(.A(new_n786_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n788_), .A2(new_n787_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n801_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n804_), .A2(new_n391_), .A3(new_n789_), .ZN(new_n805_));
  OAI21_X1  g604(.A(KEYINPUT121), .B1(new_n371_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n800_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n349_), .A2(new_n357_), .A3(KEYINPUT55), .A4(new_n354_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT117), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n350_), .A2(KEYINPUT68), .A3(new_n353_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT68), .B1(new_n350_), .B2(new_n353_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n813_), .A2(new_n814_), .A3(KEYINPUT55), .A4(new_n349_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n357_), .A2(new_n354_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n252_), .A2(KEYINPUT12), .A3(new_n325_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n347_), .B1(new_n272_), .B2(new_n326_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n816_), .B1(new_n817_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n350_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n352_), .B1(new_n820_), .B2(new_n822_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n810_), .A2(new_n815_), .A3(new_n821_), .A4(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n368_), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n824_), .A2(KEYINPUT56), .A3(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT56), .B1(new_n824_), .B2(new_n825_), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n826_), .A2(new_n827_), .A3(KEYINPUT118), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n824_), .A2(new_n825_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT56), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(KEYINPUT118), .A3(new_n830_), .ZN(new_n831_));
  OR2_X1    g630(.A1(new_n653_), .A2(new_n369_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n808_), .B1(new_n828_), .B2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n835_), .A2(KEYINPUT57), .A3(new_n650_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n829_), .A2(new_n830_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n824_), .A2(KEYINPUT56), .A3(new_n825_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n838_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n832_), .B1(new_n827_), .B2(KEYINPUT118), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n807_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n837_), .B1(new_n843_), .B2(new_n651_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n805_), .A2(new_n369_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT58), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  OAI211_X1 g647(.A(KEYINPUT58), .B(new_n845_), .C1(new_n826_), .C2(new_n827_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n299_), .A2(new_n848_), .A3(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n836_), .A2(new_n844_), .A3(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n345_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT115), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n692_), .A2(new_n853_), .A3(new_n653_), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT115), .B1(new_n345_), .B2(new_n397_), .ZN(new_n855_));
  AND4_X1   g654(.A1(new_n374_), .A2(new_n372_), .A3(new_n854_), .A4(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n293_), .A2(new_n856_), .A3(new_n298_), .ZN(new_n857_));
  XOR2_X1   g656(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n293_), .A2(new_n856_), .A3(new_n298_), .A4(new_n858_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(KEYINPUT122), .B1(new_n852_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n865_));
  AOI211_X1 g664(.A(new_n865_), .B(new_n862_), .C1(new_n851_), .C2(new_n345_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n781_), .B1(new_n864_), .B2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(G113gat), .B1(new_n868_), .B2(new_n397_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n862_), .B1(new_n851_), .B2(new_n345_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT59), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n781_), .A2(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n870_), .A2(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n873_), .B1(new_n867_), .B2(KEYINPUT59), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n397_), .A2(G113gat), .ZN(new_n875_));
  XOR2_X1   g674(.A(new_n875_), .B(KEYINPUT123), .Z(new_n876_));
  AOI21_X1  g675(.A(new_n869_), .B1(new_n874_), .B2(new_n876_), .ZN(G1340gat));
  INV_X1    g676(.A(G120gat), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n878_), .B1(new_n874_), .B2(new_n375_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n735_), .B2(KEYINPUT60), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(KEYINPUT60), .B2(new_n878_), .ZN(new_n881_));
  OR2_X1    g680(.A1(new_n867_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(KEYINPUT124), .B1(new_n879_), .B2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT124), .ZN(new_n885_));
  AOI211_X1 g684(.A(new_n735_), .B(new_n873_), .C1(new_n867_), .C2(KEYINPUT59), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n885_), .B(new_n882_), .C1(new_n886_), .C2(new_n878_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n884_), .A2(new_n887_), .ZN(G1341gat));
  INV_X1    g687(.A(G127gat), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n868_), .A2(new_n889_), .A3(new_n692_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n874_), .A2(new_n692_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n889_), .ZN(G1342gat));
  INV_X1    g691(.A(G134gat), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n868_), .A2(new_n893_), .A3(new_n651_), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n874_), .A2(new_n299_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(new_n893_), .ZN(G1343gat));
  OR2_X1    g695(.A1(new_n864_), .A2(new_n866_), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n740_), .A2(new_n469_), .A3(new_n640_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n897_), .A2(new_n638_), .A3(new_n898_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(new_n653_), .ZN(new_n900_));
  INV_X1    g699(.A(G141gat), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(G1344gat));
  NOR2_X1   g701(.A1(new_n899_), .A2(new_n735_), .ZN(new_n903_));
  INV_X1    g702(.A(G148gat), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1345gat));
  NOR2_X1   g704(.A1(new_n899_), .A2(new_n345_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT61), .B(G155gat), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n906_), .B(new_n908_), .ZN(G1346gat));
  OAI21_X1  g708(.A(G162gat), .B1(new_n899_), .B2(new_n697_), .ZN(new_n910_));
  OR2_X1    g709(.A1(new_n650_), .A2(G162gat), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n899_), .B2(new_n911_), .ZN(G1347gat));
  NOR3_X1   g711(.A1(new_n646_), .A2(new_n573_), .A3(new_n678_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n683_), .A2(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n870_), .A2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  OAI21_X1  g715(.A(G169gat), .B1(new_n916_), .B2(new_n653_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n917_), .A2(KEYINPUT62), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n917_), .A2(KEYINPUT62), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n915_), .A2(new_n540_), .A3(new_n397_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n918_), .B1(new_n919_), .B2(new_n920_), .ZN(G1348gat));
  AOI21_X1  g720(.A(G176gat), .B1(new_n915_), .B2(new_n375_), .ZN(new_n922_));
  AND3_X1   g721(.A1(new_n897_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n923_));
  AND3_X1   g722(.A1(new_n913_), .A2(G176gat), .A3(new_n375_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n922_), .B1(new_n923_), .B2(new_n924_), .ZN(G1349gat));
  AND2_X1   g724(.A1(new_n913_), .A2(new_n692_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n418_), .B1(new_n923_), .B2(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n545_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n915_), .A2(new_n692_), .A3(new_n928_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(KEYINPUT125), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n927_), .A2(new_n930_), .ZN(G1350gat));
  OAI21_X1  g730(.A(G190gat), .B1(new_n916_), .B2(new_n697_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n915_), .A2(new_n651_), .A3(new_n441_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1351gat));
  NOR3_X1   g733(.A1(new_n573_), .A2(new_n469_), .A3(new_n523_), .ZN(new_n935_));
  OAI211_X1 g734(.A(new_n638_), .B(new_n935_), .C1(new_n864_), .C2(new_n866_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n936_), .A2(new_n653_), .ZN(new_n937_));
  XOR2_X1   g736(.A(new_n937_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g737(.A1(new_n936_), .A2(new_n735_), .ZN(new_n939_));
  XOR2_X1   g738(.A(new_n939_), .B(G204gat), .Z(G1353gat));
  AOI21_X1  g739(.A(new_n345_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n941_));
  XOR2_X1   g740(.A(new_n941_), .B(KEYINPUT126), .Z(new_n942_));
  NOR2_X1   g741(.A1(new_n936_), .A2(new_n942_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n943_), .B(new_n944_), .ZN(G1354gat));
  INV_X1    g744(.A(G218gat), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n936_), .A2(new_n946_), .A3(new_n697_), .ZN(new_n947_));
  NOR3_X1   g746(.A1(new_n936_), .A2(KEYINPUT127), .A3(new_n650_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n948_), .A2(G218gat), .ZN(new_n949_));
  OAI21_X1  g748(.A(KEYINPUT127), .B1(new_n936_), .B2(new_n650_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n947_), .B1(new_n949_), .B2(new_n950_), .ZN(G1355gat));
endmodule


