//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 0 0 0 0 1 0 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n899_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n929_, new_n930_,
    new_n932_, new_n933_, new_n934_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_, new_n951_;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G29gat), .B(G36gat), .ZN(new_n203_));
  AND2_X1   g002(.A1(new_n203_), .A2(KEYINPUT68), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(KEYINPUT68), .ZN(new_n205_));
  XOR2_X1   g004(.A(G43gat), .B(G50gat), .Z(new_n206_));
  OR3_X1    g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n206_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n208_));
  AND2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G15gat), .B(G22gat), .ZN(new_n210_));
  INV_X1    g009(.A(G1gat), .ZN(new_n211_));
  INV_X1    g010(.A(G8gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT14), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G1gat), .B(G8gat), .ZN(new_n215_));
  XOR2_X1   g014(.A(new_n214_), .B(new_n215_), .Z(new_n216_));
  NAND2_X1  g015(.A1(new_n209_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n216_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n207_), .A2(new_n208_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n202_), .B1(new_n217_), .B2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n209_), .A2(KEYINPUT15), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT15), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n219_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(new_n218_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n202_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n227_), .B1(new_n209_), .B2(new_n216_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n221_), .B1(new_n226_), .B2(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n229_), .A2(KEYINPUT84), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G113gat), .B(G141gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G169gat), .B(G197gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(KEYINPUT82), .B(KEYINPUT83), .Z(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n230_), .B(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G169gat), .A2(G176gat), .ZN(new_n238_));
  INV_X1    g037(.A(G176gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT22), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT89), .B1(new_n240_), .B2(G169gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT22), .B(G169gat), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n239_), .B(new_n241_), .C1(new_n242_), .C2(KEYINPUT89), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT23), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n244_), .A2(G183gat), .A3(G190gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT90), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n244_), .B1(G183gat), .B2(G190gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(KEYINPUT85), .B(G183gat), .Z(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT87), .B(G190gat), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n238_), .B(new_n243_), .C1(new_n248_), .C2(new_n251_), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n249_), .A2(KEYINPUT86), .A3(KEYINPUT25), .ZN(new_n253_));
  AOI21_X1  g052(.A(KEYINPUT86), .B1(new_n249_), .B2(KEYINPUT25), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT26), .ZN(new_n256_));
  INV_X1    g055(.A(G190gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n258_), .B1(new_n250_), .B2(new_n256_), .ZN(new_n259_));
  INV_X1    g058(.A(G183gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n259_), .B1(KEYINPUT25), .B2(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n255_), .A2(new_n261_), .ZN(new_n262_));
  NOR3_X1   g061(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT23), .B1(new_n260_), .B2(new_n257_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n263_), .B1(new_n264_), .B2(new_n245_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT88), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n266_), .ZN(new_n268_));
  INV_X1    g067(.A(G169gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(new_n239_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n270_), .A2(KEYINPUT24), .A3(new_n238_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n267_), .A2(new_n268_), .A3(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n252_), .B1(new_n262_), .B2(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(G71gat), .B(G99gat), .Z(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT91), .B(G43gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n273_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n273_), .A2(new_n276_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G227gat), .A2(G233gat), .ZN(new_n279_));
  INV_X1    g078(.A(G15gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT30), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT31), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n277_), .A2(new_n278_), .A3(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n283_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT92), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n286_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT92), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(new_n289_), .A3(new_n284_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(G127gat), .B(G134gat), .Z(new_n292_));
  XOR2_X1   g091(.A(G113gat), .B(G120gat), .Z(new_n293_));
  XOR2_X1   g092(.A(new_n292_), .B(new_n293_), .Z(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n291_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n287_), .A2(new_n290_), .A3(new_n294_), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n296_), .A2(KEYINPUT93), .A3(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT93), .B1(new_n296_), .B2(new_n297_), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(G211gat), .B(G218gat), .Z(new_n301_));
  INV_X1    g100(.A(KEYINPUT21), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G197gat), .B(G204gat), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n301_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n303_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT21), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n305_), .A2(new_n301_), .A3(KEYINPUT21), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(G141gat), .ZN(new_n311_));
  INV_X1    g110(.A(G148gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G141gat), .A2(G148gat), .ZN(new_n314_));
  NAND3_X1  g113(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(G155gat), .B(G162gat), .Z(new_n317_));
  INV_X1    g116(.A(KEYINPUT1), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n316_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n314_), .B(KEYINPUT2), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT94), .ZN(new_n321_));
  OR4_X1    g120(.A1(new_n321_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT3), .B1(new_n313_), .B2(new_n321_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n320_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(new_n317_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n319_), .B1(new_n325_), .B2(KEYINPUT95), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT95), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n324_), .A2(new_n327_), .A3(new_n317_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n310_), .B1(new_n329_), .B2(KEYINPUT29), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G228gat), .A2(G233gat), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n331_), .B(KEYINPUT97), .Z(new_n332_));
  OR2_X1    g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G78gat), .B(G106gat), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n330_), .B1(KEYINPUT97), .B2(new_n331_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n333_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n330_), .A2(new_n332_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n331_), .A2(KEYINPUT97), .ZN(new_n339_));
  AOI211_X1 g138(.A(new_n339_), .B(new_n310_), .C1(new_n329_), .C2(KEYINPUT29), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n334_), .B1(new_n338_), .B2(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT28), .B1(new_n329_), .B2(KEYINPUT29), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT28), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT29), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n326_), .A2(new_n343_), .A3(new_n344_), .A4(new_n328_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G22gat), .B(G50gat), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n342_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n342_), .A2(new_n345_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n346_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n337_), .A2(new_n341_), .A3(new_n347_), .A4(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT96), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n342_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n346_), .B1(new_n342_), .B2(new_n345_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n353_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n350_), .A2(KEYINPUT96), .A3(new_n347_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT98), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n337_), .A2(new_n341_), .A3(new_n359_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n333_), .A2(new_n336_), .A3(KEYINPUT98), .A4(new_n335_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n358_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT99), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT99), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n358_), .A2(new_n360_), .A3(new_n364_), .A4(new_n361_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n352_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n326_), .A2(new_n328_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(new_n295_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n329_), .A2(new_n294_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G225gat), .A2(G233gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT4), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n329_), .A2(new_n374_), .A3(new_n294_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n372_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n375_), .B(new_n376_), .C1(new_n370_), .C2(new_n374_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G1gat), .B(G29gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(G85gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT0), .B(G57gat), .ZN(new_n380_));
  XOR2_X1   g179(.A(new_n379_), .B(new_n380_), .Z(new_n381_));
  AND3_X1   g180(.A1(new_n373_), .A2(new_n377_), .A3(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n381_), .B1(new_n373_), .B2(new_n377_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n242_), .A2(new_n239_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(new_n238_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT102), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n264_), .A2(new_n245_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n389_), .B1(G183gat), .B2(G190gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n263_), .ZN(new_n392_));
  XOR2_X1   g191(.A(KEYINPUT26), .B(G190gat), .Z(new_n393_));
  XOR2_X1   g192(.A(KEYINPUT25), .B(G183gat), .Z(new_n394_));
  OAI211_X1 g193(.A(new_n392_), .B(new_n271_), .C1(new_n393_), .C2(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n248_), .A2(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n396_), .A2(KEYINPUT101), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT101), .ZN(new_n398_));
  NOR3_X1   g197(.A1(new_n248_), .A2(new_n395_), .A3(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n391_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n309_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n310_), .B(new_n252_), .C1(new_n262_), .C2(new_n272_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(KEYINPUT20), .A3(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT100), .B(KEYINPUT19), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G226gat), .A2(G233gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n403_), .A2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G8gat), .B(G36gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT18), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G64gat), .B(G92gat), .ZN(new_n411_));
  XOR2_X1   g210(.A(new_n410_), .B(new_n411_), .Z(new_n412_));
  NAND2_X1  g211(.A1(new_n273_), .A2(new_n309_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n391_), .B(new_n310_), .C1(new_n397_), .C2(new_n399_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT20), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n407_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n413_), .A2(new_n414_), .A3(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n408_), .A2(new_n412_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n412_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n415_), .B1(new_n400_), .B2(new_n309_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n406_), .B1(new_n420_), .B2(new_n402_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n417_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n419_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n418_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT27), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n413_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n391_), .ZN(new_n428_));
  OR2_X1    g227(.A1(new_n309_), .A2(new_n396_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT20), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n407_), .B1(new_n427_), .B2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n431_), .B1(new_n403_), .B2(new_n407_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n419_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n433_), .A2(KEYINPUT27), .A3(new_n418_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n426_), .A2(new_n434_), .ZN(new_n435_));
  NOR3_X1   g234(.A1(new_n366_), .A2(new_n385_), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n381_), .B1(new_n371_), .B2(new_n376_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n375_), .B1(new_n370_), .B2(new_n374_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n437_), .B1(new_n376_), .B2(new_n438_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n373_), .A2(new_n377_), .A3(KEYINPUT33), .A4(new_n381_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n439_), .A2(new_n440_), .A3(new_n418_), .A4(new_n423_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n382_), .A2(KEYINPUT33), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n412_), .A2(KEYINPUT32), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n432_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n408_), .A2(new_n417_), .A3(new_n443_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  OAI22_X1  g246(.A1(new_n441_), .A2(new_n442_), .B1(new_n384_), .B2(new_n447_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n366_), .A2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n300_), .B1(new_n436_), .B2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n385_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n435_), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n451_), .A2(new_n366_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n237_), .B1(new_n450_), .B2(new_n454_), .ZN(new_n455_));
  OR2_X1    g254(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n456_));
  INV_X1    g255(.A(G106gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT64), .B(G85gat), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT9), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(G92gat), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n459_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G99gat), .A2(G106gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT6), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT6), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(G99gat), .A3(G106gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  OR2_X1    g267(.A1(G85gat), .A2(G92gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G85gat), .A2(G92gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n468_), .B1(new_n471_), .B2(new_n461_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n463_), .A2(new_n472_), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n469_), .A2(new_n470_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n466_), .B1(G99gat), .B2(G106gat), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n464_), .A2(KEYINPUT6), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT7), .ZN(new_n478_));
  INV_X1    g277(.A(G99gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n478_), .A2(new_n479_), .A3(new_n457_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n474_), .B1(new_n477_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT8), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n481_), .B(new_n480_), .C1(new_n475_), .C2(new_n476_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT8), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n486_), .A3(new_n474_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n473_), .B1(new_n484_), .B2(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n488_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n460_), .A2(new_n462_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n474_), .A2(KEYINPUT9), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n468_), .A4(new_n459_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n481_), .ZN(new_n493_));
  NOR3_X1   g292(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  AOI211_X1 g294(.A(KEYINPUT8), .B(new_n471_), .C1(new_n495_), .C2(new_n468_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n486_), .B1(new_n485_), .B2(new_n474_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n492_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G232gat), .A2(G233gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT34), .ZN(new_n500_));
  OAI22_X1  g299(.A1(new_n498_), .A2(new_n219_), .B1(KEYINPUT35), .B2(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n489_), .A2(new_n501_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n500_), .A2(KEYINPUT35), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT69), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n503_), .B1(new_n501_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n501_), .A2(new_n504_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n507_), .B(new_n503_), .C1(new_n501_), .C2(new_n489_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G190gat), .B(G218gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G134gat), .B(G162gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(new_n512_), .B(KEYINPUT36), .Z(new_n513_));
  XOR2_X1   g312(.A(new_n513_), .B(KEYINPUT71), .Z(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n509_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT72), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n512_), .A2(KEYINPUT36), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n518_), .B(KEYINPUT70), .Z(new_n519_));
  NAND3_X1  g318(.A1(new_n506_), .A2(new_n508_), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n514_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT72), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n517_), .A2(new_n520_), .A3(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n516_), .A2(new_n520_), .A3(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT74), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT74), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n516_), .A2(new_n528_), .A3(new_n520_), .A4(new_n525_), .ZN(new_n529_));
  AOI22_X1  g328(.A1(KEYINPUT37), .A2(new_n524_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(G127gat), .B(G155gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(G183gat), .B(G211gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT79), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT79), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n535_), .A2(new_n538_), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n537_), .A2(KEYINPUT17), .A3(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(KEYINPUT17), .B1(new_n537_), .B2(new_n539_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT75), .ZN(new_n543_));
  INV_X1    g342(.A(G64gat), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(G57gat), .ZN(new_n545_));
  INV_X1    g344(.A(G57gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(G64gat), .ZN(new_n547_));
  AOI21_X1  g346(.A(KEYINPUT11), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G71gat), .B(G78gat), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT65), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  AND2_X1   g349(.A1(G71gat), .A2(G78gat), .ZN(new_n551_));
  NOR2_X1   g350(.A1(G71gat), .A2(G78gat), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT65), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G57gat), .B(G64gat), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n553_), .B(new_n554_), .C1(new_n555_), .C2(KEYINPUT11), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(KEYINPUT11), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n550_), .A2(new_n556_), .A3(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n558_), .B1(new_n550_), .B2(new_n556_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(G231gat), .ZN(new_n562_));
  INV_X1    g361(.A(G233gat), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  OAI22_X1  g364(.A1(new_n559_), .A2(new_n560_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n543_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n565_), .A2(new_n566_), .A3(new_n543_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(new_n569_), .A3(new_n216_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n569_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n218_), .B1(new_n571_), .B2(new_n567_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n542_), .A2(new_n570_), .A3(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT80), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n542_), .A2(KEYINPUT80), .A3(new_n570_), .A4(new_n572_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n572_), .A2(new_n570_), .A3(KEYINPUT76), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(KEYINPUT76), .B1(new_n572_), .B2(new_n570_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT78), .B(KEYINPUT17), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n536_), .A2(new_n581_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n579_), .A2(new_n580_), .A3(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT81), .B1(new_n577_), .B2(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n580_), .A2(new_n582_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n578_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT81), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n586_), .A2(new_n587_), .A3(new_n575_), .A4(new_n576_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n584_), .A2(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(KEYINPUT12), .B1(new_n561_), .B2(new_n488_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT11), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n546_), .A2(G64gat), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n544_), .A2(G57gat), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n591_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n554_), .B1(new_n594_), .B2(new_n553_), .ZN(new_n595_));
  NOR3_X1   g394(.A1(new_n548_), .A2(KEYINPUT65), .A3(new_n549_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n557_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n550_), .A2(new_n556_), .A3(new_n558_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT12), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n599_), .A2(new_n600_), .A3(new_n498_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n590_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G230gat), .A2(G233gat), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n603_), .B1(new_n599_), .B2(new_n498_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT66), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  OAI211_X1 g405(.A(KEYINPUT66), .B(new_n603_), .C1(new_n599_), .C2(new_n498_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n602_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n603_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n561_), .A2(new_n488_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n561_), .A2(new_n488_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n609_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n608_), .A2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G120gat), .B(G148gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT5), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G176gat), .B(G204gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n614_), .A2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(KEYINPUT67), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n619_), .B1(new_n614_), .B2(new_n620_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n621_), .A2(KEYINPUT13), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(KEYINPUT13), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n530_), .A2(new_n589_), .A3(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n455_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n385_), .A2(new_n211_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT38), .ZN(new_n628_));
  OAI22_X1  g427(.A1(new_n626_), .A2(new_n627_), .B1(KEYINPUT105), .B2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(KEYINPUT105), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n629_), .B(new_n630_), .Z(new_n631_));
  NAND2_X1  g430(.A1(new_n516_), .A2(new_n520_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT103), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT103), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n516_), .A2(new_n634_), .A3(new_n520_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n636_), .B1(new_n450_), .B2(new_n454_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n577_), .A2(new_n583_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n624_), .A2(new_n639_), .A3(new_n237_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n637_), .A2(new_n640_), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n641_), .A2(KEYINPUT104), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(KEYINPUT104), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n384_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n631_), .B1(new_n211_), .B2(new_n644_), .ZN(G1324gat));
  NAND3_X1  g444(.A1(new_n637_), .A2(new_n435_), .A3(new_n640_), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n646_), .A2(KEYINPUT106), .A3(G8gat), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT106), .B1(new_n646_), .B2(G8gat), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT39), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n647_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n649_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n626_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(new_n212_), .A3(new_n435_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT40), .ZN(new_n655_));
  OR3_X1    g454(.A1(new_n650_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n655_), .B1(new_n650_), .B2(new_n654_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1325gat));
  NOR2_X1   g457(.A1(new_n298_), .A2(new_n299_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n652_), .A2(new_n280_), .A3(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n642_), .A2(new_n643_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n280_), .B1(new_n661_), .B2(new_n659_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n662_), .A2(KEYINPUT41), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(KEYINPUT41), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n660_), .B1(new_n663_), .B2(new_n664_), .ZN(G1326gat));
  INV_X1    g464(.A(G22gat), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n363_), .A2(new_n365_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(new_n351_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n652_), .A2(new_n666_), .A3(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n366_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n670_), .A2(new_n666_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT42), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n670_), .A2(KEYINPUT42), .A3(new_n666_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n669_), .B1(new_n673_), .B2(new_n674_), .ZN(G1327gat));
  INV_X1    g474(.A(new_n589_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n636_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n676_), .A2(new_n677_), .A3(new_n624_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n455_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(G29gat), .B1(new_n680_), .B2(new_n385_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n682_), .A2(KEYINPUT108), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n668_), .A2(new_n384_), .A3(new_n452_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n366_), .A2(new_n448_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n659_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n530_), .B(new_n684_), .C1(new_n687_), .C2(new_n453_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n530_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(new_n450_), .B2(new_n454_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n688_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n676_), .A2(new_n237_), .A3(new_n624_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT107), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(KEYINPUT109), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n697_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n692_), .A2(new_n699_), .A3(new_n694_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n385_), .A2(G29gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n681_), .B1(new_n701_), .B2(new_n702_), .ZN(G1328gat));
  INV_X1    g502(.A(G36gat), .ZN(new_n704_));
  AND4_X1   g503(.A1(new_n704_), .A2(new_n455_), .A3(new_n435_), .A4(new_n678_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT45), .Z(new_n706_));
  AOI21_X1  g505(.A(new_n452_), .B1(new_n698_), .B2(new_n700_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n706_), .B1(new_n707_), .B2(new_n704_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT46), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n706_), .B(KEYINPUT46), .C1(new_n707_), .C2(new_n704_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1329gat));
  XNOR2_X1  g511(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n296_), .A2(new_n297_), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n692_), .A2(new_n699_), .A3(new_n694_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n699_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n714_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(G43gat), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n679_), .A2(G43gat), .A3(new_n300_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n713_), .B1(new_n718_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n713_), .ZN(new_n722_));
  AOI211_X1 g521(.A(new_n719_), .B(new_n722_), .C1(new_n717_), .C2(G43gat), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n721_), .A2(new_n723_), .ZN(G1330gat));
  AOI21_X1  g523(.A(new_n366_), .B1(new_n698_), .B2(new_n700_), .ZN(new_n725_));
  INV_X1    g524(.A(G50gat), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n668_), .A2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT111), .ZN(new_n728_));
  OAI22_X1  g527(.A1(new_n725_), .A2(new_n726_), .B1(new_n679_), .B2(new_n728_), .ZN(G1331gat));
  NAND2_X1  g528(.A1(new_n624_), .A2(new_n237_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n730_), .B1(new_n450_), .B2(new_n454_), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n731_), .A2(new_n676_), .A3(new_n689_), .ZN(new_n732_));
  AOI21_X1  g531(.A(G57gat), .B1(new_n732_), .B2(new_n385_), .ZN(new_n733_));
  AND4_X1   g532(.A1(new_n637_), .A2(new_n237_), .A3(new_n624_), .A4(new_n676_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n546_), .B1(new_n385_), .B2(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n736_), .B1(new_n735_), .B2(new_n546_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n733_), .B1(new_n734_), .B2(new_n737_), .ZN(G1332gat));
  NAND3_X1  g537(.A1(new_n732_), .A2(new_n544_), .A3(new_n435_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT48), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n734_), .A2(new_n435_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n741_), .B2(G64gat), .ZN(new_n742_));
  AOI211_X1 g541(.A(KEYINPUT48), .B(new_n544_), .C1(new_n734_), .C2(new_n435_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n739_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT113), .ZN(G1333gat));
  INV_X1    g544(.A(G71gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n746_), .B1(new_n734_), .B2(new_n659_), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n747_), .B(KEYINPUT49), .Z(new_n748_));
  NAND3_X1  g547(.A1(new_n732_), .A2(new_n746_), .A3(new_n659_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1334gat));
  INV_X1    g549(.A(G78gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n732_), .A2(new_n751_), .A3(new_n668_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n734_), .B2(new_n668_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n753_), .A2(new_n754_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n752_), .B1(new_n755_), .B2(new_n756_), .ZN(G1335gat));
  NOR2_X1   g556(.A1(new_n676_), .A2(new_n677_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n731_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n385_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n730_), .A2(new_n676_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n692_), .A2(new_n762_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n384_), .A2(new_n460_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n761_), .B1(new_n763_), .B2(new_n764_), .ZN(G1336gat));
  INV_X1    g564(.A(G92gat), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n760_), .A2(new_n766_), .A3(new_n435_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n763_), .A2(new_n435_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(new_n766_), .ZN(G1337gat));
  AND4_X1   g568(.A1(new_n714_), .A2(new_n760_), .A3(new_n456_), .A4(new_n458_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n763_), .A2(new_n659_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(G99gat), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n772_), .B(new_n773_), .ZN(G1338gat));
  NAND3_X1  g573(.A1(new_n760_), .A2(new_n457_), .A3(new_n668_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n692_), .A2(new_n668_), .A3(new_n762_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n776_), .A2(new_n777_), .A3(G106gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n776_), .B2(G106gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g580(.A1(new_n668_), .A2(new_n435_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n384_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT118), .ZN(new_n785_));
  XOR2_X1   g584(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n786_));
  AND3_X1   g585(.A1(new_n608_), .A2(new_n785_), .A3(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n785_), .B1(new_n608_), .B2(new_n786_), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n599_), .A2(new_n600_), .A3(new_n498_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n600_), .B1(new_n599_), .B2(new_n498_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n610_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n609_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n602_), .A2(new_n606_), .A3(KEYINPUT55), .A4(new_n607_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n787_), .A2(new_n788_), .A3(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT56), .B1(new_n795_), .B2(new_n620_), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n226_), .A2(new_n217_), .A3(new_n227_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n227_), .B1(new_n217_), .B2(new_n220_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n235_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n799_), .B1(new_n229_), .B2(new_n235_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n608_), .A2(new_n786_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT118), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n792_), .A2(new_n793_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n608_), .A2(new_n785_), .A3(new_n786_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n802_), .A2(new_n803_), .A3(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT56), .ZN(new_n806_));
  INV_X1    g605(.A(new_n620_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n805_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n796_), .A2(new_n619_), .A3(new_n800_), .A4(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT58), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n805_), .A2(new_n807_), .ZN(new_n812_));
  AOI22_X1  g611(.A1(new_n812_), .A2(KEYINPUT56), .B1(new_n614_), .B2(new_n618_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n813_), .A2(KEYINPUT58), .A3(new_n800_), .A4(new_n808_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n530_), .A2(new_n811_), .A3(new_n814_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n796_), .A2(new_n236_), .A3(new_n619_), .A4(new_n808_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n800_), .A2(new_n621_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n636_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n818_), .A2(new_n819_), .A3(KEYINPUT57), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n818_), .B2(KEYINPUT57), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n815_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n816_), .A2(new_n817_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n677_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n824_), .A2(KEYINPUT119), .A3(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT119), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n818_), .B2(KEYINPUT57), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n639_), .B1(new_n822_), .B2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n584_), .A2(new_n588_), .A3(new_n237_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n527_), .A2(new_n529_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n524_), .A2(KEYINPUT37), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n834_), .A2(new_n835_), .B1(new_n623_), .B2(new_n622_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n584_), .A2(new_n588_), .A3(KEYINPUT115), .A4(new_n237_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n833_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n833_), .A2(new_n836_), .A3(new_n837_), .A4(new_n839_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n784_), .B1(new_n830_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n841_), .A2(new_n842_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n824_), .A2(new_n825_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n815_), .B(new_n847_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n846_), .B1(new_n589_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n784_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n845_), .ZN(new_n851_));
  OAI22_X1  g650(.A1(new_n844_), .A2(new_n845_), .B1(new_n849_), .B2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(G113gat), .B1(new_n852_), .B2(new_n237_), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n811_), .A2(new_n530_), .A3(new_n814_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n823_), .A2(KEYINPUT57), .A3(new_n677_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT120), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n818_), .A2(new_n819_), .A3(KEYINPUT57), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n854_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(KEYINPUT119), .B1(new_n824_), .B2(new_n825_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n818_), .A2(new_n827_), .A3(KEYINPUT57), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n638_), .B1(new_n858_), .B2(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n850_), .B1(new_n862_), .B2(new_n846_), .ZN(new_n863_));
  OR2_X1    g662(.A1(new_n237_), .A2(G113gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n853_), .B1(new_n863_), .B2(new_n864_), .ZN(G1340gat));
  XOR2_X1   g664(.A(KEYINPUT121), .B(G120gat), .Z(new_n866_));
  NAND2_X1  g665(.A1(new_n848_), .A2(new_n589_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n851_), .B1(new_n867_), .B2(new_n843_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n868_), .B1(new_n863_), .B2(KEYINPUT59), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n866_), .B1(new_n869_), .B2(new_n624_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n624_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n866_), .B1(new_n871_), .B2(KEYINPUT60), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(KEYINPUT60), .B2(new_n866_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n863_), .A2(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(KEYINPUT122), .B1(new_n870_), .B2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n866_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n852_), .B2(new_n871_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n878_));
  INV_X1    g677(.A(new_n874_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n877_), .A2(new_n878_), .A3(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n875_), .A2(new_n880_), .ZN(G1341gat));
  OAI21_X1  g680(.A(G127gat), .B1(new_n852_), .B2(new_n639_), .ZN(new_n882_));
  OR2_X1    g681(.A1(new_n589_), .A2(G127gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n863_), .B2(new_n883_), .ZN(G1342gat));
  INV_X1    g683(.A(G134gat), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n885_), .B1(new_n869_), .B2(new_n530_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n863_), .A2(G134gat), .A3(new_n677_), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT123), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(G134gat), .B1(new_n852_), .B2(new_n689_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT123), .ZN(new_n890_));
  INV_X1    g689(.A(new_n887_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n889_), .A2(new_n890_), .A3(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n888_), .A2(new_n892_), .ZN(G1343gat));
  NAND2_X1  g692(.A1(new_n830_), .A2(new_n843_), .ZN(new_n894_));
  NOR4_X1   g693(.A1(new_n659_), .A2(new_n384_), .A3(new_n366_), .A4(new_n435_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n237_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(new_n311_), .ZN(G1344gat));
  NOR2_X1   g697(.A1(new_n896_), .A2(new_n871_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n312_), .ZN(G1345gat));
  NOR2_X1   g699(.A1(new_n896_), .A2(new_n589_), .ZN(new_n901_));
  XOR2_X1   g700(.A(KEYINPUT61), .B(G155gat), .Z(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1346gat));
  INV_X1    g702(.A(G162gat), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n896_), .A2(new_n904_), .A3(new_n689_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n896_), .B2(new_n677_), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n906_), .A2(KEYINPUT124), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(KEYINPUT124), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n905_), .B1(new_n907_), .B2(new_n908_), .ZN(G1347gat));
  INV_X1    g708(.A(KEYINPUT62), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n452_), .A2(new_n385_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n659_), .A2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n366_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n849_), .A2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(new_n237_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n910_), .B1(new_n917_), .B2(new_n269_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n242_), .ZN(new_n919_));
  OAI211_X1 g718(.A(KEYINPUT62), .B(G169gat), .C1(new_n916_), .C2(new_n237_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n918_), .A2(new_n919_), .A3(new_n920_), .ZN(G1348gat));
  AOI21_X1  g720(.A(G176gat), .B1(new_n915_), .B2(new_n624_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n668_), .B1(new_n830_), .B2(new_n843_), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n912_), .A2(new_n239_), .A3(new_n871_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n922_), .B1(new_n923_), .B2(new_n924_), .ZN(G1349gat));
  NAND3_X1  g724(.A1(new_n923_), .A2(new_n676_), .A3(new_n913_), .ZN(new_n926_));
  AND2_X1   g725(.A1(new_n638_), .A2(new_n394_), .ZN(new_n927_));
  AOI22_X1  g726(.A1(new_n926_), .A2(new_n249_), .B1(new_n915_), .B2(new_n927_), .ZN(G1350gat));
  OAI21_X1  g727(.A(G190gat), .B1(new_n916_), .B2(new_n689_), .ZN(new_n929_));
  OR2_X1    g728(.A1(new_n677_), .A2(new_n393_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n916_), .B2(new_n930_), .ZN(G1351gat));
  NOR4_X1   g730(.A1(new_n659_), .A2(new_n385_), .A3(new_n366_), .A4(new_n452_), .ZN(new_n932_));
  AND2_X1   g731(.A1(new_n894_), .A2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(new_n236_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g734(.A1(new_n894_), .A2(new_n932_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n936_), .A2(new_n871_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(new_n938_), .ZN(new_n939_));
  XOR2_X1   g738(.A(KEYINPUT125), .B(G204gat), .Z(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n937_), .B2(new_n940_), .ZN(G1353gat));
  XNOR2_X1  g740(.A(KEYINPUT63), .B(G211gat), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n933_), .A2(new_n638_), .A3(new_n942_), .ZN(new_n943_));
  OAI22_X1  g742(.A1(new_n936_), .A2(new_n639_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT126), .ZN(new_n945_));
  AND3_X1   g744(.A1(new_n943_), .A2(new_n944_), .A3(new_n945_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n945_), .B1(new_n943_), .B2(new_n944_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n946_), .A2(new_n947_), .ZN(G1354gat));
  XNOR2_X1  g747(.A(KEYINPUT127), .B(G218gat), .ZN(new_n949_));
  NOR3_X1   g748(.A1(new_n936_), .A2(new_n689_), .A3(new_n949_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n933_), .A2(new_n636_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n950_), .B1(new_n951_), .B2(new_n949_), .ZN(G1355gat));
endmodule


