//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n773_, new_n774_, new_n775_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n798_, new_n799_, new_n800_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n813_, new_n814_,
    new_n815_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n931_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n961_, new_n962_,
    new_n963_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n989_, new_n990_,
    new_n992_, new_n993_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1007_, new_n1008_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G43gat), .B(G50gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT73), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n204_), .A2(KEYINPUT73), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n203_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n207_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(new_n205_), .A3(new_n202_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT15), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT79), .B(G8gat), .ZN(new_n214_));
  INV_X1    g013(.A(G1gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT14), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G15gat), .B(G22gat), .ZN(new_n217_));
  OR2_X1    g016(.A1(G1gat), .A2(G8gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G1gat), .A2(G8gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT80), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT80), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n218_), .A2(new_n222_), .A3(new_n219_), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n216_), .A2(new_n217_), .A3(new_n221_), .A4(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  AOI22_X1  g024(.A1(new_n216_), .A2(new_n217_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n208_), .A2(new_n210_), .A3(KEYINPUT15), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n213_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G229gat), .A2(G233gat), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n211_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n229_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n226_), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n233_), .A2(new_n210_), .A3(new_n208_), .A4(new_n224_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n231_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n230_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G113gat), .B(G141gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G169gat), .B(G197gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n232_), .A2(new_n237_), .A3(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n241_), .B1(new_n232_), .B2(new_n237_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT72), .ZN(new_n245_));
  AND3_X1   g044(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n246_));
  AOI21_X1  g045(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT10), .B(G99gat), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n248_), .B1(G106gat), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  OR2_X1    g050(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n252_));
  INV_X1    g051(.A(G85gat), .ZN(new_n253_));
  INV_X1    g052(.A(G92gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n252_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  OR2_X1    g056(.A1(KEYINPUT66), .A2(G92gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(KEYINPUT66), .A2(G92gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(G85gat), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n253_), .A2(new_n254_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT9), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n251_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(G57gat), .ZN(new_n266_));
  INV_X1    g065(.A(G64gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G57gat), .A2(G64gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT11), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G71gat), .B(G78gat), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT11), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n268_), .A2(new_n274_), .A3(new_n269_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n271_), .A2(new_n273_), .A3(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n270_), .A2(new_n272_), .A3(KEYINPUT11), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT8), .ZN(new_n279_));
  XOR2_X1   g078(.A(G85gat), .B(G92gat), .Z(new_n280_));
  NOR2_X1   g079(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n281_));
  NOR2_X1   g080(.A1(G99gat), .A2(G106gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  AND2_X1   g082(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  OAI22_X1  g084(.A1(KEYINPUT67), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n283_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n247_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n279_), .B(new_n280_), .C1(new_n287_), .C2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n284_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(new_n248_), .A3(new_n286_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n279_), .B1(new_n294_), .B2(new_n280_), .ZN(new_n295_));
  OAI211_X1 g094(.A(new_n265_), .B(new_n278_), .C1(new_n292_), .C2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT69), .B1(new_n292_), .B2(new_n295_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n280_), .B1(new_n287_), .B2(new_n290_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT8), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n300_), .A2(new_n301_), .A3(new_n291_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n298_), .A2(new_n302_), .A3(new_n265_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT12), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n278_), .A2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n297_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n257_), .A2(new_n260_), .B1(KEYINPUT9), .B2(new_n262_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n307_), .A2(new_n250_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n308_), .B1(new_n300_), .B2(new_n291_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n304_), .B1(new_n309_), .B2(new_n278_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT70), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G230gat), .A2(G233gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT64), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n265_), .B1(new_n292_), .B2(new_n295_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n278_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT70), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n316_), .A2(new_n317_), .A3(new_n304_), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n306_), .A2(new_n311_), .A3(new_n313_), .A4(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n313_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n316_), .B1(new_n297_), .B2(KEYINPUT68), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT68), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n296_), .A2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n320_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n319_), .A2(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(G120gat), .B(G148gat), .Z(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(G204gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT5), .B(G176gat), .ZN(new_n328_));
  XOR2_X1   g127(.A(new_n327_), .B(new_n328_), .Z(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n325_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n319_), .A2(new_n324_), .A3(new_n329_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n331_), .A2(KEYINPUT71), .A3(new_n332_), .ZN(new_n333_));
  AOI211_X1 g132(.A(KEYINPUT71), .B(new_n329_), .C1(new_n319_), .C2(new_n324_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n333_), .A2(new_n335_), .A3(KEYINPUT13), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(KEYINPUT13), .B1(new_n333_), .B2(new_n335_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n245_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n333_), .A2(new_n335_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT13), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(KEYINPUT72), .A3(new_n336_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n244_), .B1(new_n339_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G141gat), .A2(G148gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT88), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT2), .ZN(new_n347_));
  OR2_X1    g146(.A1(G141gat), .A2(G148gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT3), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT2), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n345_), .A2(KEYINPUT88), .A3(new_n350_), .ZN(new_n351_));
  OR3_X1    g150(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n347_), .A2(new_n349_), .A3(new_n351_), .A4(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(G155gat), .B(G162gat), .Z(new_n354_));
  NOR2_X1   g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  AND3_X1   g155(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n357_));
  AOI21_X1  g156(.A(KEYINPUT1), .B1(G155gat), .B2(G162gat), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n356_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n348_), .A2(new_n345_), .ZN(new_n360_));
  AOI22_X1  g159(.A1(new_n353_), .A2(new_n354_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(G113gat), .B(G120gat), .Z(new_n362_));
  XNOR2_X1  g161(.A(G127gat), .B(G134gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n361_), .B(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G225gat), .A2(G233gat), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  OR2_X1    g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G1gat), .B(G29gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(G85gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT0), .B(G57gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n353_), .A2(new_n354_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n359_), .A2(new_n360_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(new_n364_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n362_), .A2(new_n363_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n362_), .A2(new_n363_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n361_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n376_), .A2(KEYINPUT4), .A3(new_n380_), .ZN(new_n381_));
  OR3_X1    g180(.A1(new_n361_), .A2(new_n379_), .A3(KEYINPUT4), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n368_), .B(new_n372_), .C1(new_n383_), .C2(new_n366_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n372_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n366_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n365_), .A2(new_n367_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n385_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT105), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n384_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  OAI211_X1 g189(.A(KEYINPUT105), .B(new_n385_), .C1(new_n386_), .C2(new_n387_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT22), .B(G169gat), .ZN(new_n394_));
  INV_X1    g193(.A(G176gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G169gat), .A2(G176gat), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT97), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(KEYINPUT97), .A2(G169gat), .A3(G176gat), .ZN(new_n399_));
  AOI22_X1  g198(.A1(new_n394_), .A2(new_n395_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G183gat), .A2(G190gat), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT23), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n404_));
  INV_X1    g203(.A(G183gat), .ZN(new_n405_));
  INV_X1    g204(.A(G190gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n403_), .A2(new_n404_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT98), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n403_), .A2(new_n407_), .A3(KEYINPUT98), .A4(new_n404_), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n400_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n406_), .A2(KEYINPUT26), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT26), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(G190gat), .ZN(new_n415_));
  AND2_X1   g214(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n416_));
  NOR2_X1   g215(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n417_));
  OAI211_X1 g216(.A(new_n413_), .B(new_n415_), .C1(new_n416_), .C2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT95), .ZN(new_n419_));
  INV_X1    g218(.A(G169gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n395_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n421_), .A2(KEYINPUT24), .A3(new_n396_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n418_), .A2(new_n419_), .A3(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n419_), .B1(new_n418_), .B2(new_n422_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT24), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n426_), .A2(new_n420_), .A3(new_n395_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT96), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n427_), .A2(new_n403_), .A3(KEYINPUT96), .A4(new_n404_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n412_), .B1(new_n425_), .B2(new_n433_), .ZN(new_n434_));
  OR2_X1    g233(.A1(G211gat), .A2(G218gat), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT90), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G211gat), .A2(G218gat), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n435_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  AND2_X1   g237(.A1(G211gat), .A2(G218gat), .ZN(new_n439_));
  NOR2_X1   g238(.A1(G211gat), .A2(G218gat), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT90), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n438_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(G197gat), .ZN(new_n443_));
  AND2_X1   g242(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n444_));
  NOR2_X1   g243(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n443_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT21), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n447_), .B1(G197gat), .B2(G204gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(G197gat), .B1(new_n444_), .B2(new_n445_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n443_), .A2(G204gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n442_), .B(new_n449_), .C1(new_n452_), .C2(KEYINPUT21), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n452_), .A2(KEYINPUT21), .A3(new_n441_), .A4(new_n438_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n434_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT20), .ZN(new_n458_));
  OR3_X1    g257(.A1(new_n420_), .A2(KEYINPUT86), .A3(KEYINPUT22), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT86), .B1(new_n420_), .B2(KEYINPUT22), .ZN(new_n460_));
  AOI21_X1  g259(.A(G176gat), .B1(new_n420_), .B2(KEYINPUT22), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n462_), .A2(new_n396_), .A3(new_n408_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(KEYINPUT84), .A2(G183gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT25), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n413_), .A2(new_n415_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT85), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n422_), .A2(new_n427_), .A3(new_n403_), .A4(new_n404_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n468_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n464_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n455_), .A2(KEYINPUT91), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT91), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n453_), .A2(new_n475_), .A3(new_n454_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n473_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G226gat), .A2(G233gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT19), .ZN(new_n479_));
  NOR3_X1   g278(.A1(new_n458_), .A2(new_n477_), .A3(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT99), .B1(new_n434_), .B2(new_n456_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n473_), .A2(new_n474_), .A3(new_n476_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT99), .ZN(new_n483_));
  NOR3_X1   g282(.A1(new_n432_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n483_), .B(new_n455_), .C1(new_n484_), .C2(new_n412_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n481_), .A2(new_n482_), .A3(KEYINPUT20), .A4(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n479_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n480_), .B1(new_n487_), .B2(KEYINPUT100), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT100), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n486_), .A2(new_n489_), .A3(new_n479_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G8gat), .B(G36gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT102), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n492_), .B(KEYINPUT101), .Z(new_n493_));
  XOR2_X1   g292(.A(G64gat), .B(G92gat), .Z(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT18), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n493_), .B(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT32), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n488_), .A2(new_n490_), .A3(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n479_), .B1(new_n458_), .B2(new_n477_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n500_), .B(KEYINPUT104), .C1(new_n479_), .C2(new_n486_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT104), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n502_), .B(new_n479_), .C1(new_n458_), .C2(new_n477_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n501_), .A2(KEYINPUT32), .A3(new_n497_), .A4(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n393_), .A2(new_n499_), .A3(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n487_), .A2(KEYINPUT100), .ZN(new_n506_));
  INV_X1    g305(.A(new_n480_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(new_n490_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(new_n496_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n488_), .A2(new_n497_), .A3(new_n490_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n383_), .A2(new_n366_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n385_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT103), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n388_), .B(KEYINPUT33), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n505_), .B1(new_n511_), .B2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT28), .B1(new_n375_), .B2(KEYINPUT29), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n375_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G22gat), .B(G50gat), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NOR3_X1   g322(.A1(new_n520_), .A2(new_n521_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n521_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n522_), .B1(new_n525_), .B2(new_n519_), .ZN(new_n526_));
  OR2_X1    g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(G78gat), .B(G106gat), .Z(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(G228gat), .ZN(new_n530_));
  INV_X1    g329(.A(G233gat), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT29), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n533_), .B1(new_n361_), .B2(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n535_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n375_), .A2(KEYINPUT29), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n533_), .B1(new_n537_), .B2(new_n455_), .ZN(new_n538_));
  OAI211_X1 g337(.A(KEYINPUT92), .B(new_n529_), .C1(new_n536_), .C2(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n532_), .B1(new_n375_), .B2(KEYINPUT29), .ZN(new_n540_));
  INV_X1    g339(.A(new_n476_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n475_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n540_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n361_), .A2(new_n534_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n532_), .B1(new_n456_), .B2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(new_n545_), .A3(new_n528_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n539_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n543_), .A2(new_n545_), .ZN(new_n548_));
  AOI21_X1  g347(.A(KEYINPUT92), .B1(new_n548_), .B2(new_n529_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n527_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT93), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n527_), .B(KEYINPUT93), .C1(new_n547_), .C2(new_n549_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n536_), .A2(new_n538_), .ZN(new_n555_));
  OR2_X1    g354(.A1(new_n528_), .A2(KEYINPUT94), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n524_), .A2(new_n526_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n555_), .A2(new_n556_), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n557_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G71gat), .B(G99gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(G43gat), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n473_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n473_), .A2(new_n564_), .ZN(new_n567_));
  INV_X1    g366(.A(G227gat), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n364_), .B1(new_n568_), .B2(new_n531_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n531_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n379_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT30), .B(G15gat), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n573_), .B(KEYINPUT31), .Z(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n574_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n569_), .A2(new_n571_), .A3(new_n576_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n566_), .A2(new_n567_), .A3(new_n575_), .A4(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n575_), .A2(new_n577_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n567_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n579_), .B1(new_n580_), .B2(new_n565_), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n578_), .A2(new_n581_), .A3(KEYINPUT87), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT87), .B1(new_n578_), .B2(new_n581_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n554_), .A2(new_n561_), .A3(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n518_), .A2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n584_), .B1(new_n554_), .B2(new_n561_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n578_), .A2(new_n581_), .ZN(new_n589_));
  AOI211_X1 g388(.A(new_n589_), .B(new_n560_), .C1(new_n552_), .C2(new_n553_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT27), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n508_), .A2(new_n496_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n497_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n592_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n501_), .A2(new_n496_), .A3(new_n503_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n510_), .A2(KEYINPUT27), .A3(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n595_), .A2(new_n392_), .A3(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n587_), .B1(new_n591_), .B2(new_n598_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n344_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n213_), .A2(new_n228_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n300_), .A2(new_n291_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n308_), .B1(new_n602_), .B2(KEYINPUT69), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n601_), .B1(new_n603_), .B2(new_n302_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT35), .ZN(new_n605_));
  NAND2_X1  g404(.A1(G232gat), .A2(G233gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT34), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  AOI22_X1  g407(.A1(new_n309_), .A2(new_n211_), .B1(new_n605_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(KEYINPUT35), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(KEYINPUT77), .B1(new_n604_), .B2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n303_), .A2(new_n228_), .A3(new_n213_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT77), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n613_), .A2(new_n614_), .A3(new_n610_), .A4(new_n609_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n609_), .A2(KEYINPUT74), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n602_), .A2(new_n211_), .A3(new_n265_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n608_), .A2(new_n605_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT74), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n617_), .A2(new_n622_), .A3(new_n613_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n610_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n616_), .A2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G134gat), .B(G162gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT75), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G190gat), .B(G218gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT36), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n626_), .A2(new_n631_), .ZN(new_n632_));
  AOI22_X1  g431(.A1(new_n612_), .A2(new_n615_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n633_));
  XOR2_X1   g432(.A(KEYINPUT76), .B(KEYINPUT36), .Z(new_n634_));
  AND2_X1   g433(.A1(new_n630_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n632_), .A2(KEYINPUT37), .A3(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(KEYINPUT78), .B1(new_n626_), .B2(new_n631_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT78), .ZN(new_n639_));
  INV_X1    g438(.A(new_n631_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n633_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n636_), .B1(new_n638_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT37), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n637_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(G231gat), .A2(G233gat), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n233_), .A2(new_n224_), .A3(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n233_), .B2(new_n224_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n278_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  OAI211_X1 g447(.A(G231gat), .B(G233gat), .C1(new_n225_), .C2(new_n226_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n233_), .A2(new_n224_), .A3(new_n645_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n649_), .A2(new_n315_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT82), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n648_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n654_));
  XNOR2_X1  g453(.A(G127gat), .B(G155gat), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(new_n656_));
  XOR2_X1   g455(.A(G183gat), .B(G211gat), .Z(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(KEYINPUT17), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n653_), .A2(new_n660_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n648_), .A2(new_n652_), .A3(new_n659_), .A4(new_n651_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n648_), .A2(new_n651_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n658_), .A2(KEYINPUT17), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n661_), .A2(new_n662_), .A3(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT83), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n661_), .A2(new_n665_), .A3(KEYINPUT83), .A4(new_n662_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n644_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n600_), .A2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n674_), .A2(new_n215_), .A3(new_n393_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT38), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n626_), .A2(KEYINPUT78), .A3(new_n631_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n639_), .B1(new_n633_), .B2(new_n640_), .ZN(new_n679_));
  AOI22_X1  g478(.A1(new_n678_), .A2(new_n679_), .B1(new_n633_), .B2(new_n635_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n680_), .A2(new_n670_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n600_), .A2(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G1gat), .B1(new_n682_), .B2(new_n392_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n675_), .A2(new_n676_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n677_), .A2(new_n683_), .A3(new_n684_), .ZN(G1324gat));
  AND2_X1   g484(.A1(new_n596_), .A2(KEYINPUT27), .ZN(new_n686_));
  AOI22_X1  g485(.A1(new_n592_), .A2(new_n511_), .B1(new_n686_), .B2(new_n510_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n600_), .A2(new_n214_), .A3(new_n688_), .A4(new_n673_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT106), .ZN(new_n690_));
  OAI21_X1  g489(.A(G8gat), .B1(new_n682_), .B2(new_n687_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n691_), .A2(KEYINPUT39), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(KEYINPUT39), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n690_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT40), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(KEYINPUT40), .B(new_n690_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1325gat));
  OAI21_X1  g497(.A(G15gat), .B1(new_n682_), .B2(new_n585_), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n699_), .A2(KEYINPUT41), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(KEYINPUT41), .ZN(new_n701_));
  INV_X1    g500(.A(G15gat), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n674_), .A2(new_n702_), .A3(new_n584_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n700_), .A2(new_n701_), .A3(new_n703_), .ZN(G1326gat));
  AOI21_X1  g503(.A(new_n560_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n705_));
  OAI21_X1  g504(.A(G22gat), .B1(new_n682_), .B2(new_n705_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT42), .ZN(new_n707_));
  INV_X1    g506(.A(G22gat), .ZN(new_n708_));
  INV_X1    g507(.A(new_n705_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n674_), .A2(new_n708_), .A3(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n707_), .A2(new_n710_), .ZN(G1327gat));
  NOR2_X1   g510(.A1(new_n642_), .A2(new_n671_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n600_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(G29gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n714_), .A2(new_n715_), .A3(new_n393_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n344_), .A2(new_n670_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n589_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT92), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n719_), .B1(new_n555_), .B2(new_n528_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(new_n546_), .A3(new_n539_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT93), .B1(new_n721_), .B2(new_n527_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n553_), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n718_), .B(new_n561_), .C1(new_n722_), .C2(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n724_), .B1(new_n705_), .B2(new_n584_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n725_), .A2(new_n687_), .A3(new_n392_), .ZN(new_n726_));
  AOI211_X1 g525(.A(KEYINPUT43), .B(new_n644_), .C1(new_n726_), .C2(new_n587_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT43), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n632_), .A2(KEYINPUT37), .A3(new_n636_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n729_), .B1(new_n680_), .B2(KEYINPUT37), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n728_), .B1(new_n599_), .B2(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n717_), .B1(new_n727_), .B2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n733_), .A2(KEYINPUT107), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(KEYINPUT107), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n732_), .A2(new_n734_), .A3(new_n735_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n595_), .A2(new_n392_), .A3(new_n597_), .ZN(new_n737_));
  AOI22_X1  g536(.A1(new_n737_), .A2(new_n725_), .B1(new_n518_), .B2(new_n586_), .ZN(new_n738_));
  OAI21_X1  g537(.A(KEYINPUT43), .B1(new_n738_), .B2(new_n644_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n599_), .A2(new_n728_), .A3(new_n730_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n741_), .A2(KEYINPUT107), .A3(new_n733_), .A4(new_n717_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n392_), .B1(new_n736_), .B2(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n716_), .B1(new_n743_), .B2(new_n715_), .ZN(G1328gat));
  INV_X1    g543(.A(KEYINPUT46), .ZN(new_n745_));
  INV_X1    g544(.A(G36gat), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n736_), .A2(new_n742_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n747_), .B2(new_n688_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT45), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n687_), .A2(G36gat), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n344_), .A2(new_n599_), .A3(new_n712_), .A4(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT108), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n751_), .A2(KEYINPUT108), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n749_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n754_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n756_), .A2(KEYINPUT45), .A3(new_n752_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n745_), .B1(new_n748_), .B2(new_n758_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n755_), .A2(new_n757_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n687_), .B1(new_n736_), .B2(new_n742_), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n760_), .B(KEYINPUT46), .C1(new_n761_), .C2(new_n746_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n759_), .A2(new_n762_), .ZN(G1329gat));
  INV_X1    g562(.A(G43gat), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n714_), .A2(new_n764_), .A3(new_n584_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n589_), .B1(new_n736_), .B2(new_n742_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(new_n764_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n765_), .B(new_n768_), .C1(new_n766_), .C2(new_n764_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(G1330gat));
  INV_X1    g571(.A(G50gat), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n714_), .A2(new_n773_), .A3(new_n709_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n705_), .B1(new_n736_), .B2(new_n742_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(new_n773_), .ZN(G1331gat));
  INV_X1    g575(.A(new_n244_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n339_), .A2(new_n343_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n738_), .A2(new_n777_), .A3(new_n778_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n779_), .A2(new_n681_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n266_), .B1(new_n780_), .B2(new_n393_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n673_), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n782_), .A2(G57gat), .A3(new_n392_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  XOR2_X1   g583(.A(new_n784_), .B(KEYINPUT110), .Z(G1332gat));
  NAND2_X1  g584(.A1(new_n779_), .A2(new_n681_), .ZN(new_n786_));
  OAI21_X1  g585(.A(G64gat), .B1(new_n786_), .B2(new_n687_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT48), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n688_), .A2(new_n267_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n788_), .B1(new_n782_), .B2(new_n789_), .ZN(G1333gat));
  INV_X1    g589(.A(G71gat), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n791_), .B1(new_n780_), .B2(new_n584_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(KEYINPUT111), .B(KEYINPUT49), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n792_), .A2(new_n793_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n584_), .A2(new_n791_), .ZN(new_n796_));
  OAI22_X1  g595(.A1(new_n794_), .A2(new_n795_), .B1(new_n782_), .B2(new_n796_), .ZN(G1334gat));
  OAI21_X1  g596(.A(G78gat), .B1(new_n786_), .B2(new_n705_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT50), .ZN(new_n799_));
  OR2_X1    g598(.A1(new_n705_), .A2(G78gat), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n799_), .B1(new_n782_), .B2(new_n800_), .ZN(G1335gat));
  AND2_X1   g600(.A1(new_n779_), .A2(new_n712_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n393_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n253_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n741_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n739_), .A2(KEYINPUT112), .A3(new_n740_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n778_), .A2(new_n777_), .A3(new_n671_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n806_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n393_), .A2(G85gat), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n804_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(KEYINPUT113), .ZN(G1336gat));
  AOI21_X1  g611(.A(G92gat), .B1(new_n802_), .B2(new_n688_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n809_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n688_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n813_), .B1(new_n814_), .B2(new_n815_), .ZN(G1337gat));
  NAND4_X1  g615(.A1(new_n806_), .A2(new_n584_), .A3(new_n807_), .A4(new_n808_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(G99gat), .ZN(new_n818_));
  INV_X1    g617(.A(new_n249_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n802_), .A2(new_n819_), .A3(new_n718_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT51), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n818_), .A2(new_n823_), .A3(new_n820_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(G1338gat));
  NOR2_X1   g624(.A1(new_n705_), .A2(G106gat), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n779_), .A2(new_n712_), .A3(new_n826_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT114), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n741_), .A2(new_n709_), .A3(new_n808_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n829_), .A2(new_n830_), .A3(G106gat), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n830_), .B1(new_n829_), .B2(G106gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n828_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT53), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT53), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n828_), .B(new_n835_), .C1(new_n831_), .C2(new_n832_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(G1339gat));
  NAND2_X1  g636(.A1(new_n777_), .A2(new_n332_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT56), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n306_), .A2(new_n311_), .A3(new_n318_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n320_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n841_), .A2(KEYINPUT55), .A3(new_n319_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n317_), .B1(new_n316_), .B2(new_n304_), .ZN(new_n843_));
  AOI211_X1 g642(.A(KEYINPUT70), .B(KEYINPUT12), .C1(new_n314_), .C2(new_n315_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT55), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n845_), .A2(new_n846_), .A3(new_n313_), .A4(new_n306_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n330_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n839_), .B1(new_n842_), .B2(new_n848_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n847_), .A2(new_n330_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n841_), .A2(KEYINPUT55), .A3(new_n319_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n850_), .A2(KEYINPUT56), .A3(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n838_), .B1(new_n849_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n235_), .A2(new_n230_), .ZN(new_n854_));
  AOI21_X1  g653(.A(KEYINPUT117), .B1(new_n854_), .B2(new_n240_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n229_), .A2(new_n231_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n855_), .B1(new_n236_), .B2(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n854_), .A2(KEYINPUT117), .A3(new_n240_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n242_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  AND3_X1   g658(.A1(new_n333_), .A2(new_n335_), .A3(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n642_), .B1(new_n853_), .B2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  OAI211_X1 g662(.A(KEYINPUT57), .B(new_n642_), .C1(new_n853_), .C2(new_n860_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT118), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n849_), .A2(new_n865_), .A3(new_n852_), .ZN(new_n866_));
  OAI211_X1 g665(.A(KEYINPUT118), .B(new_n839_), .C1(new_n842_), .C2(new_n848_), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n859_), .A2(new_n332_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n866_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(KEYINPUT119), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n730_), .B1(new_n869_), .B2(new_n872_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n868_), .A2(new_n867_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n871_), .B1(new_n874_), .B2(new_n866_), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n863_), .B(new_n864_), .C1(new_n873_), .C2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n670_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n342_), .A2(new_n336_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n668_), .A2(new_n244_), .A3(new_n669_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(KEYINPUT115), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n879_), .B1(new_n883_), .B2(new_n730_), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n644_), .A2(new_n880_), .A3(new_n882_), .A4(new_n878_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n877_), .A2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n687_), .A2(new_n393_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(new_n724_), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n888_), .A2(KEYINPUT120), .A3(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(KEYINPUT120), .B1(new_n888_), .B2(new_n890_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n777_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(G113gat), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n890_), .A2(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n886_), .B1(new_n877_), .B2(KEYINPUT121), .ZN(new_n897_));
  INV_X1    g696(.A(new_n838_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n842_), .A2(new_n839_), .A3(new_n848_), .ZN(new_n899_));
  AOI21_X1  g698(.A(KEYINPUT56), .B1(new_n850_), .B2(new_n851_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n898_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n333_), .A2(new_n335_), .A3(new_n859_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(KEYINPUT57), .B1(new_n903_), .B2(new_n642_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n864_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n869_), .A2(new_n872_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n874_), .A2(new_n871_), .A3(new_n866_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n907_), .A2(new_n908_), .A3(new_n730_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n671_), .B1(new_n906_), .B2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT121), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n896_), .B1(new_n897_), .B2(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n895_), .B1(new_n888_), .B2(new_n890_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n244_), .A2(new_n894_), .ZN(new_n916_));
  AOI22_X1  g715(.A1(new_n893_), .A2(new_n894_), .B1(new_n915_), .B2(new_n916_), .ZN(G1340gat));
  NOR3_X1   g716(.A1(new_n913_), .A2(new_n914_), .A3(new_n778_), .ZN(new_n918_));
  INV_X1    g717(.A(G120gat), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n891_), .A2(new_n892_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n778_), .B2(KEYINPUT60), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n921_), .B1(KEYINPUT60), .B2(new_n919_), .ZN(new_n922_));
  OAI22_X1  g721(.A1(new_n918_), .A2(new_n919_), .B1(new_n920_), .B2(new_n922_), .ZN(G1341gat));
  OAI21_X1  g722(.A(new_n671_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n924_));
  INV_X1    g723(.A(G127gat), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n671_), .A2(G127gat), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(KEYINPUT122), .ZN(new_n927_));
  AOI22_X1  g726(.A1(new_n924_), .A2(new_n925_), .B1(new_n915_), .B2(new_n927_), .ZN(G1342gat));
  OAI21_X1  g727(.A(new_n680_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n929_));
  INV_X1    g728(.A(G134gat), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n644_), .A2(new_n930_), .ZN(new_n931_));
  AOI22_X1  g730(.A1(new_n929_), .A2(new_n930_), .B1(new_n915_), .B2(new_n931_), .ZN(G1343gat));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n933_));
  INV_X1    g732(.A(new_n588_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n934_), .B1(new_n877_), .B2(new_n887_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n889_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n933_), .B1(new_n935_), .B2(new_n936_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n886_), .B1(new_n876_), .B2(new_n670_), .ZN(new_n938_));
  NOR4_X1   g737(.A1(new_n938_), .A2(KEYINPUT123), .A3(new_n934_), .A4(new_n889_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n777_), .B1(new_n937_), .B2(new_n939_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(KEYINPUT124), .B(G141gat), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(new_n942_));
  OAI211_X1 g741(.A(new_n588_), .B(new_n936_), .C1(new_n910_), .C2(new_n886_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(KEYINPUT123), .ZN(new_n944_));
  NAND4_X1  g743(.A1(new_n888_), .A2(new_n933_), .A3(new_n588_), .A4(new_n936_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(new_n946_));
  INV_X1    g745(.A(new_n941_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n946_), .A2(new_n777_), .A3(new_n947_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n942_), .A2(new_n948_), .ZN(G1344gat));
  XNOR2_X1  g748(.A(KEYINPUT125), .B(G148gat), .ZN(new_n950_));
  INV_X1    g749(.A(new_n950_), .ZN(new_n951_));
  INV_X1    g750(.A(new_n778_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n951_), .B1(new_n946_), .B2(new_n952_), .ZN(new_n953_));
  AOI211_X1 g752(.A(new_n778_), .B(new_n950_), .C1(new_n944_), .C2(new_n945_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n953_), .A2(new_n954_), .ZN(G1345gat));
  XNOR2_X1  g754(.A(KEYINPUT61), .B(G155gat), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n956_), .B1(new_n946_), .B2(new_n671_), .ZN(new_n957_));
  INV_X1    g756(.A(new_n956_), .ZN(new_n958_));
  AOI211_X1 g757(.A(new_n670_), .B(new_n958_), .C1(new_n944_), .C2(new_n945_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n957_), .A2(new_n959_), .ZN(G1346gat));
  NAND2_X1  g759(.A1(new_n946_), .A2(new_n680_), .ZN(new_n961_));
  INV_X1    g760(.A(G162gat), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n644_), .A2(new_n962_), .ZN(new_n963_));
  AOI22_X1  g762(.A1(new_n961_), .A2(new_n962_), .B1(new_n946_), .B2(new_n963_), .ZN(G1347gat));
  INV_X1    g763(.A(KEYINPUT62), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n687_), .A2(new_n393_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(new_n709_), .A2(new_n585_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n966_), .A2(new_n967_), .ZN(new_n968_));
  AOI211_X1 g767(.A(new_n244_), .B(new_n968_), .C1(new_n897_), .C2(new_n912_), .ZN(new_n969_));
  OAI21_X1  g768(.A(new_n965_), .B1(new_n969_), .B2(new_n420_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n897_), .A2(new_n912_), .ZN(new_n971_));
  INV_X1    g770(.A(new_n968_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n971_), .A2(new_n972_), .ZN(new_n973_));
  OAI211_X1 g772(.A(KEYINPUT62), .B(G169gat), .C1(new_n973_), .C2(new_n244_), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n969_), .A2(new_n394_), .ZN(new_n975_));
  NAND3_X1  g774(.A1(new_n970_), .A2(new_n974_), .A3(new_n975_), .ZN(G1348gat));
  NAND2_X1  g775(.A1(new_n888_), .A2(new_n972_), .ZN(new_n977_));
  NOR3_X1   g776(.A1(new_n977_), .A2(new_n395_), .A3(new_n778_), .ZN(new_n978_));
  AOI21_X1  g777(.A(new_n968_), .B1(new_n897_), .B2(new_n912_), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n979_), .A2(new_n952_), .ZN(new_n980_));
  AOI21_X1  g779(.A(new_n978_), .B1(new_n980_), .B2(new_n395_), .ZN(G1349gat));
  NOR3_X1   g780(.A1(new_n670_), .A2(new_n417_), .A3(new_n416_), .ZN(new_n982_));
  NAND3_X1  g781(.A1(new_n971_), .A2(new_n972_), .A3(new_n982_), .ZN(new_n983_));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n983_), .A2(new_n984_), .ZN(new_n985_));
  NAND3_X1  g784(.A1(new_n979_), .A2(KEYINPUT126), .A3(new_n982_), .ZN(new_n986_));
  OAI21_X1  g785(.A(new_n405_), .B1(new_n977_), .B2(new_n670_), .ZN(new_n987_));
  AND3_X1   g786(.A1(new_n985_), .A2(new_n986_), .A3(new_n987_), .ZN(G1350gat));
  OAI21_X1  g787(.A(G190gat), .B1(new_n973_), .B2(new_n644_), .ZN(new_n989_));
  NAND3_X1  g788(.A1(new_n680_), .A2(new_n413_), .A3(new_n415_), .ZN(new_n990_));
  OAI21_X1  g789(.A(new_n989_), .B1(new_n973_), .B2(new_n990_), .ZN(G1351gat));
  AND2_X1   g790(.A1(new_n935_), .A2(new_n966_), .ZN(new_n992_));
  NAND2_X1  g791(.A1(new_n992_), .A2(new_n777_), .ZN(new_n993_));
  XNOR2_X1  g792(.A(new_n993_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g793(.A1(new_n935_), .A2(new_n952_), .A3(new_n966_), .ZN(new_n995_));
  NAND2_X1  g794(.A1(new_n995_), .A2(G204gat), .ZN(new_n996_));
  INV_X1    g795(.A(KEYINPUT127), .ZN(new_n997_));
  NAND2_X1  g796(.A1(new_n996_), .A2(new_n997_), .ZN(new_n998_));
  NAND3_X1  g797(.A1(new_n995_), .A2(KEYINPUT127), .A3(G204gat), .ZN(new_n999_));
  NOR2_X1   g798(.A1(new_n444_), .A2(new_n445_), .ZN(new_n1000_));
  OAI211_X1 g799(.A(new_n998_), .B(new_n999_), .C1(new_n1000_), .C2(new_n995_), .ZN(G1353gat));
  NAND3_X1  g800(.A1(new_n935_), .A2(new_n671_), .A3(new_n966_), .ZN(new_n1002_));
  NOR2_X1   g801(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1003_));
  AND2_X1   g802(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1004_));
  NOR3_X1   g803(.A1(new_n1002_), .A2(new_n1003_), .A3(new_n1004_), .ZN(new_n1005_));
  AOI21_X1  g804(.A(new_n1005_), .B1(new_n1002_), .B2(new_n1003_), .ZN(G1354gat));
  AOI21_X1  g805(.A(G218gat), .B1(new_n992_), .B2(new_n680_), .ZN(new_n1007_));
  AND2_X1   g806(.A1(new_n730_), .A2(G218gat), .ZN(new_n1008_));
  AOI21_X1  g807(.A(new_n1007_), .B1(new_n992_), .B2(new_n1008_), .ZN(G1355gat));
endmodule


