//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 1 1 1 0 1 0 1 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n815_, new_n816_, new_n817_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n834_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n853_, new_n855_, new_n856_, new_n857_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  INV_X1    g001(.A(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT0), .B(G57gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  NOR2_X1   g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n210_), .B1(KEYINPUT1), .B2(new_n211_), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n211_), .A2(KEYINPUT1), .ZN(new_n213_));
  AOI211_X1 g012(.A(new_n207_), .B(new_n209_), .C1(new_n212_), .C2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT87), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT84), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n217_), .A2(KEYINPUT3), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n219_), .A2(KEYINPUT84), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n207_), .B1(new_n218_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G141gat), .ZN(new_n222_));
  INV_X1    g021(.A(G148gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n219_), .A2(KEYINPUT84), .ZN(new_n225_));
  NAND2_X1  g024(.A1(KEYINPUT85), .A2(KEYINPUT2), .ZN(new_n226_));
  AOI22_X1  g025(.A1(new_n224_), .A2(new_n225_), .B1(new_n208_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n226_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(KEYINPUT85), .A2(KEYINPUT2), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n209_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n221_), .A2(new_n227_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT86), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT86), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n221_), .A2(new_n227_), .A3(new_n230_), .A4(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n211_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n235_), .A2(new_n210_), .ZN(new_n236_));
  AND4_X1   g035(.A1(new_n216_), .A2(new_n232_), .A3(new_n234_), .A4(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n236_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n238_), .B1(new_n231_), .B2(KEYINPUT86), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n216_), .B1(new_n239_), .B2(new_n234_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n215_), .B1(new_n237_), .B2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G127gat), .B(G134gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G113gat), .B(G120gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n241_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n232_), .A2(new_n234_), .A3(new_n236_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT87), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n239_), .A2(new_n216_), .A3(new_n234_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n250_), .A2(new_n244_), .A3(new_n215_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n246_), .A2(new_n251_), .A3(KEYINPUT4), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n244_), .B1(new_n250_), .B2(new_n215_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT4), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n252_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G225gat), .A2(G233gat), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n258_), .B1(new_n246_), .B2(new_n251_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n206_), .B1(new_n259_), .B2(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n257_), .B1(new_n252_), .B2(new_n255_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n206_), .ZN(new_n264_));
  NOR3_X1   g063(.A1(new_n263_), .A2(new_n264_), .A3(new_n260_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G197gat), .B(G204gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(KEYINPUT88), .A2(KEYINPUT21), .ZN(new_n269_));
  OAI21_X1  g068(.A(G211gat), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(G211gat), .ZN(new_n271_));
  INV_X1    g070(.A(new_n269_), .ZN(new_n272_));
  INV_X1    g071(.A(G204gat), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n273_), .A2(G197gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(G197gat), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n271_), .B(new_n272_), .C1(new_n274_), .C2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n270_), .A2(G218gat), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT21), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n268_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(G218gat), .B1(new_n270_), .B2(new_n276_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n214_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT29), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n282_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(G228gat), .ZN(new_n286_));
  INV_X1    g085(.A(G233gat), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n285_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n241_), .A2(KEYINPUT29), .ZN(new_n290_));
  INV_X1    g089(.A(new_n288_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n290_), .A2(new_n291_), .A3(new_n282_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G78gat), .B(G106gat), .ZN(new_n293_));
  XOR2_X1   g092(.A(new_n293_), .B(KEYINPUT89), .Z(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n289_), .A2(new_n292_), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT91), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n289_), .A2(new_n292_), .A3(KEYINPUT91), .A4(new_n295_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT28), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n283_), .A2(new_n300_), .A3(new_n284_), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n284_), .B(new_n215_), .C1(new_n237_), .C2(new_n240_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT28), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G22gat), .B(G50gat), .ZN(new_n304_));
  AND3_X1   g103(.A1(new_n301_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n304_), .B1(new_n301_), .B2(new_n303_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n291_), .B1(new_n290_), .B2(new_n282_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n281_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n309_), .A2(new_n279_), .A3(new_n277_), .ZN(new_n310_));
  AOI211_X1 g109(.A(new_n288_), .B(new_n310_), .C1(new_n241_), .C2(KEYINPUT29), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n293_), .B1(new_n308_), .B2(new_n311_), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n298_), .A2(new_n299_), .A3(new_n307_), .A4(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n294_), .B1(new_n308_), .B2(new_n311_), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n314_), .A2(KEYINPUT90), .A3(new_n296_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT90), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n289_), .A2(new_n292_), .A3(new_n316_), .A4(new_n295_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n317_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n313_), .B1(new_n315_), .B2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n244_), .B(KEYINPUT82), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G227gat), .A2(G233gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(G15gat), .B(G43gat), .Z(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT22), .B(G169gat), .ZN(new_n325_));
  INV_X1    g124(.A(G176gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G183gat), .A2(G190gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT23), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n330_), .B(new_n331_), .C1(G183gat), .C2(G190gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G169gat), .A2(G176gat), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n327_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT25), .B(G183gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT26), .B(G190gat), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  AOI22_X1  g137(.A1(new_n335_), .A2(new_n336_), .B1(new_n338_), .B2(new_n333_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT24), .ZN(new_n340_));
  INV_X1    g139(.A(G169gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(new_n341_), .A3(new_n326_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT81), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n339_), .A2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n343_), .A2(new_n344_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n334_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  XOR2_X1   g147(.A(KEYINPUT83), .B(KEYINPUT30), .Z(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT31), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n348_), .B(new_n350_), .ZN(new_n351_));
  XOR2_X1   g150(.A(G71gat), .B(G99gat), .Z(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n324_), .B(new_n353_), .ZN(new_n354_));
  NOR3_X1   g153(.A1(new_n267_), .A2(new_n319_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT27), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G226gat), .A2(G233gat), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n357_), .B(KEYINPUT19), .Z(new_n358_));
  INV_X1    g157(.A(KEYINPUT20), .ZN(new_n359_));
  INV_X1    g158(.A(new_n343_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n339_), .A2(new_n360_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n361_), .A2(new_n334_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n359_), .B1(new_n310_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT93), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n277_), .A2(new_n279_), .ZN(new_n365_));
  AND4_X1   g164(.A1(new_n364_), .A2(new_n348_), .A3(new_n365_), .A4(new_n309_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n364_), .B1(new_n282_), .B2(new_n348_), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n358_), .B(new_n363_), .C1(new_n366_), .C2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n369_));
  INV_X1    g168(.A(G92gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  XOR2_X1   g170(.A(G8gat), .B(G36gat), .Z(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT95), .B(G64gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n358_), .B(KEYINPUT92), .Z(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT20), .B1(new_n310_), .B2(new_n362_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n282_), .A2(new_n348_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n376_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n368_), .A2(new_n375_), .A3(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n375_), .B1(new_n368_), .B2(new_n379_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n356_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT100), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  OAI211_X1 g183(.A(KEYINPUT100), .B(new_n356_), .C1(new_n380_), .C2(new_n381_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n368_), .A2(new_n375_), .A3(new_n379_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT99), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n310_), .A2(new_n362_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT20), .ZN(new_n389_));
  INV_X1    g188(.A(new_n367_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n282_), .A2(new_n364_), .A3(new_n348_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n389_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  OR2_X1    g191(.A1(new_n377_), .A2(new_n378_), .ZN(new_n393_));
  OAI22_X1  g192(.A1(new_n392_), .A2(new_n358_), .B1(new_n393_), .B2(new_n376_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT98), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n375_), .B(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n356_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n384_), .A2(new_n385_), .B1(new_n387_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n355_), .A2(new_n398_), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n319_), .A2(new_n398_), .A3(new_n266_), .ZN(new_n400_));
  AOI211_X1 g199(.A(new_n245_), .B(new_n214_), .C1(new_n248_), .C2(new_n249_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n253_), .A2(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n264_), .B1(new_n402_), .B2(new_n258_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n252_), .A2(new_n257_), .A3(new_n255_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n403_), .A2(KEYINPUT96), .A3(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(KEYINPUT96), .B1(new_n403_), .B2(new_n404_), .ZN(new_n406_));
  OR2_X1    g205(.A1(new_n380_), .A2(new_n381_), .ZN(new_n407_));
  NOR3_X1   g206(.A1(new_n405_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n264_), .B1(new_n263_), .B2(new_n260_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT33), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT33), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n411_), .B(new_n264_), .C1(new_n263_), .C2(new_n260_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n408_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n368_), .A2(new_n379_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n375_), .A2(KEYINPUT32), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n417_), .B1(new_n394_), .B2(new_n416_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n418_), .B1(new_n262_), .B2(new_n265_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT97), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT97), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n421_), .B(new_n418_), .C1(new_n262_), .C2(new_n265_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n414_), .A2(new_n420_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n319_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n400_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n354_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n399_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G15gat), .B(G22gat), .ZN(new_n428_));
  INV_X1    g227(.A(G1gat), .ZN(new_n429_));
  INV_X1    g228(.A(G8gat), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT14), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G1gat), .B(G8gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G43gat), .B(G50gat), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT76), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n435_), .A2(new_n436_), .ZN(new_n438_));
  XOR2_X1   g237(.A(G29gat), .B(G36gat), .Z(new_n439_));
  OR3_X1    g238(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n439_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n434_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n441_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT15), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n442_), .B1(new_n444_), .B2(new_n434_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G229gat), .A2(G233gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  XOR2_X1   g246(.A(new_n443_), .B(new_n434_), .Z(new_n448_));
  INV_X1    g247(.A(new_n446_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n447_), .A2(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(G169gat), .B(G197gat), .Z(new_n452_));
  XNOR2_X1  g251(.A(G113gat), .B(G141gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n454_), .A2(KEYINPUT80), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n451_), .B(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G230gat), .A2(G233gat), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n457_), .B(KEYINPUT64), .Z(new_n458_));
  XNOR2_X1  g257(.A(G71gat), .B(G78gat), .ZN(new_n459_));
  XOR2_X1   g258(.A(G57gat), .B(G64gat), .Z(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n459_), .B1(new_n461_), .B2(KEYINPUT11), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n462_), .B1(KEYINPUT11), .B2(new_n461_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n459_), .A3(KEYINPUT11), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT9), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT65), .B(G92gat), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n467_), .B1(new_n468_), .B2(new_n203_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT66), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  OAI211_X1 g270(.A(KEYINPUT66), .B(new_n467_), .C1(new_n468_), .C2(new_n203_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G85gat), .B(G92gat), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n473_), .B1(KEYINPUT9), .B2(new_n370_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n471_), .A2(new_n472_), .A3(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT10), .B(G99gat), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n476_), .A2(G106gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G99gat), .A2(G106gat), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT6), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n477_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n475_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT67), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT67), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n475_), .A2(new_n486_), .A3(new_n483_), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n482_), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NOR3_X1   g290(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  AOI211_X1 g292(.A(KEYINPUT8), .B(new_n473_), .C1(new_n489_), .C2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT8), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT68), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n482_), .A2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT69), .B1(new_n491_), .B2(new_n492_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n480_), .A2(KEYINPUT68), .A3(new_n481_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(G99gat), .A2(G106gat), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT7), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT69), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(new_n503_), .A3(new_n490_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n497_), .A2(new_n498_), .A3(new_n499_), .A4(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n473_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT70), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n495_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n505_), .A2(KEYINPUT70), .A3(new_n506_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n494_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n466_), .B1(new_n488_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n509_), .A2(new_n510_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n494_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n485_), .A2(new_n487_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n515_), .A2(new_n516_), .A3(new_n465_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n458_), .B1(new_n512_), .B2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT71), .ZN(new_n519_));
  XOR2_X1   g318(.A(KEYINPUT72), .B(KEYINPUT5), .Z(new_n520_));
  XNOR2_X1  g319(.A(G120gat), .B(G148gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(G176gat), .B(G204gat), .Z(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n512_), .A2(new_n517_), .A3(KEYINPUT12), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n515_), .A2(new_n516_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT12), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n526_), .A2(new_n527_), .A3(new_n466_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n525_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n458_), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n519_), .A2(new_n524_), .A3(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n524_), .B(KEYINPUT73), .Z(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n533_), .B1(new_n519_), .B2(new_n530_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT13), .ZN(new_n535_));
  OR3_X1    g334(.A1(new_n531_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n535_), .B1(new_n531_), .B2(new_n534_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n427_), .A2(new_n456_), .A3(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n515_), .A2(new_n516_), .A3(new_n443_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT77), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT77), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n515_), .A2(new_n543_), .A3(new_n516_), .A4(new_n443_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n526_), .A2(new_n444_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n542_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G232gat), .A2(G233gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(KEYINPUT75), .B(KEYINPUT35), .Z(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n546_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n546_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n549_), .B(new_n551_), .ZN(new_n556_));
  AOI22_X1  g355(.A1(new_n554_), .A2(KEYINPUT78), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT36), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G134gat), .B(G162gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n559_), .B(new_n560_), .Z(new_n561_));
  AOI22_X1  g360(.A1(new_n541_), .A2(KEYINPUT77), .B1(new_n526_), .B2(new_n444_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n552_), .B1(new_n562_), .B2(new_n544_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT78), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n557_), .A2(new_n558_), .A3(new_n561_), .A4(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n561_), .A2(new_n558_), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n561_), .A2(new_n558_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n562_), .A2(new_n544_), .A3(new_n556_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n569_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n554_), .A2(KEYINPUT78), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n567_), .B(new_n568_), .C1(new_n570_), .C2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n566_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT37), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT79), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n434_), .B(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(new_n465_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G127gat), .B(G155gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(new_n271_), .ZN(new_n581_));
  XOR2_X1   g380(.A(KEYINPUT16), .B(G183gat), .Z(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT17), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n579_), .A2(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n583_), .B(KEYINPUT17), .Z(new_n586_));
  AOI21_X1  g385(.A(new_n585_), .B1(new_n579_), .B2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n566_), .A2(new_n572_), .A3(KEYINPUT37), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n575_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n540_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n591_), .A2(new_n429_), .A3(new_n267_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT38), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n427_), .A2(new_n573_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT101), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n456_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n587_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n538_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n596_), .A2(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n600_), .A2(new_n267_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n593_), .B1(new_n601_), .B2(new_n429_), .ZN(G1324gat));
  INV_X1    g401(.A(new_n398_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n591_), .A2(new_n430_), .A3(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n594_), .A2(new_n595_), .ZN(new_n605_));
  AOI21_X1  g404(.A(KEYINPUT101), .B1(new_n427_), .B2(new_n573_), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n603_), .B(new_n599_), .C1(new_n605_), .C2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT102), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n430_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT39), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n596_), .A2(KEYINPUT102), .A3(new_n603_), .A4(new_n599_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n609_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n610_), .B1(new_n609_), .B2(new_n611_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n604_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT40), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  OAI211_X1 g415(.A(KEYINPUT40), .B(new_n604_), .C1(new_n612_), .C2(new_n613_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1325gat));
  INV_X1    g417(.A(G15gat), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n591_), .A2(new_n619_), .A3(new_n426_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n619_), .B1(new_n600_), .B2(new_n426_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n621_), .A2(new_n622_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n620_), .B1(new_n623_), .B2(new_n624_), .ZN(G1326gat));
  INV_X1    g424(.A(G22gat), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n591_), .A2(new_n626_), .A3(new_n319_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n600_), .A2(new_n319_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(G22gat), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n629_), .A2(KEYINPUT42), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(KEYINPUT42), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n627_), .B1(new_n630_), .B2(new_n631_), .ZN(G1327gat));
  NAND4_X1  g431(.A1(new_n536_), .A2(new_n537_), .A3(new_n456_), .A4(new_n598_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT104), .Z(new_n634_));
  INV_X1    g433(.A(KEYINPUT43), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n575_), .A2(new_n588_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n427_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n635_), .B1(new_n427_), .B2(new_n636_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n634_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT44), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n634_), .B(KEYINPUT44), .C1(new_n637_), .C2(new_n638_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n641_), .A2(new_n267_), .A3(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(G29gat), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n573_), .A2(new_n587_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n540_), .A2(new_n645_), .ZN(new_n646_));
  OR3_X1    g445(.A1(new_n646_), .A2(G29gat), .A3(new_n266_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n644_), .A2(new_n647_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT105), .Z(G1328gat));
  NAND3_X1  g448(.A1(new_n641_), .A2(new_n603_), .A3(new_n642_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(KEYINPUT106), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT106), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n641_), .A2(new_n652_), .A3(new_n603_), .A4(new_n642_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n651_), .A2(G36gat), .A3(new_n653_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n646_), .A2(G36gat), .A3(new_n398_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT45), .Z(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT46), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n654_), .A2(new_n656_), .A3(KEYINPUT46), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1329gat));
  NAND3_X1  g460(.A1(new_n641_), .A2(new_n426_), .A3(new_n642_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(G43gat), .ZN(new_n663_));
  OR3_X1    g462(.A1(new_n646_), .A2(G43gat), .A3(new_n354_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g465(.A(G50gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n641_), .A2(new_n319_), .A3(new_n642_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT107), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n667_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n670_), .B1(new_n669_), .B2(new_n668_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n319_), .A2(new_n667_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT108), .Z(new_n673_));
  OAI21_X1  g472(.A(new_n671_), .B1(new_n646_), .B2(new_n673_), .ZN(G1331gat));
  INV_X1    g473(.A(KEYINPUT110), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n539_), .A2(new_n456_), .A3(new_n598_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n596_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT109), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT109), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n596_), .A2(new_n679_), .A3(new_n676_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n678_), .A2(new_n267_), .A3(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(G57gat), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n539_), .A2(new_n456_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n683_), .A2(new_n427_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n684_), .A2(new_n590_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n266_), .A2(G57gat), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n675_), .B1(new_n682_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n687_), .ZN(new_n689_));
  AOI211_X1 g488(.A(KEYINPUT110), .B(new_n689_), .C1(new_n681_), .C2(G57gat), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n688_), .A2(new_n690_), .ZN(G1332gat));
  NAND3_X1  g490(.A1(new_n678_), .A2(new_n603_), .A3(new_n680_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(G64gat), .ZN(new_n693_));
  XNOR2_X1  g492(.A(KEYINPUT111), .B(KEYINPUT48), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n692_), .A2(G64gat), .A3(new_n694_), .ZN(new_n697_));
  INV_X1    g496(.A(G64gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n685_), .A2(new_n698_), .A3(new_n603_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n696_), .A2(new_n697_), .A3(new_n699_), .ZN(G1333gat));
  INV_X1    g499(.A(G71gat), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n685_), .A2(new_n701_), .A3(new_n426_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n678_), .A2(new_n426_), .A3(new_n680_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT49), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n703_), .A2(new_n704_), .A3(G71gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n703_), .B2(G71gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n702_), .B1(new_n705_), .B2(new_n706_), .ZN(G1334gat));
  INV_X1    g506(.A(G78gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n685_), .A2(new_n708_), .A3(new_n319_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n678_), .A2(new_n319_), .A3(new_n680_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT50), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n710_), .A2(new_n711_), .A3(G78gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n710_), .B2(G78gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n709_), .B1(new_n712_), .B2(new_n713_), .ZN(G1335gat));
  AND2_X1   g513(.A1(new_n684_), .A2(new_n645_), .ZN(new_n715_));
  AOI21_X1  g514(.A(G85gat), .B1(new_n715_), .B2(new_n267_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n427_), .A2(new_n636_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT43), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n427_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n720_), .A2(KEYINPUT112), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(KEYINPUT112), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n683_), .A2(new_n598_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n721_), .A2(new_n722_), .A3(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n266_), .A2(new_n203_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT113), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n716_), .B1(new_n726_), .B2(new_n728_), .ZN(G1336gat));
  AOI21_X1  g528(.A(G92gat), .B1(new_n715_), .B2(new_n603_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n398_), .A2(new_n468_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n726_), .B2(new_n731_), .ZN(G1337gat));
  OAI21_X1  g531(.A(G99gat), .B1(new_n725_), .B2(new_n354_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n354_), .A2(new_n476_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n715_), .A2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT114), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n733_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT51), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT51), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n733_), .A2(new_n739_), .A3(new_n736_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(G1338gat));
  AOI211_X1 g540(.A(new_n424_), .B(new_n723_), .C1(new_n718_), .C2(new_n719_), .ZN(new_n742_));
  INV_X1    g541(.A(G106gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(KEYINPUT115), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n720_), .A2(new_n319_), .A3(new_n724_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT115), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n745_), .A2(new_n746_), .A3(G106gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n744_), .A2(new_n747_), .A3(KEYINPUT52), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n715_), .A2(new_n743_), .A3(new_n319_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT52), .B1(new_n744_), .B2(new_n747_), .ZN(new_n751_));
  OAI21_X1  g550(.A(KEYINPUT53), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n751_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT53), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n753_), .A2(new_n754_), .A3(new_n749_), .A4(new_n748_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n752_), .A2(new_n755_), .ZN(G1339gat));
  NOR2_X1   g555(.A1(new_n319_), .A2(new_n354_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n603_), .A2(new_n266_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n458_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n525_), .A2(new_n759_), .A3(new_n528_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT55), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n759_), .B1(new_n525_), .B2(new_n528_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT55), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n529_), .A2(new_n764_), .A3(new_n458_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n532_), .ZN(new_n766_));
  OAI21_X1  g565(.A(KEYINPUT56), .B1(new_n763_), .B2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n530_), .A2(KEYINPUT55), .A3(new_n760_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT56), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n768_), .A2(new_n769_), .A3(new_n532_), .A4(new_n765_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n519_), .A2(new_n524_), .A3(new_n530_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n767_), .A2(new_n770_), .A3(new_n456_), .A4(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n447_), .A2(new_n454_), .A3(new_n450_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n445_), .A2(new_n449_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n454_), .B1(new_n448_), .B2(new_n446_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n775_), .B1(new_n778_), .B2(KEYINPUT118), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n779_), .B1(KEYINPUT118), .B2(new_n778_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n780_), .B1(new_n531_), .B2(new_n534_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n781_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n573_), .B1(new_n774_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT57), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n767_), .A2(new_n770_), .A3(new_n780_), .A4(new_n771_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT119), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n786_), .A2(KEYINPUT58), .ZN(new_n787_));
  AOI22_X1  g586(.A1(new_n786_), .A2(KEYINPUT58), .B1(new_n575_), .B2(new_n588_), .ZN(new_n788_));
  AOI22_X1  g587(.A1(new_n783_), .A2(new_n784_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  OAI211_X1 g588(.A(KEYINPUT57), .B(new_n573_), .C1(new_n774_), .C2(new_n782_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n587_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n536_), .A2(new_n537_), .A3(new_n597_), .ZN(new_n792_));
  XOR2_X1   g591(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  OR3_X1    g593(.A1(new_n589_), .A2(new_n792_), .A3(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n794_), .B1(new_n589_), .B2(new_n792_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n757_), .B(new_n758_), .C1(new_n791_), .C2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(G113gat), .B1(new_n799_), .B2(new_n456_), .ZN(new_n800_));
  OR2_X1    g599(.A1(new_n798_), .A2(KEYINPUT59), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n798_), .A2(KEYINPUT59), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n456_), .A2(G113gat), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n800_), .B1(new_n803_), .B2(new_n804_), .ZN(G1340gat));
  NAND3_X1  g604(.A1(new_n801_), .A2(new_n538_), .A3(new_n802_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(G120gat), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT60), .ZN(new_n808_));
  AOI21_X1  g607(.A(G120gat), .B1(new_n538_), .B2(new_n808_), .ZN(new_n809_));
  OR2_X1    g608(.A1(new_n809_), .A2(KEYINPUT120), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(KEYINPUT120), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n808_), .A2(G120gat), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n810_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n807_), .B1(new_n798_), .B2(new_n813_), .ZN(G1341gat));
  AOI21_X1  g613(.A(G127gat), .B1(new_n799_), .B2(new_n587_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n598_), .A2(KEYINPUT121), .ZN(new_n816_));
  MUX2_X1   g615(.A(KEYINPUT121), .B(new_n816_), .S(G127gat), .Z(new_n817_));
  AOI21_X1  g616(.A(new_n815_), .B1(new_n803_), .B2(new_n817_), .ZN(G1342gat));
  INV_X1    g617(.A(new_n573_), .ZN(new_n819_));
  AOI21_X1  g618(.A(G134gat), .B1(new_n799_), .B2(new_n819_), .ZN(new_n820_));
  XOR2_X1   g619(.A(KEYINPUT122), .B(G134gat), .Z(new_n821_));
  NAND2_X1  g620(.A1(new_n636_), .A2(new_n821_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(KEYINPUT123), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n820_), .B1(new_n803_), .B2(new_n823_), .ZN(G1343gat));
  NAND2_X1  g623(.A1(new_n783_), .A2(new_n784_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n787_), .A2(new_n788_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n790_), .A3(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n797_), .B1(new_n827_), .B2(new_n598_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n828_), .A2(new_n266_), .A3(new_n603_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n424_), .A2(new_n426_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n831_), .A2(new_n597_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(new_n222_), .ZN(G1344gat));
  NOR2_X1   g632(.A1(new_n831_), .A2(new_n539_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(new_n223_), .ZN(G1345gat));
  AND2_X1   g634(.A1(new_n829_), .A2(new_n830_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n587_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(KEYINPUT61), .B(G155gat), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n837_), .B(new_n838_), .ZN(G1346gat));
  AND3_X1   g638(.A1(new_n836_), .A2(G162gat), .A3(new_n636_), .ZN(new_n840_));
  AOI21_X1  g639(.A(G162gat), .B1(new_n836_), .B2(new_n819_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n840_), .A2(new_n841_), .ZN(G1347gat));
  INV_X1    g641(.A(KEYINPUT62), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n828_), .A2(new_n398_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n355_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n845_), .A2(new_n597_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n843_), .B1(new_n846_), .B2(new_n341_), .ZN(new_n847_));
  OAI211_X1 g646(.A(KEYINPUT62), .B(G169gat), .C1(new_n845_), .C2(new_n597_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n325_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n847_), .A2(new_n848_), .A3(new_n849_), .ZN(G1348gat));
  NOR2_X1   g649(.A1(new_n845_), .A2(new_n539_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(new_n326_), .ZN(G1349gat));
  NOR2_X1   g651(.A1(new_n845_), .A2(new_n598_), .ZN(new_n853_));
  MUX2_X1   g652(.A(G183gat), .B(new_n335_), .S(new_n853_), .Z(G1350gat));
  INV_X1    g653(.A(new_n636_), .ZN(new_n855_));
  OAI21_X1  g654(.A(G190gat), .B1(new_n845_), .B2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n819_), .A2(new_n336_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n845_), .B2(new_n857_), .ZN(G1351gat));
  NOR2_X1   g657(.A1(new_n424_), .A2(new_n267_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n354_), .ZN(new_n860_));
  NOR4_X1   g659(.A1(new_n828_), .A2(new_n398_), .A3(new_n597_), .A4(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT125), .B1(new_n861_), .B2(KEYINPUT124), .ZN(new_n862_));
  AOI21_X1  g661(.A(G197gat), .B1(new_n861_), .B2(KEYINPUT124), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT124), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT125), .ZN(new_n865_));
  INV_X1    g664(.A(new_n860_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n603_), .B(new_n866_), .C1(new_n791_), .C2(new_n797_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n864_), .B(new_n865_), .C1(new_n867_), .C2(new_n597_), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n862_), .A2(new_n863_), .A3(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n863_), .B1(new_n862_), .B2(new_n868_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1352gat));
  INV_X1    g670(.A(new_n867_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n538_), .ZN(new_n873_));
  AND2_X1   g672(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n874_));
  NOR2_X1   g673(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n873_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n873_), .B2(new_n874_), .ZN(G1353gat));
  NOR2_X1   g676(.A1(new_n867_), .A2(new_n598_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n878_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n879_));
  XOR2_X1   g678(.A(KEYINPUT63), .B(G211gat), .Z(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n878_), .B2(new_n880_), .ZN(G1354gat));
  XNOR2_X1  g680(.A(KEYINPUT127), .B(G218gat), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n867_), .A2(new_n855_), .A3(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n872_), .A2(new_n819_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n883_), .B1(new_n884_), .B2(new_n882_), .ZN(G1355gat));
endmodule


