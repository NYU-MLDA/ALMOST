//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 0 0 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT66), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT7), .ZN(new_n204_));
  AOI211_X1 g003(.A(G99gat), .B(G106gat), .C1(new_n203_), .C2(new_n204_), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n205_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT6), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT65), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n206_), .A2(new_n208_), .A3(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G85gat), .A2(G92gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n211_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT8), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT8), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n211_), .A2(new_n218_), .A3(new_n215_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n214_), .B1(new_n213_), .B2(KEYINPUT9), .ZN(new_n220_));
  NOR3_X1   g019(.A1(new_n213_), .A2(KEYINPUT64), .A3(KEYINPUT9), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT9), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n222_), .B1(new_n212_), .B2(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n220_), .B1(new_n221_), .B2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT10), .B(G99gat), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n226_), .A2(G106gat), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n227_), .A2(new_n208_), .ZN(new_n228_));
  AOI22_X1  g027(.A1(new_n217_), .A2(new_n219_), .B1(new_n225_), .B2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G57gat), .B(G64gat), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n230_), .A2(KEYINPUT11), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(KEYINPUT11), .ZN(new_n232_));
  XOR2_X1   g031(.A(G71gat), .B(G78gat), .Z(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n232_), .A2(new_n233_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n229_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n228_), .A2(new_n225_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n219_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n218_), .B1(new_n211_), .B2(new_n215_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n238_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n236_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n237_), .A2(new_n243_), .A3(KEYINPUT12), .ZN(new_n244_));
  OR3_X1    g043(.A1(new_n229_), .A2(KEYINPUT12), .A3(new_n236_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G230gat), .A2(G233gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n237_), .A2(new_n243_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(G230gat), .A3(G233gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(G120gat), .B(G148gat), .Z(new_n252_));
  XNOR2_X1  g051(.A(G176gat), .B(G204gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n251_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n248_), .A2(new_n250_), .A3(new_n256_), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n258_), .A2(KEYINPUT13), .A3(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT13), .B1(new_n258_), .B2(new_n259_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  XOR2_X1   g062(.A(G15gat), .B(G22gat), .Z(new_n264_));
  NAND2_X1  g063(.A1(G1gat), .A2(G8gat), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n265_), .A2(KEYINPUT14), .ZN(new_n266_));
  OR3_X1    g065(.A1(new_n264_), .A2(KEYINPUT75), .A3(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT75), .B1(new_n264_), .B2(new_n266_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n265_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(G1gat), .A2(G8gat), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n269_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n270_), .A2(new_n271_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n267_), .A2(new_n273_), .A3(new_n268_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(G29gat), .B(G36gat), .Z(new_n276_));
  XOR2_X1   g075(.A(G43gat), .B(G50gat), .Z(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT15), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n275_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n272_), .A2(new_n278_), .A3(new_n274_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G229gat), .A2(G233gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT80), .B1(new_n282_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT80), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n280_), .A2(new_n286_), .A3(new_n283_), .A4(new_n281_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT79), .ZN(new_n289_));
  INV_X1    g088(.A(new_n281_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n278_), .B1(new_n272_), .B2(new_n274_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n289_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n291_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(KEYINPUT79), .A3(new_n281_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n283_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n288_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G113gat), .B(G141gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G169gat), .B(G197gat), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n297_), .B(new_n298_), .Z(new_n299_));
  NAND2_X1  g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n299_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n301_), .B1(new_n288_), .B2(new_n295_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n263_), .A2(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(G127gat), .B(G155gat), .Z(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G183gat), .B(G211gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G231gat), .A2(G233gat), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n236_), .B(new_n311_), .Z(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(new_n275_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n310_), .B1(new_n313_), .B2(KEYINPUT17), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n314_), .B1(KEYINPUT17), .B2(new_n310_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT77), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n315_), .B(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n305_), .A2(new_n318_), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n319_), .B(KEYINPUT103), .Z(new_n320_));
  NAND2_X1  g119(.A1(G225gat), .A2(G233gat), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT2), .ZN(new_n323_));
  AND3_X1   g122(.A1(KEYINPUT85), .A2(G141gat), .A3(G148gat), .ZN(new_n324_));
  AOI21_X1  g123(.A(KEYINPUT85), .B1(G141gat), .B2(G148gat), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n323_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT87), .ZN(new_n327_));
  NAND3_X1  g126(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT88), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(KEYINPUT88), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n331_));
  INV_X1    g130(.A(G141gat), .ZN(new_n332_));
  INV_X1    g131(.A(G148gat), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(new_n333_), .A3(KEYINPUT3), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT3), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n335_), .B1(G141gat), .B2(G148gat), .ZN(new_n336_));
  AOI22_X1  g135(.A1(new_n330_), .A2(new_n331_), .B1(new_n334_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT87), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n338_), .B(new_n323_), .C1(new_n324_), .C2(new_n325_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n327_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G155gat), .A2(G162gat), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(G155gat), .A2(G162gat), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n340_), .A2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n341_), .B1(new_n343_), .B2(KEYINPUT1), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT86), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  OAI211_X1 g147(.A(KEYINPUT86), .B(new_n341_), .C1(new_n343_), .C2(KEYINPUT1), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n341_), .A2(KEYINPUT1), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n348_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n324_), .A2(new_n325_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n352_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n345_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT89), .ZN(new_n356_));
  AOI22_X1  g155(.A1(new_n340_), .A2(new_n344_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT89), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  XOR2_X1   g158(.A(G127gat), .B(G134gat), .Z(new_n360_));
  XOR2_X1   g159(.A(G113gat), .B(G120gat), .Z(new_n361_));
  XOR2_X1   g160(.A(new_n360_), .B(new_n361_), .Z(new_n362_));
  NAND3_X1  g161(.A1(new_n356_), .A2(new_n359_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n362_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n357_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n363_), .A2(KEYINPUT4), .A3(new_n365_), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n345_), .A2(new_n358_), .A3(new_n354_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n358_), .B1(new_n345_), .B2(new_n354_), .ZN(new_n368_));
  NOR3_X1   g167(.A1(new_n367_), .A2(new_n368_), .A3(new_n364_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT4), .ZN(new_n370_));
  AOI21_X1  g169(.A(KEYINPUT98), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n356_), .A2(new_n370_), .A3(new_n359_), .A4(new_n362_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT98), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n322_), .B(new_n366_), .C1(new_n371_), .C2(new_n374_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n363_), .A2(new_n365_), .A3(new_n321_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G1gat), .B(G29gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(G85gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(KEYINPUT0), .B(G57gat), .ZN(new_n381_));
  XOR2_X1   g180(.A(new_n380_), .B(new_n381_), .Z(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n378_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT101), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n372_), .B(KEYINPUT98), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n366_), .A2(new_n322_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n377_), .B(new_n382_), .C1(new_n386_), .C2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n384_), .A2(new_n385_), .A3(new_n388_), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n366_), .A2(new_n322_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n369_), .A2(KEYINPUT98), .A3(new_n370_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n372_), .A2(new_n373_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  AOI211_X1 g192(.A(new_n376_), .B(new_n383_), .C1(new_n390_), .C2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n382_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT101), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n389_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n356_), .A2(KEYINPUT29), .A3(new_n359_), .ZN(new_n398_));
  AND2_X1   g197(.A1(G228gat), .A2(G233gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G211gat), .B(G218gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT92), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT21), .ZN(new_n402_));
  INV_X1    g201(.A(G197gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(G204gat), .ZN(new_n404_));
  INV_X1    g203(.A(G204gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(G197gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT93), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n402_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n401_), .B(new_n409_), .C1(new_n408_), .C2(new_n407_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n404_), .A2(new_n406_), .A3(KEYINPUT91), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n411_), .B(KEYINPUT21), .C1(KEYINPUT91), .C2(new_n404_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n404_), .A2(new_n406_), .A3(new_n402_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n412_), .A2(new_n413_), .A3(new_n400_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n399_), .B1(new_n410_), .B2(new_n414_), .ZN(new_n415_));
  XOR2_X1   g214(.A(new_n400_), .B(KEYINPUT92), .Z(new_n416_));
  OAI21_X1  g215(.A(new_n409_), .B1(new_n408_), .B2(new_n407_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n414_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT29), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n418_), .B1(new_n357_), .B2(new_n419_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n398_), .A2(new_n415_), .B1(new_n399_), .B2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G78gat), .B(G106gat), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT94), .B1(new_n421_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n356_), .A2(new_n359_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n419_), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(KEYINPUT29), .B1(new_n356_), .B2(new_n359_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n429_), .A2(new_n426_), .ZN(new_n430_));
  XOR2_X1   g229(.A(G22gat), .B(G50gat), .Z(new_n431_));
  NOR3_X1   g230(.A1(new_n428_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n431_), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n429_), .A2(new_n426_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n433_), .B1(new_n434_), .B2(new_n427_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n424_), .B1(new_n432_), .B2(new_n435_), .ZN(new_n436_));
  OR2_X1    g235(.A1(new_n421_), .A2(new_n423_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n421_), .A2(new_n423_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n436_), .A2(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n431_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n434_), .A2(new_n433_), .A3(new_n427_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n443_), .A2(new_n438_), .A3(new_n437_), .A4(new_n424_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n440_), .A2(new_n444_), .ZN(new_n445_));
  XOR2_X1   g244(.A(G8gat), .B(G36gat), .Z(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT18), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G64gat), .B(G92gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT22), .B(G169gat), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT97), .ZN(new_n452_));
  OR2_X1    g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(KEYINPUT83), .B(G176gat), .Z(new_n454_));
  NAND2_X1  g253(.A1(new_n451_), .A2(new_n452_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n453_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G183gat), .A2(G190gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT23), .ZN(new_n458_));
  OR2_X1    g257(.A1(G183gat), .A2(G190gat), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n458_), .A2(new_n459_), .B1(G169gat), .B2(G176gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n456_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n462_));
  NOR3_X1   g261(.A1(KEYINPUT82), .A2(G169gat), .A3(G176gat), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT82), .B1(G169gat), .B2(G176gat), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n462_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G169gat), .A2(G176gat), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n464_), .A2(new_n462_), .A3(new_n465_), .A4(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT26), .B(G190gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT25), .B(G183gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n468_), .A2(new_n458_), .A3(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n461_), .B1(new_n466_), .B2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT20), .B1(new_n473_), .B2(new_n418_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n454_), .A2(new_n451_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n460_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(G183gat), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT25), .B1(new_n477_), .B2(KEYINPUT81), .ZN(new_n478_));
  OR2_X1    g277(.A1(new_n477_), .A2(KEYINPUT25), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n469_), .B(new_n478_), .C1(new_n479_), .C2(KEYINPUT81), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n464_), .A2(KEYINPUT24), .A3(new_n465_), .A4(new_n467_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT24), .ZN(new_n482_));
  INV_X1    g281(.A(new_n465_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n482_), .B1(new_n483_), .B2(new_n463_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n480_), .A2(new_n481_), .A3(new_n458_), .A4(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n476_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n418_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G226gat), .A2(G233gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  NOR3_X1   g290(.A1(new_n474_), .A2(new_n488_), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n491_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT20), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n494_), .B1(new_n473_), .B2(new_n418_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n410_), .A2(new_n414_), .A3(new_n485_), .A4(new_n476_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n493_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n450_), .B1(new_n492_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n473_), .A2(new_n418_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n499_), .A2(new_n496_), .A3(KEYINPUT20), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n491_), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n473_), .A2(new_n418_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n502_), .A2(new_n487_), .A3(KEYINPUT20), .A4(new_n493_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n501_), .A2(new_n503_), .A3(new_n449_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n498_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT27), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n491_), .B1(new_n474_), .B2(new_n488_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n508_), .B1(new_n491_), .B2(new_n500_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n450_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n510_), .A2(KEYINPUT27), .A3(new_n504_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n507_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT30), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n486_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n486_), .A2(new_n513_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT84), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G71gat), .B(G99gat), .ZN(new_n519_));
  INV_X1    g318(.A(G43gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G227gat), .A2(G233gat), .ZN(new_n522_));
  INV_X1    g321(.A(G15gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n521_), .B(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n518_), .A2(new_n525_), .ZN(new_n526_));
  NOR3_X1   g325(.A1(new_n515_), .A2(KEYINPUT84), .A3(new_n516_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n525_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n362_), .B(KEYINPUT31), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  OR3_X1    g330(.A1(new_n526_), .A2(new_n529_), .A3(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n531_), .B1(new_n526_), .B2(new_n529_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n512_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n397_), .A2(new_n445_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n449_), .A2(KEYINPUT32), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n537_), .B1(new_n492_), .B2(new_n497_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n538_), .B1(new_n509_), .B2(new_n537_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n539_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT100), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT99), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT33), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n543_), .B1(new_n388_), .B2(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n376_), .B1(new_n390_), .B2(new_n393_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n546_), .A2(KEYINPUT99), .A3(KEYINPUT33), .A4(new_n382_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n388_), .A2(new_n544_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n393_), .A2(new_n321_), .A3(new_n366_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n363_), .A2(new_n365_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n382_), .B1(new_n550_), .B2(new_n322_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n505_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n545_), .A2(new_n547_), .A3(new_n548_), .A4(new_n552_), .ZN(new_n553_));
  OAI211_X1 g352(.A(KEYINPUT100), .B(new_n539_), .C1(new_n394_), .C2(new_n395_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n542_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(new_n445_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n512_), .B1(new_n440_), .B2(new_n444_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n397_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n532_), .A2(new_n533_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n536_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n278_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n563_), .B(new_n238_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n564_), .B1(new_n229_), .B2(new_n279_), .ZN(new_n565_));
  XOR2_X1   g364(.A(KEYINPUT68), .B(KEYINPUT34), .Z(new_n566_));
  NAND2_X1  g365(.A1(G232gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT35), .ZN(new_n569_));
  AOI21_X1  g368(.A(KEYINPUT70), .B1(new_n565_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n565_), .A2(KEYINPUT70), .A3(new_n569_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT35), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n568_), .A2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(KEYINPUT69), .B1(new_n565_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n279_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n241_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT69), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n568_), .A2(new_n573_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n577_), .A2(new_n578_), .A3(new_n564_), .A4(new_n579_), .ZN(new_n580_));
  AOI22_X1  g379(.A1(new_n571_), .A2(new_n572_), .B1(new_n575_), .B2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G190gat), .B(G218gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G134gat), .B(G162gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n584_), .B(KEYINPUT36), .Z(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(KEYINPUT72), .B1(new_n581_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT72), .ZN(new_n588_));
  INV_X1    g387(.A(new_n572_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n589_), .A2(new_n570_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n575_), .A2(new_n580_), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n588_), .B(new_n585_), .C1(new_n590_), .C2(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n584_), .A2(KEYINPUT36), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n581_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n587_), .A2(new_n592_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n562_), .A2(new_n596_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n320_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT104), .ZN(new_n599_));
  INV_X1    g398(.A(new_n397_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n202_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  AOI22_X1  g400(.A1(new_n555_), .A2(new_n445_), .B1(new_n397_), .B2(new_n557_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n535_), .B1(new_n602_), .B2(new_n560_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(new_n303_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT102), .ZN(new_n605_));
  XOR2_X1   g404(.A(KEYINPUT73), .B(KEYINPUT37), .Z(new_n606_));
  NAND4_X1  g405(.A1(new_n587_), .A2(new_n592_), .A3(new_n594_), .A4(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT74), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n571_), .A2(new_n572_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n575_), .A2(new_n580_), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n609_), .A2(new_n610_), .A3(new_n593_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n585_), .B(KEYINPUT71), .Z(new_n612_));
  AOI21_X1  g411(.A(new_n612_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n613_));
  OAI21_X1  g412(.A(KEYINPUT37), .B1(new_n611_), .B2(new_n613_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n607_), .A2(new_n608_), .A3(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n608_), .B1(new_n607_), .B2(new_n614_), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n262_), .B(new_n318_), .C1(new_n615_), .C2(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT78), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n605_), .A2(new_n618_), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n619_), .A2(G1gat), .A3(new_n397_), .ZN(new_n620_));
  OAI21_X1  g419(.A(KEYINPUT38), .B1(new_n601_), .B2(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n621_), .B1(KEYINPUT38), .B2(new_n620_), .ZN(G1324gat));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n598_), .A2(new_n512_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n623_), .B1(new_n624_), .B2(G8gat), .ZN(new_n625_));
  INV_X1    g424(.A(G8gat), .ZN(new_n626_));
  AOI211_X1 g425(.A(KEYINPUT39), .B(new_n626_), .C1(new_n598_), .C2(new_n512_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n619_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n629_), .A2(new_n626_), .A3(new_n512_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(G1325gat));
  NAND3_X1  g432(.A1(new_n629_), .A2(new_n523_), .A3(new_n560_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n523_), .B1(new_n599_), .B2(new_n560_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n635_), .A2(KEYINPUT41), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(KEYINPUT41), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n634_), .B1(new_n636_), .B2(new_n637_), .ZN(G1326gat));
  INV_X1    g437(.A(G22gat), .ZN(new_n639_));
  INV_X1    g438(.A(new_n445_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n629_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n639_), .B1(new_n599_), .B2(new_n640_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT42), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n642_), .A2(new_n643_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n641_), .B1(new_n644_), .B2(new_n645_), .ZN(G1327gat));
  NOR2_X1   g445(.A1(new_n318_), .A2(new_n595_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n647_), .A2(new_n262_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n605_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(G29gat), .B1(new_n650_), .B2(new_n600_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT44), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT43), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n615_), .A2(new_n616_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n603_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n653_), .B1(new_n603_), .B2(new_n654_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n318_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n305_), .A2(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n652_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n654_), .ZN(new_n661_));
  OAI21_X1  g460(.A(KEYINPUT43), .B1(new_n562_), .B2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n603_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n664_), .A2(KEYINPUT44), .A3(new_n305_), .A4(new_n658_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n660_), .A2(new_n665_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n600_), .A2(G29gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n651_), .B1(new_n666_), .B2(new_n667_), .ZN(G1328gat));
  INV_X1    g467(.A(KEYINPUT107), .ZN(new_n669_));
  AOI21_X1  g468(.A(G36gat), .B1(new_n507_), .B2(new_n511_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n605_), .A2(new_n648_), .A3(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT45), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT45), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n605_), .A2(new_n673_), .A3(new_n648_), .A4(new_n670_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n660_), .A2(new_n665_), .A3(new_n512_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(G36gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n669_), .B1(new_n675_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n675_), .A2(new_n677_), .A3(new_n669_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n679_), .A2(new_n680_), .A3(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n680_), .B1(new_n679_), .B2(new_n681_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1329gat));
  NAND3_X1  g483(.A1(new_n666_), .A2(G43gat), .A3(new_n560_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n520_), .B1(new_n649_), .B2(new_n561_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g487(.A(G50gat), .B1(new_n650_), .B2(new_n640_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n640_), .A2(G50gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n666_), .B2(new_n690_), .ZN(G1331gat));
  AND4_X1   g490(.A1(new_n597_), .A2(new_n304_), .A3(new_n263_), .A4(new_n318_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n692_), .A2(G57gat), .A3(new_n600_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n693_), .A2(KEYINPUT108), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n693_), .A2(KEYINPUT108), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n263_), .A2(new_n304_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n562_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n607_), .A2(new_n614_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT74), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n607_), .A2(new_n608_), .A3(new_n614_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n658_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n697_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(G57gat), .B1(new_n703_), .B2(new_n600_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n694_), .A2(new_n695_), .A3(new_n704_), .ZN(G1332gat));
  INV_X1    g504(.A(G64gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n692_), .B2(new_n512_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n707_), .B(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n703_), .A2(new_n706_), .A3(new_n512_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT110), .Z(G1333gat));
  NAND2_X1  g511(.A1(new_n692_), .A2(new_n560_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(G71gat), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT49), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n561_), .A2(G71gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n715_), .B1(new_n702_), .B2(new_n716_), .ZN(G1334gat));
  INV_X1    g516(.A(G78gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n692_), .B2(new_n640_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n719_), .B(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n703_), .A2(new_n718_), .A3(new_n640_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1335gat));
  NAND2_X1  g522(.A1(new_n697_), .A2(new_n647_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT112), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n697_), .A2(KEYINPUT112), .A3(new_n647_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(G85gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n728_), .A2(new_n729_), .A3(new_n600_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n263_), .A2(new_n304_), .A3(new_n658_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(G85gat), .B1(new_n733_), .B2(new_n397_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n730_), .A2(new_n734_), .ZN(G1336gat));
  AOI21_X1  g534(.A(G92gat), .B1(new_n728_), .B2(new_n512_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n512_), .A2(G92gat), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT113), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n736_), .B1(new_n732_), .B2(new_n738_), .ZN(G1337gat));
  NAND2_X1  g538(.A1(new_n732_), .A2(new_n560_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(G99gat), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT114), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n561_), .A2(new_n226_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT115), .ZN(new_n744_));
  AOI22_X1  g543(.A1(new_n728_), .A2(new_n743_), .B1(new_n744_), .B2(KEYINPUT51), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n742_), .A2(new_n745_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n744_), .A2(KEYINPUT51), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n746_), .B(new_n747_), .Z(G1338gat));
  XNOR2_X1  g547(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n749_));
  INV_X1    g548(.A(new_n731_), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n640_), .B(new_n750_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n751_));
  OAI21_X1  g550(.A(G106gat), .B1(new_n751_), .B2(KEYINPUT116), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT116), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n732_), .B2(new_n640_), .ZN(new_n754_));
  OAI21_X1  g553(.A(KEYINPUT52), .B1(new_n752_), .B2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n732_), .A2(new_n753_), .A3(new_n640_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n751_), .A2(KEYINPUT116), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT52), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n756_), .A2(new_n757_), .A3(new_n758_), .A4(G106gat), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n755_), .A2(new_n759_), .ZN(new_n760_));
  AOI211_X1 g559(.A(G106gat), .B(new_n445_), .C1(new_n726_), .C2(new_n727_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT118), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT118), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n760_), .A2(new_n765_), .A3(new_n762_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n749_), .B1(new_n764_), .B2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n765_), .B1(new_n760_), .B2(new_n762_), .ZN(new_n768_));
  AOI211_X1 g567(.A(KEYINPUT118), .B(new_n761_), .C1(new_n755_), .C2(new_n759_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n749_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n768_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n767_), .A2(new_n771_), .ZN(G1339gat));
  INV_X1    g571(.A(KEYINPUT125), .ZN(new_n773_));
  INV_X1    g572(.A(G113gat), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n534_), .A2(new_n600_), .A3(new_n445_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(KEYINPUT119), .B(KEYINPUT54), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n778_), .B1(new_n617_), .B2(new_n303_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT121), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT121), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n781_), .B(new_n778_), .C1(new_n617_), .C2(new_n303_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n701_), .A2(new_n304_), .A3(new_n262_), .A4(new_n777_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT120), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n617_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n787_), .A2(KEYINPUT120), .A3(new_n304_), .A4(new_n777_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n783_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n246_), .A2(KEYINPUT55), .ZN(new_n791_));
  NAND3_X1  g590(.A1(KEYINPUT122), .A2(G230gat), .A3(G233gat), .ZN(new_n792_));
  AOI22_X1  g591(.A1(new_n244_), .A2(new_n245_), .B1(G230gat), .B2(G233gat), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n791_), .B(new_n792_), .C1(new_n793_), .C2(KEYINPUT55), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n792_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n256_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT56), .B1(new_n794_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n794_), .A2(KEYINPUT56), .A3(new_n798_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n284_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n301_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n805_), .B1(new_n296_), .B2(new_n299_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n806_), .A2(new_n259_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n802_), .A2(KEYINPUT58), .A3(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT58), .B1(new_n802_), .B2(new_n807_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n801_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n303_), .B(new_n259_), .C1(new_n811_), .C2(new_n799_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n258_), .A2(new_n259_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n813_), .A2(new_n806_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n596_), .B1(new_n812_), .B2(new_n815_), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n810_), .A2(new_n654_), .B1(KEYINPUT57), .B2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(KEYINPUT57), .B2(new_n816_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n658_), .ZN(new_n819_));
  AOI211_X1 g618(.A(KEYINPUT59), .B(new_n776_), .C1(new_n790_), .C2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT124), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT123), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n822_), .B1(new_n816_), .B2(KEYINPUT57), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n303_), .A2(new_n259_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n824_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n595_), .B1(new_n825_), .B2(new_n814_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(KEYINPUT123), .A3(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n817_), .A2(new_n823_), .A3(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n658_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n776_), .B1(new_n790_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT59), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n821_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n783_), .A2(new_n789_), .B1(new_n829_), .B2(new_n658_), .ZN(new_n834_));
  OAI211_X1 g633(.A(KEYINPUT124), .B(KEYINPUT59), .C1(new_n834_), .C2(new_n776_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n820_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n774_), .B1(new_n836_), .B2(new_n303_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n831_), .A2(new_n774_), .A3(new_n303_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n773_), .B1(new_n837_), .B2(new_n839_), .ZN(new_n840_));
  AOI211_X1 g639(.A(new_n304_), .B(new_n820_), .C1(new_n833_), .C2(new_n835_), .ZN(new_n841_));
  OAI211_X1 g640(.A(KEYINPUT125), .B(new_n838_), .C1(new_n841_), .C2(new_n774_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(G1340gat));
  INV_X1    g642(.A(G120gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n262_), .B2(KEYINPUT60), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n831_), .B(new_n845_), .C1(KEYINPUT60), .C2(new_n844_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n836_), .A2(new_n263_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n847_), .B2(new_n844_), .ZN(G1341gat));
  INV_X1    g647(.A(G127gat), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n831_), .A2(new_n849_), .A3(new_n318_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n836_), .A2(new_n318_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n849_), .ZN(G1342gat));
  INV_X1    g651(.A(G134gat), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n831_), .A2(new_n853_), .A3(new_n596_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n836_), .A2(new_n654_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n853_), .ZN(G1343gat));
  NOR2_X1   g655(.A1(new_n834_), .A2(new_n560_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n397_), .A2(new_n445_), .A3(new_n512_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n304_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(new_n332_), .ZN(G1344gat));
  NAND3_X1  g660(.A1(new_n857_), .A2(new_n263_), .A3(new_n858_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g662(.A1(new_n859_), .A2(new_n658_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT61), .B(G155gat), .ZN(new_n865_));
  XOR2_X1   g664(.A(new_n864_), .B(new_n865_), .Z(G1346gat));
  OAI21_X1  g665(.A(G162gat), .B1(new_n859_), .B2(new_n661_), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n595_), .A2(G162gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n859_), .B2(new_n868_), .ZN(G1347gat));
  INV_X1    g668(.A(KEYINPUT62), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n640_), .B1(new_n790_), .B2(new_n819_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n397_), .A2(new_n512_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n872_), .A2(new_n561_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n874_), .A2(new_n304_), .ZN(new_n875_));
  INV_X1    g674(.A(G169gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n870_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n875_), .A2(new_n453_), .A3(new_n455_), .ZN(new_n878_));
  OAI211_X1 g677(.A(KEYINPUT62), .B(G169gat), .C1(new_n874_), .C2(new_n304_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n877_), .A2(new_n878_), .A3(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT126), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n877_), .A2(new_n878_), .A3(KEYINPUT126), .A4(new_n879_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1348gat));
  INV_X1    g683(.A(new_n874_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n263_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n834_), .A2(new_n640_), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n873_), .A2(G176gat), .A3(new_n263_), .ZN(new_n888_));
  AOI22_X1  g687(.A1(new_n886_), .A2(new_n454_), .B1(new_n887_), .B2(new_n888_), .ZN(G1349gat));
  NAND3_X1  g688(.A1(new_n887_), .A2(new_n318_), .A3(new_n873_), .ZN(new_n890_));
  NOR4_X1   g689(.A1(new_n872_), .A2(new_n658_), .A3(new_n470_), .A4(new_n561_), .ZN(new_n891_));
  AOI22_X1  g690(.A1(new_n890_), .A2(new_n477_), .B1(new_n871_), .B2(new_n891_), .ZN(G1350gat));
  OAI21_X1  g691(.A(G190gat), .B1(new_n874_), .B2(new_n661_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n596_), .A2(new_n469_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n874_), .B2(new_n894_), .ZN(G1351gat));
  NAND4_X1  g694(.A1(new_n857_), .A2(new_n397_), .A3(new_n640_), .A4(new_n512_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n304_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(new_n403_), .ZN(G1352gat));
  NOR2_X1   g697(.A1(new_n896_), .A2(new_n262_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n405_), .ZN(G1353gat));
  INV_X1    g699(.A(KEYINPUT63), .ZN(new_n901_));
  INV_X1    g700(.A(G211gat), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n318_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(KEYINPUT127), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n896_), .A2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n905_), .B(new_n906_), .ZN(G1354gat));
  OAI21_X1  g706(.A(G218gat), .B1(new_n896_), .B2(new_n661_), .ZN(new_n908_));
  OR2_X1    g707(.A1(new_n595_), .A2(G218gat), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n896_), .B2(new_n909_), .ZN(G1355gat));
endmodule


