//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n642_,
    new_n643_, new_n644_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n854_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n904_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(KEYINPUT84), .ZN(new_n205_));
  INV_X1    g004(.A(G204gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n206_), .A2(KEYINPUT84), .A3(G197gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT21), .ZN(new_n208_));
  OAI221_X1 g007(.A(new_n202_), .B1(KEYINPUT21), .B2(new_n204_), .C1(new_n205_), .C2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT21), .ZN(new_n210_));
  AOI211_X1 g009(.A(new_n210_), .B(new_n202_), .C1(KEYINPUT85), .C2(new_n203_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n211_), .B1(KEYINPUT85), .B2(new_n203_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT82), .B1(G155gat), .B2(G162gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NOR3_X1   g014(.A1(KEYINPUT82), .A2(G155gat), .A3(G162gat), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(new_n222_), .B(KEYINPUT83), .Z(new_n223_));
  NOR2_X1   g022(.A1(G141gat), .A2(G148gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n225_));
  OAI22_X1  g024(.A1(new_n224_), .A2(new_n225_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n226_), .B1(new_n225_), .B2(new_n224_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n219_), .B1(new_n223_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n224_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(new_n220_), .ZN(new_n230_));
  XOR2_X1   g029(.A(new_n218_), .B(KEYINPUT1), .Z(new_n231_));
  AOI21_X1  g030(.A(new_n230_), .B1(new_n231_), .B2(new_n217_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n228_), .A2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(KEYINPUT86), .B(KEYINPUT29), .Z(new_n234_));
  OAI21_X1  g033(.A(new_n213_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(G228gat), .A3(G233gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G228gat), .A2(G233gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT29), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n237_), .B(new_n213_), .C1(new_n233_), .C2(new_n238_), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n236_), .A2(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(G78gat), .B(G106gat), .Z(new_n241_));
  NOR2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT88), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n233_), .A2(new_n238_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT28), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G22gat), .B(G50gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n240_), .A2(new_n241_), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n243_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n242_), .A2(KEYINPUT88), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n240_), .A2(new_n241_), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT87), .B1(new_n240_), .B2(new_n241_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n247_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT87), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n242_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n248_), .ZN(new_n256_));
  AOI22_X1  g055(.A1(new_n249_), .A2(new_n250_), .B1(new_n253_), .B2(new_n256_), .ZN(new_n257_));
  XOR2_X1   g056(.A(G127gat), .B(G134gat), .Z(new_n258_));
  XNOR2_X1  g057(.A(G113gat), .B(G120gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n233_), .B(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G225gat), .A2(G233gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT99), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n261_), .A2(KEYINPUT4), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n262_), .B(KEYINPUT97), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n268_), .B(new_n260_), .C1(new_n228_), .C2(new_n232_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n266_), .A2(new_n267_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT98), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT98), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n266_), .A2(new_n272_), .A3(new_n267_), .A4(new_n269_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n265_), .A2(new_n271_), .A3(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G1gat), .B(G29gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(G85gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT0), .B(G57gat), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n276_), .B(new_n277_), .Z(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n274_), .A2(new_n279_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n265_), .A2(new_n278_), .A3(new_n271_), .A4(new_n273_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n257_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT103), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT27), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G226gat), .A2(G233gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(new_n288_), .B(KEYINPUT90), .Z(new_n289_));
  NOR2_X1   g088(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(G169gat), .ZN(new_n291_));
  INV_X1    g090(.A(G183gat), .ZN(new_n292_));
  INV_X1    g091(.A(G190gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT23), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT80), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  OR3_X1    g095(.A1(new_n292_), .A2(new_n293_), .A3(KEYINPUT23), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(G183gat), .A2(G190gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n291_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT95), .ZN(new_n301_));
  XOR2_X1   g100(.A(KEYINPUT26), .B(G190gat), .Z(new_n302_));
  XOR2_X1   g101(.A(new_n302_), .B(KEYINPUT93), .Z(new_n303_));
  XOR2_X1   g102(.A(KEYINPUT25), .B(G183gat), .Z(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT92), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307_));
  INV_X1    g106(.A(G169gat), .ZN(new_n308_));
  INV_X1    g107(.A(G176gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT24), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT94), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n307_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n312_), .B1(new_n311_), .B2(new_n310_), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n297_), .A2(new_n294_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT24), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n307_), .A2(new_n316_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n306_), .A2(new_n313_), .A3(new_n315_), .A4(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n301_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n213_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n291_), .B1(new_n314_), .B2(new_n299_), .ZN(new_n321_));
  OAI221_X1 g120(.A(new_n317_), .B1(new_n310_), .B2(new_n307_), .C1(new_n304_), .C2(new_n302_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n321_), .B1(new_n298_), .B2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT20), .B1(new_n213_), .B2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT91), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n289_), .B1(new_n320_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n213_), .A2(new_n323_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n288_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n327_), .A2(KEYINPUT20), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n319_), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n209_), .A2(new_n212_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n329_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n326_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G8gat), .B(G36gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT18), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G64gat), .B(G92gat), .ZN(new_n336_));
  XOR2_X1   g135(.A(new_n335_), .B(new_n336_), .Z(new_n337_));
  AOI21_X1  g136(.A(new_n285_), .B1(new_n333_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n331_), .A2(new_n300_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(new_n318_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT20), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT102), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n341_), .A2(KEYINPUT102), .A3(KEYINPUT20), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n344_), .A2(new_n327_), .A3(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(new_n288_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n320_), .A2(new_n325_), .A3(new_n289_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n337_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n284_), .B1(new_n339_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n333_), .A2(new_n337_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n337_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n352_), .B1(new_n326_), .B2(new_n332_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(KEYINPUT96), .A3(new_n353_), .ZN(new_n354_));
  OR3_X1    g153(.A1(new_n333_), .A2(KEYINPUT96), .A3(new_n337_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(new_n355_), .A3(new_n285_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n347_), .A2(new_n348_), .ZN(new_n357_));
  OAI211_X1 g156(.A(KEYINPUT103), .B(new_n338_), .C1(new_n357_), .C2(new_n337_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n283_), .A2(new_n350_), .A3(new_n356_), .A4(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n266_), .A2(new_n262_), .A3(new_n269_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n278_), .B1(new_n261_), .B2(new_n267_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT33), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n362_), .B1(new_n281_), .B2(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n364_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT100), .B(KEYINPUT33), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n281_), .A2(KEYINPUT101), .A3(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(KEYINPUT101), .B1(new_n281_), .B2(new_n366_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n337_), .A2(KEYINPUT32), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n370_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n371_), .B1(new_n370_), .B2(new_n333_), .ZN(new_n372_));
  AOI22_X1  g171(.A1(new_n365_), .A2(new_n369_), .B1(new_n372_), .B2(new_n282_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n257_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n359_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G71gat), .B(G99gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(G43gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n323_), .B(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G227gat), .A2(G233gat), .ZN(new_n379_));
  INV_X1    g178(.A(G15gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT30), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n378_), .B(new_n382_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n383_), .A2(KEYINPUT81), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(KEYINPUT81), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n260_), .B(KEYINPUT31), .ZN(new_n386_));
  OR3_X1    g185(.A1(new_n384_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n383_), .A2(KEYINPUT81), .A3(new_n386_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n350_), .A2(new_n356_), .A3(new_n257_), .A4(new_n358_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n389_), .A2(new_n282_), .ZN(new_n392_));
  AOI22_X1  g191(.A1(new_n375_), .A2(new_n389_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G229gat), .A2(G233gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n380_), .A2(KEYINPUT75), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT75), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(G15gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(G22gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT75), .B(G15gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(G22gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(G1gat), .ZN(new_n404_));
  INV_X1    g203(.A(G8gat), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT14), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n403_), .A2(new_n406_), .ZN(new_n407_));
  XOR2_X1   g206(.A(G1gat), .B(G8gat), .Z(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n403_), .A2(new_n408_), .A3(new_n406_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G29gat), .B(G36gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G43gat), .B(G50gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n413_), .A2(new_n415_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n417_), .A2(KEYINPUT77), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT77), .B1(new_n417_), .B2(new_n418_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n394_), .B1(new_n412_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n417_), .A2(new_n418_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT15), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n403_), .A2(new_n408_), .A3(new_n406_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n408_), .B1(new_n403_), .B2(new_n406_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT78), .B1(new_n425_), .B2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n423_), .B(KEYINPUT15), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT78), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n430_), .A2(new_n431_), .A3(new_n412_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n422_), .B1(new_n429_), .B2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n428_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n412_), .A2(new_n421_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n394_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  OR2_X1    g235(.A1(new_n433_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT79), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G113gat), .B(G141gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G169gat), .B(G197gat), .ZN(new_n441_));
  XOR2_X1   g240(.A(new_n440_), .B(new_n441_), .Z(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n439_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n437_), .A2(new_n438_), .A3(new_n442_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G99gat), .A2(G106gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT6), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT6), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(G99gat), .A3(G106gat), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n448_), .A2(new_n450_), .A3(KEYINPUT67), .ZN(new_n451_));
  AOI21_X1  g250(.A(KEYINPUT67), .B1(new_n448_), .B2(new_n450_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G85gat), .A2(G92gat), .ZN(new_n454_));
  AND2_X1   g253(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n455_));
  NOR2_X1   g254(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n454_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(G85gat), .ZN(new_n458_));
  INV_X1    g257(.A(G92gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n461_), .A2(KEYINPUT66), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(KEYINPUT66), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n457_), .B(new_n460_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n453_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT64), .ZN(new_n466_));
  OR2_X1    g265(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n466_), .B1(new_n469_), .B2(G106gat), .ZN(new_n470_));
  INV_X1    g269(.A(G106gat), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n467_), .A2(KEYINPUT64), .A3(new_n471_), .A4(new_n468_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n448_), .A2(new_n450_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT67), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT7), .ZN(new_n477_));
  INV_X1    g276(.A(G99gat), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(new_n478_), .A3(new_n471_), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n448_), .A2(new_n450_), .A3(KEYINPUT67), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n476_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n460_), .A2(new_n454_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT8), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n484_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n474_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(new_n485_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT8), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n465_), .A2(new_n473_), .B1(new_n489_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT35), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G232gat), .A2(G233gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  AOI22_X1  g296(.A1(new_n493_), .A2(new_n423_), .B1(new_n494_), .B2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n487_), .B1(new_n453_), .B2(new_n482_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n486_), .B1(new_n490_), .B2(new_n485_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT69), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT69), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n489_), .A2(new_n492_), .A3(new_n502_), .ZN(new_n503_));
  AOI22_X1  g302(.A1(new_n501_), .A2(new_n503_), .B1(new_n473_), .B2(new_n465_), .ZN(new_n504_));
  NOR3_X1   g303(.A1(new_n504_), .A2(KEYINPUT73), .A3(new_n425_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT73), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n473_), .A2(new_n453_), .A3(new_n464_), .ZN(new_n507_));
  NOR3_X1   g306(.A1(new_n499_), .A2(KEYINPUT69), .A3(new_n500_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n502_), .B1(new_n489_), .B2(new_n492_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n507_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n506_), .B1(new_n510_), .B2(new_n430_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n498_), .B1(new_n505_), .B2(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n497_), .A2(new_n494_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  OAI221_X1 g313(.A(new_n498_), .B1(new_n494_), .B2(new_n497_), .C1(new_n505_), .C2(new_n511_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(new_n515_), .A3(KEYINPUT74), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G190gat), .B(G218gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G134gat), .B(G162gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n519_), .A2(KEYINPUT36), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n516_), .A2(new_n521_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n514_), .A2(new_n515_), .A3(KEYINPUT74), .A4(new_n520_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n514_), .A2(new_n515_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n525_), .A2(KEYINPUT36), .A3(new_n519_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT37), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT71), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n507_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G57gat), .B(G64gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT11), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT68), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT11), .ZN(new_n534_));
  INV_X1    g333(.A(G57gat), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n535_), .A2(G64gat), .ZN(new_n536_));
  INV_X1    g335(.A(G64gat), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n537_), .A2(G57gat), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n534_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(G71gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(G78gat), .ZN(new_n541_));
  INV_X1    g340(.A(G78gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(G71gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n533_), .B1(new_n539_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n537_), .A2(G57gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n535_), .A2(G64gat), .ZN(new_n547_));
  AOI21_X1  g346(.A(KEYINPUT11), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G71gat), .B(G78gat), .ZN(new_n549_));
  NOR3_X1   g348(.A1(new_n548_), .A2(KEYINPUT68), .A3(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n532_), .B1(new_n545_), .B2(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(KEYINPUT68), .B1(new_n548_), .B2(new_n549_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n544_), .B(new_n533_), .C1(new_n531_), .C2(KEYINPUT11), .ZN(new_n553_));
  INV_X1    g352(.A(new_n532_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n551_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n530_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT12), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  AND2_X1   g358(.A1(G230gat), .A2(G233gat), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n554_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n560_), .B1(new_n493_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT70), .ZN(new_n565_));
  NOR3_X1   g364(.A1(new_n561_), .A2(new_n562_), .A3(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT70), .B1(new_n551_), .B2(new_n555_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT12), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n559_), .B(new_n564_), .C1(new_n568_), .C2(new_n504_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n493_), .A2(new_n563_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(new_n557_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(new_n560_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G120gat), .B(G148gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT5), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G176gat), .B(G204gat), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n574_), .B(new_n575_), .Z(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n569_), .A2(new_n572_), .A3(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n577_), .B1(new_n569_), .B2(new_n572_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n529_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n569_), .A2(new_n572_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n576_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n569_), .A2(new_n572_), .A3(new_n577_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(KEYINPUT71), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n580_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT13), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G127gat), .B(G155gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT16), .ZN(new_n589_));
  XOR2_X1   g388(.A(G183gat), .B(G211gat), .Z(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT17), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT76), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G231gat), .A2(G233gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n428_), .B(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(new_n563_), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n596_), .A2(new_n563_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n594_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n565_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n551_), .A2(KEYINPUT70), .A3(new_n555_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  AOI211_X1 g401(.A(new_n592_), .B(new_n591_), .C1(new_n596_), .C2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n603_), .B1(new_n602_), .B2(new_n596_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n599_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT37), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n524_), .A2(new_n607_), .A3(new_n526_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n528_), .A2(new_n587_), .A3(new_n606_), .A4(new_n608_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n393_), .A2(new_n446_), .A3(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT104), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n611_), .A2(new_n404_), .A3(new_n282_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT38), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n393_), .A2(new_n527_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n587_), .ZN(new_n616_));
  NOR3_X1   g415(.A1(new_n616_), .A2(new_n446_), .A3(new_n605_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n404_), .B1(new_n618_), .B2(new_n282_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n614_), .A2(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n620_), .B1(new_n613_), .B2(new_n612_), .ZN(G1324gat));
  INV_X1    g420(.A(KEYINPUT105), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n350_), .A2(new_n358_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(new_n356_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n618_), .A2(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n622_), .B1(new_n625_), .B2(G8gat), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n611_), .A2(new_n405_), .A3(new_n624_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  AOI211_X1 g429(.A(KEYINPUT105), .B(new_n405_), .C1(new_n618_), .C2(new_n624_), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n626_), .A2(new_n631_), .A3(new_n627_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT40), .ZN(G1325gat));
  INV_X1    g433(.A(new_n389_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n380_), .B1(new_n618_), .B2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT106), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n637_), .A2(KEYINPUT41), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(KEYINPUT41), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n611_), .A2(new_n380_), .A3(new_n635_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n638_), .A2(new_n639_), .A3(new_n640_), .ZN(G1326gat));
  AOI21_X1  g440(.A(new_n399_), .B1(new_n618_), .B2(new_n374_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT42), .Z(new_n643_));
  NAND3_X1  g442(.A1(new_n611_), .A2(new_n399_), .A3(new_n374_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(G1327gat));
  NOR2_X1   g444(.A1(new_n393_), .A2(new_n446_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n527_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n616_), .A2(new_n647_), .A3(new_n606_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(G29gat), .B1(new_n649_), .B2(new_n282_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n375_), .A2(new_n389_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n391_), .A2(new_n392_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n528_), .A2(new_n608_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT43), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT108), .B1(new_n653_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT108), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n393_), .A2(new_n659_), .A3(new_n656_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT107), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n654_), .B1(new_n393_), .B2(new_n662_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n651_), .A2(new_n662_), .A3(new_n652_), .ZN(new_n664_));
  OAI21_X1  g463(.A(KEYINPUT43), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n661_), .A2(new_n665_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n616_), .A2(new_n446_), .A3(new_n606_), .ZN(new_n667_));
  AOI21_X1  g466(.A(KEYINPUT44), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n669_));
  INV_X1    g468(.A(new_n667_), .ZN(new_n670_));
  AOI211_X1 g469(.A(new_n669_), .B(new_n670_), .C1(new_n661_), .C2(new_n665_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n668_), .A2(new_n671_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n282_), .A2(G29gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n650_), .B1(new_n672_), .B2(new_n673_), .ZN(G1328gat));
  INV_X1    g473(.A(G36gat), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n649_), .A2(new_n675_), .A3(new_n624_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT45), .Z(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n624_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n668_), .A2(new_n671_), .A3(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n678_), .B1(new_n680_), .B2(new_n675_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT46), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n678_), .B(KEYINPUT46), .C1(new_n675_), .C2(new_n680_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1329gat));
  NAND3_X1  g484(.A1(new_n672_), .A2(G43gat), .A3(new_n635_), .ZN(new_n686_));
  INV_X1    g485(.A(G43gat), .ZN(new_n687_));
  INV_X1    g486(.A(new_n649_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n687_), .B1(new_n688_), .B2(new_n389_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n686_), .A2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT47), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT47), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n686_), .A2(new_n692_), .A3(new_n689_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1330gat));
  AOI21_X1  g493(.A(G50gat), .B1(new_n649_), .B2(new_n374_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n374_), .A2(G50gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n672_), .B2(new_n696_), .ZN(G1331gat));
  NAND2_X1  g496(.A1(new_n653_), .A2(new_n446_), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n698_), .A2(KEYINPUT109), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(KEYINPUT109), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n699_), .A2(new_n616_), .A3(new_n700_), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n528_), .A2(new_n606_), .A3(new_n608_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n282_), .A2(new_n535_), .ZN(new_n704_));
  AND4_X1   g503(.A1(new_n446_), .A2(new_n615_), .A3(new_n616_), .A4(new_n606_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n705_), .A2(new_n282_), .ZN(new_n706_));
  OAI22_X1  g505(.A1(new_n703_), .A2(new_n704_), .B1(new_n535_), .B2(new_n706_), .ZN(G1332gat));
  AOI21_X1  g506(.A(new_n537_), .B1(new_n705_), .B2(new_n624_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n708_), .B(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n624_), .A2(new_n537_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n710_), .B1(new_n703_), .B2(new_n711_), .ZN(G1333gat));
  AOI21_X1  g511(.A(new_n540_), .B1(new_n705_), .B2(new_n635_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT49), .Z(new_n714_));
  NAND2_X1  g513(.A1(new_n635_), .A2(new_n540_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n714_), .B1(new_n703_), .B2(new_n715_), .ZN(G1334gat));
  AOI21_X1  g515(.A(new_n542_), .B1(new_n705_), .B2(new_n374_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT50), .Z(new_n718_));
  NAND2_X1  g517(.A1(new_n374_), .A2(new_n542_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n703_), .B2(new_n719_), .ZN(G1335gat));
  INV_X1    g519(.A(new_n446_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n587_), .A2(new_n721_), .A3(new_n606_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n666_), .A2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n282_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(G85gat), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n647_), .A2(new_n606_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n699_), .A2(new_n616_), .A3(new_n726_), .A4(new_n700_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n728_), .A2(new_n458_), .A3(new_n282_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n725_), .A2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT111), .ZN(G1336gat));
  NAND3_X1  g530(.A1(new_n728_), .A2(new_n459_), .A3(new_n624_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n723_), .A2(new_n624_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(new_n459_), .ZN(G1337gat));
  AOI21_X1  g533(.A(new_n478_), .B1(new_n723_), .B2(new_n635_), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n389_), .A2(new_n469_), .ZN(new_n736_));
  OAI21_X1  g535(.A(KEYINPUT112), .B1(new_n727_), .B2(new_n736_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n735_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT51), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n738_), .B(new_n739_), .ZN(G1338gat));
  NOR2_X1   g539(.A1(new_n257_), .A2(G106gat), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  OR3_X1    g541(.A1(new_n727_), .A2(KEYINPUT113), .A3(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(KEYINPUT113), .B1(new_n727_), .B2(new_n742_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n666_), .A2(new_n374_), .A3(new_n722_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(G106gat), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n746_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n745_), .A2(new_n749_), .A3(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT53), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT53), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n745_), .A2(new_n753_), .A3(new_n749_), .A4(new_n750_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(G1339gat));
  INV_X1    g554(.A(KEYINPUT119), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT57), .ZN(new_n757_));
  INV_X1    g556(.A(new_n394_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n758_), .B1(new_n412_), .B2(new_n421_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n429_), .B2(new_n432_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n758_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n443_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n442_), .B1(new_n433_), .B2(new_n436_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n580_), .A2(new_n584_), .A3(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT56), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n569_), .A2(KEYINPUT55), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT12), .B1(new_n530_), .B2(new_n556_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n558_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(new_n510_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT55), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n770_), .A2(new_n771_), .A3(new_n564_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n559_), .B(new_n570_), .C1(new_n568_), .C2(new_n504_), .ZN(new_n773_));
  AOI22_X1  g572(.A1(new_n767_), .A2(new_n772_), .B1(new_n560_), .B2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n766_), .B1(new_n774_), .B2(new_n577_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n577_), .A2(new_n766_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(KEYINPUT114), .B1(new_n774_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n773_), .A2(new_n560_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n569_), .A2(KEYINPUT55), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n771_), .B1(new_n770_), .B2(new_n564_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n779_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT114), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(new_n783_), .A3(new_n776_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n775_), .A2(new_n778_), .A3(new_n784_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n446_), .A2(new_n578_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n765_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n757_), .B1(new_n787_), .B2(new_n527_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT115), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT115), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n790_), .B(new_n757_), .C1(new_n787_), .C2(new_n527_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT118), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n775_), .B1(new_n774_), .B2(new_n777_), .ZN(new_n794_));
  OR2_X1    g593(.A1(KEYINPUT117), .A2(KEYINPUT58), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT116), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n764_), .A2(new_n796_), .A3(new_n583_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n764_), .B2(new_n583_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n794_), .A2(new_n795_), .A3(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n795_), .B1(new_n794_), .B2(new_n799_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n787_), .A2(new_n527_), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n803_), .A2(new_n654_), .B1(new_n804_), .B2(KEYINPUT57), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n792_), .A2(new_n793_), .A3(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n793_), .B1(new_n792_), .B2(new_n805_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n806_), .A2(new_n807_), .A3(new_n606_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n702_), .A2(new_n809_), .A3(new_n446_), .A4(new_n587_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT54), .B1(new_n609_), .B2(new_n721_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n756_), .B1(new_n808_), .B2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n792_), .A2(new_n805_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT118), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n792_), .A2(new_n805_), .A3(new_n793_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n605_), .A3(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n812_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(KEYINPUT119), .A3(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n813_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n391_), .A2(new_n282_), .A3(new_n635_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(G113gat), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n822_), .A2(new_n823_), .A3(new_n721_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n822_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n805_), .A2(new_n788_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n818_), .B1(new_n826_), .B2(new_n606_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n821_), .A2(KEYINPUT59), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n825_), .A2(KEYINPUT59), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n829_), .A2(new_n721_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n824_), .B1(new_n830_), .B2(new_n823_), .ZN(G1340gat));
  INV_X1    g630(.A(G120gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n832_), .B1(new_n587_), .B2(KEYINPUT60), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n822_), .B(new_n833_), .C1(KEYINPUT60), .C2(new_n832_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(KEYINPUT120), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n829_), .A2(new_n616_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(new_n832_), .ZN(G1341gat));
  INV_X1    g636(.A(G127gat), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n822_), .A2(new_n838_), .A3(new_n606_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n829_), .A2(new_n606_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(new_n838_), .ZN(G1342gat));
  INV_X1    g640(.A(G134gat), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n822_), .A2(new_n842_), .A3(new_n527_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n829_), .A2(new_n654_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(new_n842_), .ZN(G1343gat));
  AND4_X1   g644(.A1(new_n374_), .A2(new_n679_), .A3(new_n282_), .A4(new_n389_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n813_), .A2(new_n819_), .A3(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n813_), .A2(KEYINPUT121), .A3(new_n819_), .A4(new_n846_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n721_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n616_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(G148gat), .ZN(G1345gat));
  AOI21_X1  g654(.A(new_n606_), .B1(new_n814_), .B2(KEYINPUT118), .ZN(new_n856_));
  AOI211_X1 g655(.A(new_n756_), .B(new_n812_), .C1(new_n856_), .C2(new_n816_), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT119), .B1(new_n817_), .B2(new_n818_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(KEYINPUT121), .B1(new_n859_), .B2(new_n846_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n850_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n606_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT122), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT122), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n851_), .A2(new_n864_), .A3(new_n606_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(KEYINPUT61), .B(G155gat), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n863_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n866_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n864_), .B1(new_n851_), .B2(new_n606_), .ZN(new_n869_));
  AOI211_X1 g668(.A(KEYINPUT122), .B(new_n605_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n868_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n867_), .A2(new_n871_), .ZN(G1346gat));
  INV_X1    g671(.A(G162gat), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n851_), .A2(new_n873_), .A3(new_n527_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n851_), .A2(new_n654_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(new_n873_), .ZN(G1347gat));
  NAND2_X1  g675(.A1(new_n624_), .A2(new_n392_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(new_n374_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n827_), .A2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n721_), .ZN(new_n880_));
  OAI21_X1  g679(.A(KEYINPUT62), .B1(new_n880_), .B2(KEYINPUT22), .ZN(new_n881_));
  OAI21_X1  g680(.A(G169gat), .B1(new_n880_), .B2(KEYINPUT62), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n308_), .B2(new_n881_), .ZN(G1348gat));
  AOI21_X1  g683(.A(G176gat), .B1(new_n879_), .B2(new_n616_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n820_), .A2(new_n374_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n877_), .A2(new_n309_), .A3(new_n587_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n885_), .B1(new_n886_), .B2(new_n887_), .ZN(G1349gat));
  NAND4_X1  g687(.A1(new_n886_), .A2(new_n624_), .A3(new_n392_), .A4(new_n606_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n292_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n305_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n879_), .A2(new_n891_), .A3(new_n606_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(KEYINPUT123), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT123), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n890_), .A2(new_n895_), .A3(new_n892_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(G1350gat));
  AOI21_X1  g696(.A(new_n293_), .B1(new_n879_), .B2(new_n654_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(KEYINPUT124), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n879_), .A2(new_n303_), .A3(new_n527_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(G1351gat));
  NAND3_X1  g700(.A1(new_n624_), .A2(new_n283_), .A3(new_n389_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n820_), .A2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n721_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g704(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT125), .B(G204gat), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n903_), .A2(new_n616_), .ZN(new_n908_));
  MUX2_X1   g707(.A(new_n906_), .B(new_n907_), .S(new_n908_), .Z(G1353gat));
  NAND2_X1  g708(.A1(new_n903_), .A2(new_n606_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n911_));
  AND2_X1   g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n910_), .A2(new_n911_), .A3(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n910_), .A2(new_n911_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n910_), .A2(KEYINPUT126), .A3(new_n911_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n913_), .B1(new_n916_), .B2(new_n917_), .ZN(G1354gat));
  NOR3_X1   g717(.A1(new_n820_), .A2(new_n647_), .A3(new_n902_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT127), .ZN(new_n920_));
  OR2_X1    g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  AOI21_X1  g720(.A(G218gat), .B1(new_n919_), .B2(new_n920_), .ZN(new_n922_));
  AND2_X1   g721(.A1(new_n654_), .A2(G218gat), .ZN(new_n923_));
  AOI22_X1  g722(.A1(new_n921_), .A2(new_n922_), .B1(new_n903_), .B2(new_n923_), .ZN(G1355gat));
endmodule


