//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 0 0 1 1 1 1 0 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n683_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n832_, new_n833_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_;
  INV_X1    g000(.A(KEYINPUT78), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT26), .B(G190gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT77), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT76), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT25), .ZN(new_n206_));
  AOI21_X1  g005(.A(new_n205_), .B1(new_n206_), .B2(G183gat), .ZN(new_n207_));
  INV_X1    g006(.A(G183gat), .ZN(new_n208_));
  NOR3_X1   g007(.A1(new_n208_), .A2(KEYINPUT76), .A3(KEYINPUT25), .ZN(new_n209_));
  OAI22_X1  g008(.A1(new_n203_), .A2(new_n204_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT26), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(new_n204_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT75), .B(G183gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n213_), .B1(new_n214_), .B2(new_n206_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n202_), .B1(new_n210_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT26), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(G190gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n212_), .A2(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT76), .B1(new_n208_), .B2(KEYINPUT25), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n205_), .A2(new_n206_), .A3(G183gat), .ZN(new_n221_));
  AOI22_X1  g020(.A1(new_n219_), .A2(KEYINPUT77), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  AND2_X1   g021(.A1(KEYINPUT75), .A2(G183gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(KEYINPUT75), .A2(G183gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  AOI22_X1  g024(.A1(new_n225_), .A2(KEYINPUT25), .B1(new_n204_), .B2(new_n212_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n222_), .A2(new_n226_), .A3(KEYINPUT78), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT23), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n231_));
  INV_X1    g030(.A(G169gat), .ZN(new_n232_));
  INV_X1    g031(.A(G176gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n230_), .B(new_n231_), .C1(new_n234_), .C2(KEYINPUT24), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G169gat), .A2(G176gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n234_), .A2(KEYINPUT24), .A3(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT79), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n234_), .A2(KEYINPUT79), .A3(KEYINPUT24), .A4(new_n236_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n235_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n216_), .A2(new_n227_), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT81), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n230_), .A2(new_n231_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n244_), .B1(G190gat), .B2(new_n214_), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT80), .B1(new_n232_), .B2(KEYINPUT22), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT22), .B(G169gat), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n233_), .B(new_n246_), .C1(new_n247_), .C2(KEYINPUT80), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n245_), .A2(new_n248_), .A3(new_n236_), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n242_), .A2(new_n243_), .A3(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n243_), .B1(new_n242_), .B2(new_n249_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G71gat), .B(G99gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(G43gat), .ZN(new_n254_));
  XOR2_X1   g053(.A(new_n254_), .B(KEYINPUT30), .Z(new_n255_));
  XNOR2_X1  g054(.A(new_n252_), .B(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(KEYINPUT82), .B(G15gat), .Z(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT83), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G127gat), .B(G134gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G113gat), .B(G120gat), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n260_), .A2(new_n261_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n259_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT83), .B1(new_n260_), .B2(new_n261_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n266_), .B(KEYINPUT31), .Z(new_n267_));
  NAND2_X1  g066(.A1(G227gat), .A2(G233gat), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n267_), .B(new_n268_), .Z(new_n269_));
  XNOR2_X1  g068(.A(new_n258_), .B(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G8gat), .B(G36gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT18), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G64gat), .B(G92gat), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n272_), .B(new_n273_), .Z(new_n274_));
  XOR2_X1   g073(.A(new_n274_), .B(KEYINPUT101), .Z(new_n275_));
  INV_X1    g074(.A(new_n251_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n242_), .A2(new_n243_), .A3(new_n249_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT92), .ZN(new_n278_));
  INV_X1    g077(.A(G197gat), .ZN(new_n279_));
  INV_X1    g078(.A(G204gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT90), .B(G204gat), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n278_), .B(new_n281_), .C1(new_n282_), .C2(new_n279_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT91), .ZN(new_n285_));
  INV_X1    g084(.A(G218gat), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n286_), .A2(G211gat), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n286_), .A2(G211gat), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n285_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G211gat), .B(G218gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT91), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n289_), .A2(new_n291_), .A3(KEYINPUT21), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n284_), .A2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n281_), .B1(new_n282_), .B2(new_n279_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT92), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n282_), .A2(G197gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT89), .B1(new_n279_), .B2(G204gat), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT89), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(new_n280_), .A3(G197gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT21), .B1(new_n296_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT21), .ZN(new_n302_));
  AOI22_X1  g101(.A1(new_n294_), .A2(new_n302_), .B1(new_n289_), .B2(new_n291_), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n293_), .A2(new_n295_), .B1(new_n301_), .B2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n276_), .A2(new_n277_), .A3(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G226gat), .A2(G233gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT19), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT25), .B(G183gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT96), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(new_n203_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n235_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n312_), .A2(new_n237_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n244_), .B1(G183gat), .B2(G190gat), .ZN(new_n314_));
  INV_X1    g113(.A(new_n236_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n315_), .B1(new_n247_), .B2(new_n233_), .ZN(new_n316_));
  AOI22_X1  g115(.A1(new_n311_), .A2(new_n313_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT20), .B1(new_n304_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n305_), .A2(new_n308_), .A3(new_n319_), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n289_), .A2(new_n291_), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n321_), .A2(new_n295_), .A3(KEYINPUT21), .A4(new_n283_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n289_), .A2(new_n291_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n294_), .A2(new_n302_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n301_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n322_), .A2(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT20), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n328_), .B1(new_n304_), .B2(new_n317_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n308_), .B1(new_n327_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT99), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n320_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  AOI211_X1 g131(.A(KEYINPUT99), .B(new_n308_), .C1(new_n327_), .C2(new_n329_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n275_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  NOR3_X1   g133(.A1(new_n250_), .A2(new_n251_), .A3(new_n326_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n307_), .B1(new_n335_), .B2(new_n318_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n327_), .A2(new_n308_), .A3(new_n329_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(new_n274_), .A3(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n334_), .A2(KEYINPUT27), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT95), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G228gat), .A2(G233gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G78gat), .B(G106gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT93), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT1), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n344_), .A2(KEYINPUT84), .A3(G155gat), .A4(G162gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G141gat), .A2(G148gat), .ZN(new_n346_));
  INV_X1    g145(.A(G141gat), .ZN(new_n347_));
  INV_X1    g146(.A(G148gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n345_), .A2(new_n346_), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G155gat), .A2(G162gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT1), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n344_), .A2(G155gat), .A3(G162gat), .ZN(new_n353_));
  OR2_X1    g152(.A1(G155gat), .A2(G162gat), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT84), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .A4(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n350_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT3), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n358_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT2), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n346_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n359_), .A2(new_n361_), .A3(new_n362_), .A4(new_n363_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n354_), .A2(new_n351_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n357_), .A2(new_n366_), .ZN(new_n367_));
  AOI221_X4 g166(.A(new_n343_), .B1(new_n367_), .B2(KEYINPUT29), .C1(new_n322_), .C2(new_n325_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n343_), .ZN(new_n369_));
  AOI22_X1  g168(.A1(new_n350_), .A2(new_n356_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT29), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n369_), .B1(new_n326_), .B2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n341_), .B1(new_n368_), .B2(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n343_), .B1(new_n304_), .B2(new_n372_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n341_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n326_), .A2(new_n373_), .A3(new_n369_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n376_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n375_), .A2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G22gat), .B(G50gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT87), .B(KEYINPUT88), .ZN(new_n382_));
  XOR2_X1   g181(.A(new_n381_), .B(new_n382_), .Z(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT85), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n385_), .B1(new_n367_), .B2(KEYINPUT29), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n370_), .A2(KEYINPUT85), .A3(new_n371_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n386_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n388_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n384_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n386_), .A2(new_n387_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n388_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n395_), .A2(new_n389_), .A3(new_n383_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n392_), .A2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n340_), .B1(new_n380_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n375_), .A2(new_n379_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n392_), .A2(new_n396_), .ZN(new_n400_));
  NOR3_X1   g199(.A1(new_n399_), .A2(new_n400_), .A3(KEYINPUT95), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n399_), .A2(new_n400_), .A3(KEYINPUT94), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT94), .B1(new_n399_), .B2(new_n400_), .ZN(new_n403_));
  OAI22_X1  g202(.A1(new_n398_), .A2(new_n401_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n274_), .ZN(new_n405_));
  AND3_X1   g204(.A1(new_n327_), .A2(new_n308_), .A3(new_n329_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n308_), .B1(new_n305_), .B2(new_n319_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n405_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n338_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT27), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(KEYINPUT98), .B(KEYINPUT4), .Z(new_n412_));
  NAND4_X1  g211(.A1(new_n367_), .A2(new_n264_), .A3(new_n265_), .A4(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G225gat), .A2(G233gat), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n260_), .B(new_n261_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT97), .B1(new_n418_), .B2(new_n367_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n367_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT97), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n370_), .A2(new_n421_), .A3(new_n417_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n419_), .A2(new_n420_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT4), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n416_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n419_), .A2(new_n420_), .A3(new_n414_), .A4(new_n422_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G1gat), .B(G29gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(G85gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT0), .B(G57gat), .ZN(new_n430_));
  XOR2_X1   g229(.A(new_n429_), .B(new_n430_), .Z(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n427_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n425_), .A2(new_n426_), .A3(new_n431_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n339_), .A2(new_n404_), .A3(new_n411_), .A4(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n274_), .A2(KEYINPUT32), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n336_), .A2(new_n438_), .A3(new_n337_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n439_), .A2(new_n435_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n438_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n441_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT33), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n434_), .A2(new_n444_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n425_), .A2(KEYINPUT33), .A3(new_n426_), .A4(new_n431_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n414_), .B(new_n413_), .C1(new_n423_), .C2(new_n424_), .ZN(new_n447_));
  OAI211_X1 g246(.A(new_n447_), .B(new_n432_), .C1(new_n414_), .C2(new_n423_), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n445_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(new_n338_), .A3(new_n408_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n404_), .B1(new_n443_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT100), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n437_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  AOI211_X1 g252(.A(KEYINPUT100), .B(new_n404_), .C1(new_n443_), .C2(new_n450_), .ZN(new_n454_));
  OAI211_X1 g253(.A(KEYINPUT102), .B(new_n270_), .C1(new_n453_), .C2(new_n454_), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n339_), .A2(new_n411_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n404_), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n270_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(new_n436_), .A3(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n455_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n409_), .ZN(new_n462_));
  AOI22_X1  g261(.A1(new_n462_), .A2(new_n449_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT100), .B1(new_n463_), .B2(new_n404_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n451_), .A2(new_n452_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(new_n465_), .A3(new_n437_), .ZN(new_n466_));
  AOI21_X1  g265(.A(KEYINPUT102), .B1(new_n466_), .B2(new_n270_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n461_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G29gat), .B(G36gat), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT67), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G43gat), .B(G50gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT15), .ZN(new_n474_));
  XOR2_X1   g273(.A(G85gat), .B(G92gat), .Z(new_n475_));
  NOR2_X1   g274(.A1(G99gat), .A2(G106gat), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT7), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G99gat), .A2(G106gat), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n475_), .B1(new_n478_), .B2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT8), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT64), .B(G92gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(G85gat), .ZN(new_n486_));
  OR3_X1    g285(.A1(new_n485_), .A2(KEYINPUT9), .A3(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n481_), .B1(KEYINPUT9), .B2(new_n475_), .ZN(new_n488_));
  XOR2_X1   g287(.A(KEYINPUT10), .B(G99gat), .Z(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n487_), .B(new_n488_), .C1(G106gat), .C2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n483_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT65), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT65), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n483_), .A2(new_n494_), .A3(new_n491_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n474_), .A2(new_n493_), .A3(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G232gat), .A2(G233gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT34), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n483_), .A2(new_n473_), .A3(new_n491_), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n499_), .A2(KEYINPUT68), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(KEYINPUT68), .ZN(new_n501_));
  OAI221_X1 g300(.A(new_n496_), .B1(KEYINPUT35), .B2(new_n498_), .C1(new_n500_), .C2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n498_), .A2(KEYINPUT35), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G190gat), .B(G218gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G134gat), .B(G162gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT36), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n504_), .A2(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n507_), .A2(KEYINPUT36), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n504_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n468_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT103), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n514_), .A2(KEYINPUT103), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G57gat), .B(G64gat), .ZN(new_n519_));
  OR2_X1    g318(.A1(new_n519_), .A2(KEYINPUT11), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(KEYINPUT11), .ZN(new_n521_));
  XOR2_X1   g320(.A(G71gat), .B(G78gat), .Z(new_n522_));
  NAND3_X1  g321(.A1(new_n520_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n521_), .A2(new_n522_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n483_), .A2(new_n491_), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT12), .ZN(new_n528_));
  INV_X1    g327(.A(new_n525_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n492_), .A2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n527_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G230gat), .A2(G233gat), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n493_), .A2(KEYINPUT12), .A3(new_n495_), .A4(new_n529_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n530_), .A2(new_n526_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n534_), .B1(new_n532_), .B2(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(G120gat), .B(G148gat), .Z(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT66), .B(KEYINPUT5), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G176gat), .B(G204gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n536_), .B(new_n542_), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n543_), .A2(KEYINPUT13), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(KEYINPUT13), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(G15gat), .B(G22gat), .Z(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT69), .B(G8gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(G1gat), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n548_), .B1(new_n550_), .B2(KEYINPUT14), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT70), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G1gat), .B(G8gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT70), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n551_), .B(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n553_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n554_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n473_), .ZN(new_n560_));
  OR3_X1    g359(.A1(new_n559_), .A2(KEYINPUT72), .A3(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT72), .B1(new_n559_), .B2(new_n560_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G229gat), .A2(G233gat), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n474_), .A2(new_n559_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT73), .ZN(new_n567_));
  AOI22_X1  g366(.A1(new_n561_), .A2(new_n562_), .B1(new_n560_), .B2(new_n559_), .ZN(new_n568_));
  OAI22_X1  g367(.A1(new_n565_), .A2(new_n567_), .B1(new_n568_), .B2(new_n564_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G113gat), .B(G141gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G169gat), .B(G197gat), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n570_), .B(new_n571_), .Z(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n569_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT74), .ZN(new_n575_));
  OAI221_X1 g374(.A(new_n572_), .B1(new_n568_), .B2(new_n564_), .C1(new_n565_), .C2(new_n567_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n574_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n569_), .A2(KEYINPUT74), .A3(new_n573_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G231gat), .A2(G233gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n525_), .B(new_n580_), .Z(new_n581_));
  XNOR2_X1  g380(.A(new_n559_), .B(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(G127gat), .B(G155gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT71), .B(KEYINPUT16), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G183gat), .B(G211gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n582_), .A2(KEYINPUT17), .A3(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(KEYINPUT17), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n582_), .A2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n547_), .A2(new_n579_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n518_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(G1gat), .B1(new_n596_), .B2(new_n436_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n468_), .A2(new_n579_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT37), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n512_), .B(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n600_), .A2(new_n592_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n598_), .A2(new_n546_), .A3(new_n601_), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n602_), .A2(G1gat), .A3(new_n436_), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n603_), .B(KEYINPUT38), .Z(new_n604_));
  NAND2_X1  g403(.A1(new_n597_), .A2(new_n604_), .ZN(G1324gat));
  OR3_X1    g404(.A1(new_n602_), .A2(new_n456_), .A3(new_n549_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n456_), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n607_), .B(new_n593_), .C1(new_n516_), .C2(new_n517_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT39), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n608_), .A2(new_n609_), .A3(G8gat), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n609_), .B1(new_n608_), .B2(G8gat), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n606_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT40), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  OAI211_X1 g413(.A(KEYINPUT40), .B(new_n606_), .C1(new_n610_), .C2(new_n611_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(G1325gat));
  INV_X1    g415(.A(G15gat), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n617_), .B1(new_n595_), .B2(new_n459_), .ZN(new_n618_));
  XOR2_X1   g417(.A(KEYINPUT104), .B(KEYINPUT41), .Z(new_n619_));
  OR2_X1    g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n619_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n459_), .A2(new_n617_), .ZN(new_n622_));
  OAI211_X1 g421(.A(new_n620_), .B(new_n621_), .C1(new_n602_), .C2(new_n622_), .ZN(G1326gat));
  NAND2_X1  g422(.A1(new_n595_), .A2(new_n404_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT42), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n624_), .A2(new_n625_), .A3(G22gat), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n625_), .B1(new_n624_), .B2(G22gat), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n457_), .A2(G22gat), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT105), .Z(new_n629_));
  OAI22_X1  g428(.A1(new_n626_), .A2(new_n627_), .B1(new_n602_), .B2(new_n629_), .ZN(G1327gat));
  NOR2_X1   g429(.A1(new_n512_), .A2(new_n591_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n632_), .A2(new_n547_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n598_), .A2(new_n633_), .ZN(new_n634_));
  OR3_X1    g433(.A1(new_n634_), .A2(G29gat), .A3(new_n436_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT107), .ZN(new_n636_));
  INV_X1    g435(.A(new_n579_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n637_), .A2(new_n546_), .A3(new_n592_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n600_), .B1(new_n461_), .B2(new_n467_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT43), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n642_), .B(new_n600_), .C1(new_n461_), .C2(new_n467_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n638_), .B1(new_n641_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT44), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n636_), .B1(new_n646_), .B2(new_n435_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n638_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n643_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n640_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n270_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT102), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n653_), .A2(new_n460_), .A3(new_n455_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n650_), .B1(new_n654_), .B2(new_n600_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n648_), .B1(new_n649_), .B2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(new_n645_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n644_), .A2(KEYINPUT44), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n657_), .A2(new_n658_), .A3(new_n636_), .A4(new_n435_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(G29gat), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n635_), .B1(new_n647_), .B2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT108), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT108), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n663_), .B(new_n635_), .C1(new_n647_), .C2(new_n660_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(G1328gat));
  NAND3_X1  g464(.A1(new_n657_), .A2(new_n607_), .A3(new_n658_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(G36gat), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT45), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n456_), .A2(G36gat), .ZN(new_n669_));
  OR3_X1    g468(.A1(new_n634_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n668_), .B1(new_n634_), .B2(new_n669_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT109), .B1(new_n667_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT46), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(G1329gat));
  NAND3_X1  g474(.A1(new_n646_), .A2(G43gat), .A3(new_n459_), .ZN(new_n676_));
  INV_X1    g475(.A(G43gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n677_), .B1(new_n634_), .B2(new_n270_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g479(.A(G50gat), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n457_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n598_), .A2(new_n404_), .A3(new_n633_), .ZN(new_n683_));
  AOI22_X1  g482(.A1(new_n646_), .A2(new_n682_), .B1(new_n681_), .B2(new_n683_), .ZN(G1331gat));
  NOR2_X1   g483(.A1(new_n468_), .A2(new_n637_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT110), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n686_), .A2(new_n547_), .A3(new_n601_), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n687_), .A2(KEYINPUT111), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(KEYINPUT111), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n436_), .A2(G57gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n688_), .A2(new_n689_), .A3(new_n690_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n637_), .A2(new_n546_), .A3(new_n592_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n692_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n693_));
  OAI21_X1  g492(.A(G57gat), .B1(new_n693_), .B2(new_n436_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n691_), .A2(new_n694_), .ZN(G1332gat));
  NOR2_X1   g494(.A1(new_n456_), .A2(G64gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n688_), .A2(new_n689_), .A3(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(G64gat), .B1(new_n693_), .B2(new_n456_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n698_), .A2(KEYINPUT48), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n698_), .A2(KEYINPUT48), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n697_), .B1(new_n699_), .B2(new_n700_), .ZN(G1333gat));
  NOR2_X1   g500(.A1(new_n270_), .A2(G71gat), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n688_), .A2(new_n689_), .A3(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(G71gat), .B1(new_n693_), .B2(new_n270_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n704_), .A2(KEYINPUT49), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(KEYINPUT49), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n703_), .B1(new_n705_), .B2(new_n706_), .ZN(G1334gat));
  NOR2_X1   g506(.A1(new_n457_), .A2(G78gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n688_), .A2(new_n689_), .A3(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G78gat), .B1(new_n693_), .B2(new_n457_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n710_), .A2(KEYINPUT50), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(KEYINPUT50), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n709_), .B1(new_n711_), .B2(new_n712_), .ZN(G1335gat));
  NAND2_X1  g512(.A1(new_n686_), .A2(new_n547_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n714_), .A2(new_n632_), .ZN(new_n715_));
  AOI21_X1  g514(.A(G85gat), .B1(new_n715_), .B2(new_n435_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n547_), .A2(new_n592_), .A3(new_n579_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n717_), .B1(new_n641_), .B2(new_n643_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT112), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n436_), .A2(new_n486_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n716_), .B1(new_n719_), .B2(new_n720_), .ZN(G1336gat));
  AOI21_X1  g520(.A(G92gat), .B1(new_n715_), .B2(new_n607_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n456_), .A2(new_n485_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n719_), .B2(new_n723_), .ZN(G1337gat));
  INV_X1    g523(.A(KEYINPUT113), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT51), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT114), .Z(new_n727_));
  NOR4_X1   g526(.A1(new_n714_), .A2(new_n490_), .A3(new_n270_), .A4(new_n632_), .ZN(new_n728_));
  INV_X1    g527(.A(G99gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n729_), .B1(new_n718_), .B2(new_n459_), .ZN(new_n730_));
  OAI221_X1 g529(.A(new_n727_), .B1(new_n725_), .B2(KEYINPUT51), .C1(new_n728_), .C2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n727_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n270_), .A2(new_n490_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n730_), .B1(new_n715_), .B2(new_n733_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n725_), .A2(KEYINPUT51), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n732_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n731_), .A2(new_n736_), .ZN(G1338gat));
  NOR2_X1   g536(.A1(new_n457_), .A2(G106gat), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n686_), .A2(new_n547_), .A3(new_n631_), .A4(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n717_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n404_), .B(new_n740_), .C1(new_n649_), .C2(new_n655_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT115), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n741_), .A2(new_n742_), .A3(G106gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n741_), .B2(G106gat), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n743_), .A2(new_n744_), .A3(KEYINPUT52), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n746_));
  AOI211_X1 g545(.A(new_n457_), .B(new_n717_), .C1(new_n641_), .C2(new_n643_), .ZN(new_n747_));
  INV_X1    g546(.A(G106gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(KEYINPUT115), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n741_), .A2(new_n742_), .A3(G106gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n739_), .B1(new_n745_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT53), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT53), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n754_), .B(new_n739_), .C1(new_n745_), .C2(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1339gat));
  NAND3_X1  g555(.A1(new_n458_), .A2(new_n435_), .A3(new_n459_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT120), .ZN(new_n758_));
  INV_X1    g557(.A(new_n564_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n563_), .A2(new_n759_), .ZN(new_n760_));
  OAI221_X1 g559(.A(new_n573_), .B1(new_n568_), .B2(new_n759_), .C1(new_n760_), .C2(new_n567_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n543_), .A2(KEYINPUT116), .A3(new_n576_), .A4(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n543_), .A2(new_n576_), .A3(new_n761_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT116), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n536_), .A2(new_n542_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n577_), .A2(new_n766_), .A3(new_n578_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n532_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n534_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n531_), .A2(new_n533_), .A3(KEYINPUT55), .A4(new_n532_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n541_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT56), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n772_), .B(new_n773_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n762_), .B(new_n765_), .C1(new_n767_), .C2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n512_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT57), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n758_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n775_), .A2(KEYINPUT120), .A3(KEYINPUT57), .A4(new_n512_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n512_), .B(KEYINPUT37), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT58), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n770_), .A2(new_n771_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n542_), .ZN(new_n784_));
  OAI21_X1  g583(.A(KEYINPUT117), .B1(new_n784_), .B2(new_n773_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT118), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n784_), .A2(new_n786_), .A3(new_n773_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT117), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n772_), .A2(new_n788_), .A3(KEYINPUT56), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT118), .B1(new_n772_), .B2(KEYINPUT56), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n785_), .A2(new_n787_), .A3(new_n789_), .A4(new_n790_), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n576_), .A2(new_n761_), .A3(new_n766_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n782_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n791_), .A2(new_n792_), .A3(new_n782_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n781_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT119), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n780_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n776_), .A2(new_n777_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n799_), .B1(new_n796_), .B2(KEYINPUT119), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n592_), .B1(new_n798_), .B2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n781_), .A2(new_n591_), .A3(new_n546_), .ZN(new_n802_));
  OAI21_X1  g601(.A(KEYINPUT54), .B1(new_n802_), .B2(new_n637_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n601_), .A2(new_n804_), .A3(new_n546_), .A4(new_n579_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n803_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n757_), .B1(new_n801_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT59), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n791_), .A2(new_n792_), .A3(new_n782_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n600_), .B1(new_n810_), .B2(new_n793_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n799_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT121), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT121), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n811_), .A2(new_n799_), .A3(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n813_), .A2(new_n780_), .A3(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n806_), .B1(new_n816_), .B2(new_n592_), .ZN(new_n817_));
  OR2_X1    g616(.A1(new_n757_), .A2(KEYINPUT59), .ZN(new_n818_));
  OAI22_X1  g617(.A1(new_n808_), .A2(new_n809_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(G113gat), .B1(new_n819_), .B2(new_n579_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n808_), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n579_), .A2(G113gat), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n820_), .B1(new_n821_), .B2(new_n822_), .ZN(G1340gat));
  INV_X1    g622(.A(KEYINPUT60), .ZN(new_n824_));
  AOI21_X1  g623(.A(G120gat), .B1(new_n547_), .B2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n825_), .B1(new_n824_), .B2(G120gat), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n808_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT122), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n827_), .B(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(G120gat), .B1(new_n819_), .B2(new_n546_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(G1341gat));
  OAI21_X1  g630(.A(G127gat), .B1(new_n819_), .B2(new_n592_), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n592_), .A2(G127gat), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n832_), .B1(new_n821_), .B2(new_n833_), .ZN(G1342gat));
  OAI21_X1  g633(.A(G134gat), .B1(new_n819_), .B2(new_n781_), .ZN(new_n835_));
  OR2_X1    g634(.A1(new_n512_), .A2(G134gat), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n821_), .B2(new_n836_), .ZN(G1343gat));
  AOI21_X1  g636(.A(new_n459_), .B1(new_n801_), .B2(new_n807_), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n607_), .A2(new_n436_), .A3(new_n457_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n840_), .A2(new_n579_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(new_n347_), .ZN(G1344gat));
  NOR2_X1   g641(.A1(new_n840_), .A2(new_n546_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(new_n348_), .ZN(G1345gat));
  NAND3_X1  g643(.A1(new_n838_), .A2(new_n591_), .A3(new_n839_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(KEYINPUT61), .B(G155gat), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n845_), .B(new_n846_), .ZN(G1346gat));
  OAI21_X1  g646(.A(G162gat), .B1(new_n840_), .B2(new_n781_), .ZN(new_n848_));
  INV_X1    g647(.A(G162gat), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n513_), .A2(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n848_), .B1(new_n840_), .B2(new_n850_), .ZN(G1347gat));
  NOR3_X1   g650(.A1(new_n270_), .A2(new_n456_), .A3(new_n435_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(new_n404_), .ZN(new_n854_));
  AOI22_X1  g653(.A1(new_n812_), .A2(KEYINPUT121), .B1(new_n778_), .B2(new_n779_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n591_), .B1(new_n855_), .B2(new_n815_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n637_), .B(new_n854_), .C1(new_n856_), .C2(new_n806_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(G169gat), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT123), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n857_), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(KEYINPUT62), .A3(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n247_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n857_), .A2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(KEYINPUT123), .B1(new_n857_), .B2(G169gat), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT62), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n864_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n862_), .A2(new_n867_), .ZN(G1348gat));
  INV_X1    g667(.A(new_n854_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n817_), .A2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(G176gat), .B1(new_n870_), .B2(new_n547_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n404_), .B1(new_n801_), .B2(new_n807_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n853_), .A2(new_n233_), .A3(new_n546_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n871_), .B1(new_n872_), .B2(new_n873_), .ZN(G1349gat));
  NOR2_X1   g673(.A1(new_n592_), .A2(new_n310_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n870_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n853_), .A2(new_n592_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n214_), .B1(new_n872_), .B2(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(KEYINPUT124), .B1(new_n877_), .B2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n872_), .A2(new_n878_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n881_), .B(new_n876_), .C1(new_n882_), .C2(new_n214_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n880_), .A2(new_n883_), .ZN(G1350gat));
  NOR2_X1   g683(.A1(new_n512_), .A2(new_n219_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n870_), .A2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n211_), .B1(new_n870_), .B2(new_n600_), .ZN(new_n888_));
  OAI21_X1  g687(.A(KEYINPUT125), .B1(new_n887_), .B2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT125), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n817_), .A2(new_n781_), .A3(new_n869_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n886_), .B(new_n890_), .C1(new_n211_), .C2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n889_), .A2(new_n892_), .ZN(G1351gat));
  NAND2_X1  g692(.A1(new_n404_), .A2(new_n436_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n456_), .A2(new_n894_), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n838_), .A2(G197gat), .A3(new_n637_), .A4(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT126), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n896_), .A2(new_n897_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n895_), .ZN(new_n900_));
  AOI211_X1 g699(.A(new_n459_), .B(new_n900_), .C1(new_n801_), .C2(new_n807_), .ZN(new_n901_));
  AOI21_X1  g700(.A(G197gat), .B1(new_n901_), .B2(new_n637_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n898_), .A2(new_n899_), .A3(new_n902_), .ZN(G1352gat));
  INV_X1    g702(.A(new_n901_), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n904_), .A2(new_n282_), .A3(new_n546_), .ZN(new_n905_));
  AOI21_X1  g704(.A(G204gat), .B1(new_n901_), .B2(new_n547_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1353gat));
  XNOR2_X1  g706(.A(KEYINPUT63), .B(G211gat), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n904_), .A2(new_n592_), .A3(new_n908_), .ZN(new_n909_));
  AOI211_X1 g708(.A(KEYINPUT63), .B(G211gat), .C1(new_n901_), .C2(new_n591_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1354gat));
  OAI21_X1  g710(.A(G218gat), .B1(new_n904_), .B2(new_n781_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n901_), .A2(new_n286_), .A3(new_n513_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1355gat));
endmodule


