//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 0 1 0 0 0 1 1 1 0 1 1 0 1 0 0 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n913_, new_n914_, new_n916_, new_n917_, new_n918_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_;
  INV_X1    g000(.A(KEYINPUT23), .ZN(new_n202_));
  AOI21_X1  g001(.A(new_n202_), .B1(G183gat), .B2(G190gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT84), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n203_), .B1(new_n205_), .B2(new_n202_), .ZN(new_n206_));
  NOR3_X1   g005(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT85), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT25), .B(G183gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT26), .B(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G169gat), .ZN(new_n215_));
  INV_X1    g014(.A(G176gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  AND2_X1   g016(.A1(new_n212_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n209_), .A2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n208_), .A2(KEYINPUT85), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n222_), .B1(new_n205_), .B2(KEYINPUT23), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n223_), .B1(G183gat), .B2(G190gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(G169gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n221_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G227gat), .A2(G233gat), .ZN(new_n229_));
  INV_X1    g028(.A(G15gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n228_), .B(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(new_n232_), .B(KEYINPUT31), .Z(new_n233_));
  XNOR2_X1  g032(.A(G71gat), .B(G99gat), .ZN(new_n234_));
  INV_X1    g033(.A(G43gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT86), .B(KEYINPUT30), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(G127gat), .B(G134gat), .Z(new_n239_));
  XOR2_X1   g038(.A(G113gat), .B(G120gat), .Z(new_n240_));
  XOR2_X1   g039(.A(new_n239_), .B(new_n240_), .Z(new_n241_));
  XNOR2_X1  g040(.A(new_n238_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n233_), .B(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(G141gat), .A2(G148gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT3), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G141gat), .A2(G148gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT2), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT87), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G155gat), .A2(G162gat), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(G155gat), .A2(G162gat), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n250_), .A2(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n253_), .B1(KEYINPUT1), .B2(new_n251_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n257_), .B1(KEYINPUT1), .B2(new_n251_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n244_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(new_n259_), .A3(new_n246_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n256_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT29), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(G228gat), .ZN(new_n265_));
  INV_X1    g064(.A(G233gat), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(G204gat), .ZN(new_n268_));
  OR3_X1    g067(.A1(new_n268_), .A2(KEYINPUT89), .A3(G197gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT89), .B1(new_n268_), .B2(G197gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT88), .B(G204gat), .ZN(new_n271_));
  INV_X1    g070(.A(G197gat), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n269_), .B(new_n270_), .C1(new_n271_), .C2(new_n272_), .ZN(new_n273_));
  OR2_X1    g072(.A1(new_n273_), .A2(KEYINPUT21), .ZN(new_n274_));
  XOR2_X1   g073(.A(G211gat), .B(G218gat), .Z(new_n275_));
  OR2_X1    g074(.A1(new_n271_), .A2(G197gat), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT21), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n277_), .B1(G197gat), .B2(G204gat), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n275_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n275_), .A2(KEYINPUT21), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n274_), .A2(new_n279_), .B1(new_n273_), .B2(new_n280_), .ZN(new_n281_));
  OR3_X1    g080(.A1(new_n264_), .A2(new_n267_), .A3(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n267_), .B1(new_n264_), .B2(new_n281_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G78gat), .B(G106gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT90), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n282_), .A2(new_n283_), .A3(new_n285_), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n286_), .A2(KEYINPUT91), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n262_), .A2(new_n263_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT28), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G22gat), .B(G50gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n286_), .A2(KEYINPUT91), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n282_), .A2(new_n283_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n284_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n287_), .A2(new_n291_), .A3(new_n292_), .A4(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n290_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n289_), .B(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n285_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n286_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n297_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n295_), .A2(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n241_), .B1(new_n256_), .B2(new_n261_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT93), .ZN(new_n303_));
  INV_X1    g102(.A(new_n241_), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n304_), .B(new_n260_), .C1(new_n250_), .C2(new_n255_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n302_), .A2(new_n303_), .A3(new_n305_), .ZN(new_n306_));
  OAI211_X1 g105(.A(KEYINPUT93), .B(new_n241_), .C1(new_n256_), .C2(new_n261_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT4), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT94), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G225gat), .A2(G233gat), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n312_), .B(KEYINPUT95), .Z(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT96), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n308_), .A2(KEYINPUT94), .A3(KEYINPUT4), .ZN(new_n315_));
  OR2_X1    g114(.A1(new_n302_), .A2(KEYINPUT4), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n311_), .A2(new_n314_), .A3(new_n315_), .A4(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n308_), .A2(new_n313_), .ZN(new_n318_));
  XOR2_X1   g117(.A(G1gat), .B(G29gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT97), .B(G85gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT0), .B(G57gat), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n321_), .B(new_n322_), .Z(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n317_), .A2(new_n318_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT33), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT98), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G8gat), .B(G36gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT18), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G64gat), .B(G92gat), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n330_), .B(new_n331_), .Z(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n281_), .B1(new_n221_), .B2(new_n227_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G226gat), .A2(G233gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT19), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n210_), .B(KEYINPUT92), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n211_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n207_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n338_), .A2(new_n223_), .A3(new_n339_), .A4(new_n217_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(G183gat), .A2(G190gat), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n226_), .B1(new_n206_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n281_), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT20), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NOR3_X1   g144(.A1(new_n334_), .A2(new_n336_), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT20), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n347_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n227_), .B(new_n281_), .C1(new_n219_), .C2(new_n220_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n336_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n333_), .B1(new_n346_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n336_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n345_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n354_), .B(new_n355_), .C1(new_n228_), .C2(new_n281_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n356_), .A2(new_n332_), .A3(new_n351_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n353_), .A2(new_n357_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n311_), .A2(new_n313_), .A3(new_n315_), .A4(new_n316_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n324_), .B1(new_n308_), .B2(new_n314_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n358_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n317_), .A2(KEYINPUT33), .A3(new_n318_), .A4(new_n324_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT98), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n325_), .A2(new_n364_), .A3(new_n326_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n328_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n317_), .A2(new_n318_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(new_n323_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(new_n325_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n332_), .A2(KEYINPUT32), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NOR3_X1   g170(.A1(new_n346_), .A2(new_n352_), .A3(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n336_), .B1(new_n334_), .B2(new_n345_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT99), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n348_), .A2(new_n349_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n354_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT100), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n375_), .A2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n372_), .B1(new_n380_), .B2(new_n371_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n369_), .A2(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n301_), .B1(new_n366_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT27), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n358_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT101), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT101), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n358_), .A2(new_n387_), .A3(new_n384_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n380_), .A2(new_n333_), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n357_), .A2(KEYINPUT27), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n389_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n301_), .ZN(new_n394_));
  NOR3_X1   g193(.A1(new_n393_), .A2(new_n394_), .A3(new_n369_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n243_), .B1(new_n383_), .B2(new_n395_), .ZN(new_n396_));
  NOR4_X1   g195(.A1(new_n243_), .A2(new_n393_), .A3(new_n301_), .A4(new_n369_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(G85gat), .ZN(new_n400_));
  INV_X1    g199(.A(G92gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT9), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G85gat), .A2(G92gat), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT64), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n402_), .B(new_n403_), .C1(new_n405_), .C2(new_n406_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n402_), .A2(KEYINPUT64), .A3(KEYINPUT9), .A4(new_n404_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G99gat), .A2(G106gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT6), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT6), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(G99gat), .A3(G106gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  OR2_X1    g212(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n414_));
  INV_X1    g213(.A(G106gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n414_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n407_), .A2(new_n408_), .A3(new_n413_), .A4(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT65), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  AND2_X1   g219(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n421_));
  NOR2_X1   g220(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n423_), .A2(new_n415_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n424_), .A2(KEYINPUT65), .A3(new_n407_), .A4(new_n408_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n420_), .A2(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n402_), .A2(new_n404_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n410_), .A2(new_n412_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT7), .ZN(new_n429_));
  INV_X1    g228(.A(G99gat), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n429_), .A2(new_n430_), .A3(new_n415_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n427_), .B1(new_n428_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT8), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n413_), .A2(new_n432_), .A3(new_n431_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT8), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n437_), .A3(new_n427_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n426_), .B1(new_n435_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G57gat), .B(G64gat), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n441_), .A2(KEYINPUT11), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(KEYINPUT11), .ZN(new_n443_));
  XOR2_X1   g242(.A(G71gat), .B(G78gat), .Z(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n443_), .A2(new_n444_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n440_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT66), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n439_), .A2(new_n447_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G230gat), .A2(G233gat), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n452_), .B(new_n454_), .C1(new_n450_), .C2(new_n449_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n436_), .A2(new_n437_), .A3(new_n427_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n437_), .B1(new_n436_), .B2(new_n427_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT67), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT67), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n435_), .A2(new_n459_), .A3(new_n438_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n426_), .ZN(new_n462_));
  AOI21_X1  g261(.A(KEYINPUT68), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT68), .ZN(new_n464_));
  AOI211_X1 g263(.A(new_n464_), .B(new_n426_), .C1(new_n458_), .C2(new_n460_), .ZN(new_n465_));
  OAI211_X1 g264(.A(KEYINPUT12), .B(new_n448_), .C1(new_n463_), .C2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n451_), .A2(KEYINPUT12), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(new_n449_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n466_), .A2(new_n468_), .A3(new_n453_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n455_), .A2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G120gat), .B(G148gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT5), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G176gat), .B(G204gat), .ZN(new_n473_));
  XOR2_X1   g272(.A(new_n472_), .B(new_n473_), .Z(new_n474_));
  NAND2_X1  g273(.A1(new_n470_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n474_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n455_), .A2(new_n469_), .A3(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT13), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n475_), .A2(KEYINPUT13), .A3(new_n477_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G29gat), .B(G36gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G43gat), .B(G50gat), .ZN(new_n484_));
  XOR2_X1   g283(.A(new_n483_), .B(new_n484_), .Z(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT15), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G15gat), .B(G22gat), .ZN(new_n488_));
  INV_X1    g287(.A(G1gat), .ZN(new_n489_));
  INV_X1    g288(.A(G8gat), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT14), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G1gat), .B(G8gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n487_), .A2(KEYINPUT81), .A3(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n485_), .B(KEYINPUT80), .Z(new_n496_));
  INV_X1    g295(.A(new_n494_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT81), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n499_), .B1(new_n486_), .B2(new_n497_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n495_), .A2(new_n498_), .A3(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G229gat), .A2(G233gat), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n502_), .B(KEYINPUT82), .Z(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  OR3_X1    g303(.A1(new_n501_), .A2(KEYINPUT83), .A3(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT83), .B1(new_n501_), .B2(new_n504_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n496_), .B(new_n497_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n507_), .A2(G229gat), .A3(G233gat), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n505_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G113gat), .B(G141gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G169gat), .B(G197gat), .ZN(new_n511_));
  XOR2_X1   g310(.A(new_n510_), .B(new_n511_), .Z(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n509_), .A2(new_n513_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n505_), .A2(new_n506_), .A3(new_n508_), .A4(new_n512_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n482_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n399_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G231gat), .A2(G233gat), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n447_), .B(new_n520_), .Z(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT77), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(new_n494_), .ZN(new_n523_));
  XOR2_X1   g322(.A(G127gat), .B(G155gat), .Z(new_n524_));
  XNOR2_X1  g323(.A(G183gat), .B(G211gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT17), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n528_), .A2(KEYINPUT17), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n523_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n531_), .A2(KEYINPUT79), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n531_), .B(KEYINPUT79), .C1(new_n529_), .C2(new_n523_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n440_), .A2(new_n485_), .ZN(new_n536_));
  XOR2_X1   g335(.A(KEYINPUT69), .B(KEYINPUT34), .Z(new_n537_));
  NAND2_X1  g336(.A1(G232gat), .A2(G233gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n539_), .A2(KEYINPUT35), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT72), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n536_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n539_), .A2(KEYINPUT35), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n543_), .B(KEYINPUT73), .Z(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n487_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT70), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NOR3_X1   g347(.A1(new_n456_), .A2(new_n457_), .A3(KEYINPUT67), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n459_), .B1(new_n435_), .B2(new_n438_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n462_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n464_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n461_), .A2(KEYINPUT68), .A3(new_n462_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n554_), .A2(KEYINPUT70), .A3(new_n487_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n545_), .B1(new_n548_), .B2(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(KEYINPUT70), .B1(new_n554_), .B2(new_n487_), .ZN(new_n557_));
  AOI211_X1 g356(.A(new_n547_), .B(new_n486_), .C1(new_n552_), .C2(new_n553_), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT71), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT71), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n548_), .A2(new_n555_), .A3(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n559_), .A2(new_n542_), .A3(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n543_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n556_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G190gat), .B(G218gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G134gat), .B(G162gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n567_), .B(KEYINPUT36), .Z(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n564_), .A2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n567_), .A2(KEYINPUT36), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  AOI211_X1 g371(.A(new_n556_), .B(new_n572_), .C1(new_n562_), .C2(new_n563_), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT37), .B1(new_n570_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(KEYINPUT74), .ZN(new_n575_));
  INV_X1    g374(.A(new_n542_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n548_), .A2(new_n555_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n576_), .B1(new_n577_), .B2(KEYINPUT71), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n543_), .B1(new_n578_), .B2(new_n561_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n568_), .B1(new_n579_), .B2(new_n556_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n564_), .A2(new_n571_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT74), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(new_n583_), .A3(KEYINPUT37), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n562_), .A2(new_n563_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n556_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n569_), .B1(new_n587_), .B2(KEYINPUT75), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT75), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n585_), .A2(new_n589_), .A3(new_n586_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n573_), .B1(new_n588_), .B2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT76), .B(KEYINPUT37), .ZN(new_n592_));
  AOI22_X1  g391(.A1(new_n575_), .A2(new_n584_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n519_), .A2(new_n535_), .A3(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n369_), .B(KEYINPUT102), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n594_), .A2(new_n489_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT38), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n568_), .B1(new_n564_), .B2(new_n589_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n579_), .A2(KEYINPUT75), .A3(new_n556_), .ZN(new_n600_));
  OAI211_X1 g399(.A(KEYINPUT103), .B(new_n581_), .C1(new_n599_), .C2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(KEYINPUT75), .B1(new_n579_), .B2(new_n556_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(new_n568_), .A3(new_n590_), .ZN(new_n604_));
  AOI21_X1  g403(.A(KEYINPUT103), .B1(new_n604_), .B2(new_n581_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n519_), .A2(new_n535_), .A3(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n489_), .B1(new_n608_), .B2(new_n369_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n598_), .A2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n610_), .B1(new_n597_), .B2(new_n596_), .ZN(G1324gat));
  NAND3_X1  g410(.A1(new_n594_), .A2(new_n490_), .A3(new_n393_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n607_), .A2(new_n535_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n399_), .A2(new_n613_), .A3(new_n518_), .A4(new_n393_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT104), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n615_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT39), .ZN(new_n619_));
  OAI21_X1  g418(.A(G8gat), .B1(new_n619_), .B2(KEYINPUT105), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n618_), .A2(new_n621_), .B1(KEYINPUT105), .B2(new_n619_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n619_), .A2(KEYINPUT105), .ZN(new_n623_));
  AOI211_X1 g422(.A(new_n623_), .B(new_n620_), .C1(new_n616_), .C2(new_n617_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n612_), .B1(new_n622_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT40), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  OAI211_X1 g426(.A(KEYINPUT40), .B(new_n612_), .C1(new_n622_), .C2(new_n624_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(G1325gat));
  INV_X1    g428(.A(new_n243_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n230_), .B1(new_n608_), .B2(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT41), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n594_), .A2(new_n230_), .A3(new_n630_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(G1326gat));
  INV_X1    g433(.A(G22gat), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n608_), .B2(new_n301_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT42), .Z(new_n637_));
  NAND3_X1  g436(.A1(new_n594_), .A2(new_n635_), .A3(new_n301_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(G1327gat));
  NOR3_X1   g438(.A1(new_n519_), .A2(new_n534_), .A3(new_n606_), .ZN(new_n640_));
  INV_X1    g439(.A(G29gat), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(new_n641_), .A3(new_n369_), .ZN(new_n642_));
  XOR2_X1   g441(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n369_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n645_), .A2(new_n301_), .A3(new_n389_), .A4(new_n392_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n364_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n361_), .A2(new_n362_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  AOI22_X1  g448(.A1(new_n649_), .A2(new_n365_), .B1(new_n369_), .B2(new_n381_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n646_), .B1(new_n650_), .B2(new_n301_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n397_), .B1(new_n651_), .B2(new_n243_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n604_), .A2(new_n581_), .A3(new_n592_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n583_), .B1(new_n582_), .B2(KEYINPUT37), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT37), .ZN(new_n655_));
  AOI211_X1 g454(.A(KEYINPUT74), .B(new_n655_), .C1(new_n580_), .C2(new_n581_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n653_), .B1(new_n654_), .B2(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n644_), .B1(new_n652_), .B2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n399_), .A2(new_n593_), .A3(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n535_), .A2(new_n518_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(KEYINPUT44), .B1(new_n661_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n661_), .A2(KEYINPUT44), .A3(new_n663_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n665_), .A2(new_n595_), .A3(new_n666_), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n667_), .A2(KEYINPUT107), .A3(G29gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(KEYINPUT107), .B1(new_n667_), .B2(G29gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n642_), .B1(new_n668_), .B2(new_n669_), .ZN(G1328gat));
  INV_X1    g469(.A(KEYINPUT46), .ZN(new_n671_));
  INV_X1    g470(.A(G36gat), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673_));
  AOI211_X1 g472(.A(new_n673_), .B(new_n662_), .C1(new_n658_), .C2(new_n660_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n664_), .A2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n672_), .B1(new_n675_), .B2(new_n393_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n640_), .A2(new_n672_), .A3(new_n393_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT45), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n677_), .B(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n671_), .B1(new_n676_), .B2(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n677_), .B(KEYINPUT45), .ZN(new_n681_));
  INV_X1    g480(.A(new_n393_), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n664_), .A2(new_n674_), .A3(new_n682_), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n681_), .B(KEYINPUT46), .C1(new_n672_), .C2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n680_), .A2(new_n684_), .ZN(G1329gat));
  NAND2_X1  g484(.A1(new_n640_), .A2(new_n630_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(new_n235_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n665_), .A2(new_n666_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n243_), .A2(new_n235_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n687_), .B1(new_n688_), .B2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(KEYINPUT47), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT47), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n693_), .B(new_n687_), .C1(new_n688_), .C2(new_n690_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(G1330gat));
  INV_X1    g494(.A(G50gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n640_), .A2(new_n696_), .A3(new_n301_), .ZN(new_n697_));
  AOI211_X1 g496(.A(KEYINPUT108), .B(new_n696_), .C1(new_n675_), .C2(new_n301_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT108), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n665_), .A2(new_n301_), .A3(new_n666_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n700_), .B2(G50gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n697_), .B1(new_n698_), .B2(new_n701_), .ZN(G1331gat));
  INV_X1    g501(.A(new_n595_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n652_), .A2(new_n516_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n593_), .A2(new_n535_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(new_n482_), .A3(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT109), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n703_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n708_), .B1(new_n707_), .B2(new_n706_), .ZN(new_n709_));
  INV_X1    g508(.A(G57gat), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n709_), .A2(KEYINPUT110), .A3(new_n710_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n482_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n534_), .A2(new_n517_), .ZN(new_n716_));
  NOR4_X1   g515(.A1(new_n652_), .A2(new_n715_), .A3(new_n607_), .A4(new_n716_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n645_), .A2(new_n710_), .ZN(new_n718_));
  AOI22_X1  g517(.A1(new_n713_), .A2(new_n714_), .B1(new_n717_), .B2(new_n718_), .ZN(G1332gat));
  INV_X1    g518(.A(G64gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n720_), .B1(new_n717_), .B2(new_n393_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT48), .Z(new_n722_));
  INV_X1    g521(.A(new_n706_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n723_), .A2(new_n720_), .A3(new_n393_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(G1333gat));
  INV_X1    g524(.A(G71gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n726_), .B1(new_n717_), .B2(new_n630_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT49), .Z(new_n728_));
  NAND3_X1  g527(.A1(new_n723_), .A2(new_n726_), .A3(new_n630_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1334gat));
  INV_X1    g529(.A(G78gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n717_), .B2(new_n301_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT50), .Z(new_n733_));
  NAND3_X1  g532(.A1(new_n723_), .A2(new_n731_), .A3(new_n301_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1335gat));
  NOR2_X1   g534(.A1(new_n715_), .A2(new_n534_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n704_), .A2(new_n607_), .A3(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(new_n400_), .A3(new_n595_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n517_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n658_), .B2(new_n660_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n740_), .A2(new_n369_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n738_), .B1(new_n741_), .B2(new_n400_), .ZN(G1336gat));
  AOI21_X1  g541(.A(new_n401_), .B1(new_n740_), .B2(new_n393_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n682_), .A2(G92gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n737_), .B2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n745_), .B(new_n746_), .ZN(G1337gat));
  AOI21_X1  g546(.A(new_n430_), .B1(new_n740_), .B2(new_n630_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n243_), .A2(new_n422_), .A3(new_n421_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n737_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n750_), .B(new_n751_), .ZN(G1338gat));
  NAND3_X1  g551(.A1(new_n737_), .A2(new_n415_), .A3(new_n301_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n740_), .A2(new_n301_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n755_), .B2(G106gat), .ZN(new_n756_));
  AOI211_X1 g555(.A(KEYINPUT52), .B(new_n415_), .C1(new_n740_), .C2(new_n301_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT53), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT53), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n760_), .B(new_n753_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1339gat));
  INV_X1    g561(.A(KEYINPUT115), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n581_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT103), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n453_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n469_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n466_), .A2(new_n468_), .A3(KEYINPUT55), .A4(new_n453_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT56), .B1(new_n771_), .B2(new_n474_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT56), .ZN(new_n773_));
  AOI211_X1 g572(.A(new_n773_), .B(new_n476_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n516_), .B(new_n477_), .C1(new_n772_), .C2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n512_), .B1(new_n507_), .B2(new_n503_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n776_), .B1(new_n503_), .B2(new_n501_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n515_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n478_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n775_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT57), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT113), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n766_), .A2(new_n601_), .A3(new_n780_), .A4(new_n782_), .ZN(new_n783_));
  OR3_X1    g582(.A1(new_n772_), .A2(new_n774_), .A3(KEYINPUT114), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n772_), .A2(KEYINPUT114), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n778_), .A2(new_n477_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n784_), .A2(KEYINPUT58), .A3(new_n785_), .A4(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT58), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n785_), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n772_), .A2(new_n774_), .A3(KEYINPUT114), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n788_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n787_), .A2(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n783_), .B1(new_n657_), .B2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n782_), .B1(new_n606_), .B2(new_n780_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n535_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n715_), .A2(new_n534_), .A3(new_n517_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n575_), .A2(new_n584_), .ZN(new_n798_));
  AOI211_X1 g597(.A(new_n796_), .B(new_n797_), .C1(new_n798_), .C2(new_n653_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n796_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n797_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n657_), .B2(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n799_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n795_), .A2(new_n803_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n393_), .A2(new_n301_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n595_), .A2(new_n630_), .A3(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n763_), .B1(new_n804_), .B2(new_n807_), .ZN(new_n808_));
  AOI211_X1 g607(.A(KEYINPUT115), .B(new_n806_), .C1(new_n795_), .C2(new_n803_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(G113gat), .B1(new_n810_), .B2(new_n516_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT59), .B1(new_n804_), .B2(new_n807_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT59), .ZN(new_n814_));
  AOI211_X1 g613(.A(new_n814_), .B(new_n806_), .C1(new_n795_), .C2(new_n803_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n812_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n796_), .B1(new_n593_), .B2(new_n797_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n657_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n766_), .A2(new_n601_), .A3(new_n780_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n820_), .A2(KEYINPUT113), .A3(new_n781_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n798_), .A2(new_n653_), .A3(new_n791_), .A4(new_n787_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n821_), .A2(new_n822_), .A3(new_n783_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n819_), .B1(new_n535_), .B2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n814_), .B1(new_n824_), .B2(new_n806_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n804_), .A2(KEYINPUT59), .A3(new_n807_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(KEYINPUT116), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n816_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(G113gat), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n829_), .B1(new_n516_), .B2(KEYINPUT117), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n830_), .B1(KEYINPUT117), .B2(new_n829_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n811_), .B1(new_n828_), .B2(new_n831_), .ZN(G1340gat));
  AOI21_X1  g631(.A(new_n715_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n833_));
  INV_X1    g632(.A(G120gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT115), .B1(new_n824_), .B2(new_n806_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n804_), .A2(new_n763_), .A3(new_n807_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n834_), .B1(new_n715_), .B2(KEYINPUT60), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(KEYINPUT60), .B2(new_n834_), .ZN(new_n839_));
  OAI22_X1  g638(.A1(new_n833_), .A2(new_n834_), .B1(new_n837_), .B2(new_n839_), .ZN(G1341gat));
  INV_X1    g639(.A(G127gat), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n535_), .A2(new_n841_), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n813_), .A2(new_n815_), .A3(new_n812_), .ZN(new_n843_));
  AOI21_X1  g642(.A(KEYINPUT116), .B1(new_n825_), .B2(new_n826_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n842_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n841_), .B1(new_n837_), .B2(new_n535_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(KEYINPUT118), .A3(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n848_));
  INV_X1    g647(.A(new_n842_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n849_), .B1(new_n816_), .B2(new_n827_), .ZN(new_n850_));
  AOI21_X1  g649(.A(G127gat), .B1(new_n810_), .B2(new_n534_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n848_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n847_), .A2(new_n852_), .ZN(G1342gat));
  INV_X1    g652(.A(G134gat), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n837_), .B2(new_n606_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  OAI211_X1 g656(.A(KEYINPUT119), .B(new_n854_), .C1(new_n837_), .C2(new_n606_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n593_), .A2(G134gat), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  AOI22_X1  g659(.A1(new_n857_), .A2(new_n858_), .B1(new_n828_), .B2(new_n860_), .ZN(G1343gat));
  NOR2_X1   g660(.A1(new_n824_), .A2(new_n630_), .ZN(new_n862_));
  NOR3_X1   g661(.A1(new_n703_), .A2(new_n394_), .A3(new_n393_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(KEYINPUT121), .B1(new_n864_), .B2(new_n517_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n862_), .A2(new_n866_), .A3(new_n516_), .A4(new_n863_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT120), .B(G141gat), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n865_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1344gat));
  NOR2_X1   g670(.A1(new_n864_), .A2(new_n715_), .ZN(new_n872_));
  XOR2_X1   g671(.A(new_n872_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g672(.A1(new_n864_), .A2(new_n535_), .ZN(new_n874_));
  XOR2_X1   g673(.A(KEYINPUT61), .B(G155gat), .Z(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1346gat));
  OAI21_X1  g675(.A(G162gat), .B1(new_n864_), .B2(new_n657_), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n606_), .A2(G162gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n864_), .B2(new_n878_), .ZN(G1347gat));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n301_), .B1(new_n795_), .B2(new_n803_), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n595_), .A2(new_n243_), .A3(new_n682_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n516_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n880_), .B1(new_n885_), .B2(G169gat), .ZN(new_n886_));
  AOI211_X1 g685(.A(KEYINPUT62), .B(new_n215_), .C1(new_n884_), .C2(new_n516_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n883_), .A2(KEYINPUT122), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n889_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n888_), .A2(new_n890_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT22), .B(G169gat), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n516_), .A2(new_n892_), .ZN(new_n893_));
  OAI22_X1  g692(.A1(new_n886_), .A2(new_n887_), .B1(new_n891_), .B2(new_n893_), .ZN(G1348gat));
  OAI21_X1  g693(.A(new_n216_), .B1(new_n891_), .B2(new_n715_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n881_), .B(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n715_), .A2(new_n216_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n897_), .A2(new_n882_), .A3(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(KEYINPUT124), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT124), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n897_), .A2(new_n901_), .A3(new_n882_), .A4(new_n898_), .ZN(new_n902_));
  AND3_X1   g701(.A1(new_n895_), .A2(new_n900_), .A3(new_n902_), .ZN(G1349gat));
  NAND3_X1  g702(.A1(new_n897_), .A2(new_n534_), .A3(new_n882_), .ZN(new_n904_));
  INV_X1    g703(.A(G183gat), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n535_), .A2(new_n337_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n907_), .B1(new_n888_), .B2(new_n890_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT125), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  OAI211_X1 g709(.A(KEYINPUT125), .B(new_n907_), .C1(new_n888_), .C2(new_n890_), .ZN(new_n911_));
  AND3_X1   g710(.A1(new_n906_), .A2(new_n910_), .A3(new_n911_), .ZN(G1350gat));
  OAI21_X1  g711(.A(G190gat), .B1(new_n891_), .B2(new_n657_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n607_), .A2(new_n211_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n891_), .B2(new_n914_), .ZN(G1351gat));
  NOR3_X1   g714(.A1(new_n682_), .A2(new_n394_), .A3(new_n369_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n862_), .A2(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n917_), .A2(new_n517_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(new_n272_), .ZN(G1352gat));
  NOR2_X1   g718(.A1(new_n917_), .A2(new_n715_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(G204gat), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n921_), .B1(new_n271_), .B2(new_n920_), .ZN(G1353gat));
  AOI21_X1  g721(.A(new_n535_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n923_));
  INV_X1    g722(.A(new_n923_), .ZN(new_n924_));
  OAI21_X1  g723(.A(KEYINPUT126), .B1(new_n917_), .B2(new_n924_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n927_));
  NAND4_X1  g726(.A1(new_n862_), .A2(new_n927_), .A3(new_n916_), .A4(new_n923_), .ZN(new_n928_));
  AND3_X1   g727(.A1(new_n925_), .A2(new_n926_), .A3(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n926_), .B1(new_n925_), .B2(new_n928_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n929_), .A2(new_n930_), .ZN(G1354gat));
  OAI21_X1  g730(.A(G218gat), .B1(new_n917_), .B2(new_n657_), .ZN(new_n932_));
  OR2_X1    g731(.A1(new_n606_), .A2(G218gat), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n917_), .B2(new_n933_), .ZN(G1355gat));
endmodule


