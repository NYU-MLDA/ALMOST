//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n622_, new_n623_,
    new_n624_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n785_, new_n787_, new_n788_, new_n789_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n802_, new_n803_, new_n804_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n841_, new_n843_, new_n844_, new_n845_,
    new_n847_, new_n848_, new_n849_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT34), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT35), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT72), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G92gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT9), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(KEYINPUT65), .A3(G85gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n207_), .B1(new_n209_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n207_), .A2(G85gat), .ZN(new_n213_));
  INV_X1    g012(.A(G85gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(G92gat), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n210_), .B1(new_n213_), .B2(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT66), .B1(new_n212_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n218_), .A2(KEYINPUT9), .ZN(new_n219_));
  OAI21_X1  g018(.A(G92gat), .B1(new_n219_), .B2(new_n208_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n214_), .A2(G92gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n207_), .A2(G85gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT9), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n220_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G99gat), .A2(G106gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT6), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  XOR2_X1   g029(.A(KEYINPUT10), .B(G99gat), .Z(new_n231_));
  INV_X1    g030(.A(G106gat), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n230_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n217_), .A2(new_n225_), .A3(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT7), .ZN(new_n235_));
  INV_X1    g034(.A(G99gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n236_), .A3(new_n232_), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n237_), .A2(new_n228_), .A3(new_n229_), .A4(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n213_), .A2(new_n215_), .ZN(new_n240_));
  AOI21_X1  g039(.A(KEYINPUT67), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT8), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n239_), .A2(KEYINPUT67), .A3(new_n240_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT8), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n234_), .B(new_n243_), .C1(new_n241_), .C2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G29gat), .B(G36gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G43gat), .B(G50gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT15), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n246_), .A2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT73), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n203_), .A2(KEYINPUT35), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n239_), .A2(new_n240_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(KEYINPUT8), .A3(new_n244_), .ZN(new_n257_));
  AND3_X1   g056(.A1(new_n257_), .A2(new_n243_), .A3(new_n234_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n253_), .B1(new_n258_), .B2(new_n249_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT74), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n252_), .A2(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n259_), .A2(new_n260_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n206_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n251_), .A2(KEYINPUT73), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n251_), .A2(KEYINPUT73), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n259_), .B(new_n205_), .C1(new_n265_), .C2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT76), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n252_), .A2(KEYINPUT76), .A3(new_n205_), .A4(new_n259_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n264_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G190gat), .B(G218gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(G162gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT75), .B(G134gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n273_), .B(new_n274_), .Z(new_n275_));
  INV_X1    g074(.A(KEYINPUT36), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  OR2_X1    g076(.A1(new_n275_), .A2(new_n276_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n271_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n269_), .A2(new_n270_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n280_), .A2(new_n276_), .A3(new_n275_), .A4(new_n264_), .ZN(new_n281_));
  AND3_X1   g080(.A1(new_n279_), .A2(KEYINPUT37), .A3(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT37), .B1(new_n279_), .B2(new_n281_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(G15gat), .B(G22gat), .Z(new_n285_));
  XOR2_X1   g084(.A(KEYINPUT77), .B(G1gat), .Z(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(G8gat), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n285_), .B1(new_n287_), .B2(KEYINPUT14), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G1gat), .B(G8gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G231gat), .A2(G233gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(G57gat), .ZN(new_n293_));
  INV_X1    g092(.A(G64gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT11), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G57gat), .A2(G64gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n295_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT68), .ZN(new_n299_));
  INV_X1    g098(.A(G71gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(G78gat), .ZN(new_n301_));
  INV_X1    g100(.A(G78gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(G71gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  AND3_X1   g103(.A1(new_n298_), .A2(new_n299_), .A3(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n299_), .B1(new_n298_), .B2(new_n304_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n296_), .B1(new_n295_), .B2(new_n297_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NOR3_X1   g107(.A1(new_n305_), .A2(new_n306_), .A3(new_n308_), .ZN(new_n309_));
  AND2_X1   g108(.A1(G57gat), .A2(G64gat), .ZN(new_n310_));
  NOR2_X1   g109(.A1(G57gat), .A2(G64gat), .ZN(new_n311_));
  NOR3_X1   g110(.A1(new_n310_), .A2(new_n311_), .A3(KEYINPUT11), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G71gat), .B(G78gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT68), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n298_), .A2(new_n299_), .A3(new_n304_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n307_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n309_), .A2(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n292_), .B(new_n317_), .Z(new_n318_));
  XNOR2_X1  g117(.A(G183gat), .B(G211gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G127gat), .B(G155gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  XOR2_X1   g122(.A(KEYINPUT79), .B(KEYINPUT17), .Z(new_n324_));
  NAND3_X1  g123(.A1(new_n318_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT69), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(new_n309_), .B2(new_n316_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n308_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n314_), .A2(new_n307_), .A3(new_n315_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n328_), .A2(KEYINPUT69), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n327_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n292_), .B(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n323_), .B(KEYINPUT17), .Z(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n325_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n284_), .A2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT80), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G155gat), .A2(G162gat), .ZN(new_n338_));
  OR2_X1    g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339_));
  NOR2_X1   g138(.A1(G141gat), .A2(G148gat), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT3), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G141gat), .A2(G148gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT2), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n338_), .B(new_n339_), .C1(new_n342_), .C2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n338_), .A2(KEYINPUT1), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT89), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n338_), .A2(KEYINPUT1), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT89), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n338_), .A2(new_n350_), .A3(KEYINPUT1), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n348_), .A2(new_n349_), .A3(new_n351_), .A4(new_n339_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(new_n343_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n346_), .B1(new_n353_), .B2(new_n340_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n354_), .A2(KEYINPUT29), .ZN(new_n355_));
  INV_X1    g154(.A(G50gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT28), .B(G22gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G211gat), .B(G218gat), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT92), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G197gat), .B(G204gat), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT91), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n362_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT21), .ZN(new_n367_));
  INV_X1    g166(.A(new_n362_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(new_n363_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT93), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n354_), .A2(KEYINPUT29), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n367_), .A2(KEYINPUT93), .A3(new_n369_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n372_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(G233gat), .ZN(new_n376_));
  NOR2_X1   g175(.A1(KEYINPUT90), .A2(G228gat), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(KEYINPUT90), .A2(G228gat), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n376_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n370_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n380_), .B1(new_n354_), .B2(KEYINPUT29), .ZN(new_n382_));
  AOI22_X1  g181(.A1(new_n375_), .A2(new_n380_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(G78gat), .B(G106gat), .Z(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n383_), .A2(new_n384_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n359_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n387_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n359_), .A2(KEYINPUT94), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(new_n385_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n386_), .A2(KEYINPUT94), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n388_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(G169gat), .A2(G176gat), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT82), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G169gat), .A2(G176gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT83), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(KEYINPUT24), .A3(new_n399_), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n400_), .A2(KEYINPUT84), .ZN(new_n401_));
  XOR2_X1   g200(.A(KEYINPUT26), .B(G190gat), .Z(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT25), .B(G183gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n400_), .A2(KEYINPUT84), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n397_), .A2(KEYINPUT24), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G183gat), .A2(G190gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT23), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT23), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n410_), .A2(G183gat), .A3(G190gat), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n407_), .A2(new_n412_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n401_), .A2(new_n405_), .A3(new_n406_), .A4(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n409_), .A2(KEYINPUT86), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n415_), .B1(new_n412_), .B2(KEYINPUT86), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n416_), .B1(G183gat), .B2(G190gat), .ZN(new_n417_));
  INV_X1    g216(.A(G169gat), .ZN(new_n418_));
  OR3_X1    g217(.A1(new_n418_), .A2(KEYINPUT85), .A3(KEYINPUT22), .ZN(new_n419_));
  INV_X1    g218(.A(G176gat), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT22), .B1(new_n418_), .B2(KEYINPUT85), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n419_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n417_), .A2(new_n399_), .A3(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n414_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT30), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT87), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G227gat), .A2(G233gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(new_n300_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(new_n236_), .ZN(new_n430_));
  XOR2_X1   g229(.A(G15gat), .B(G43gat), .Z(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n427_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT88), .B(KEYINPUT31), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n434_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n427_), .A2(new_n436_), .A3(new_n432_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n426_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT87), .ZN(new_n440_));
  XOR2_X1   g239(.A(G113gat), .B(G120gat), .Z(new_n441_));
  XNOR2_X1  g240(.A(G127gat), .B(G134gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n439_), .A2(new_n440_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n443_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n445_), .B1(new_n426_), .B2(KEYINPUT87), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n438_), .A2(new_n447_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n435_), .A2(new_n444_), .A3(new_n446_), .A4(new_n437_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n394_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n393_), .A2(new_n450_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G226gat), .A2(G233gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT19), .ZN(new_n456_));
  INV_X1    g255(.A(new_n395_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n416_), .B1(KEYINPUT24), .B2(new_n457_), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n397_), .A2(KEYINPUT24), .A3(new_n398_), .ZN(new_n459_));
  OR2_X1    g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT95), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n404_), .B(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n462_), .A2(new_n402_), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT96), .B1(new_n460_), .B2(new_n463_), .ZN(new_n464_));
  NOR3_X1   g263(.A1(new_n463_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT96), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n412_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n468_), .B1(G183gat), .B2(G190gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT22), .B(G169gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n420_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n469_), .A2(new_n399_), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT97), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n472_), .A2(KEYINPUT97), .ZN(new_n474_));
  AOI22_X1  g273(.A1(new_n464_), .A2(new_n467_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n456_), .B1(new_n475_), .B2(new_n370_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n381_), .A2(new_n424_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n476_), .A2(KEYINPUT20), .A3(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G8gat), .B(G36gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(G92gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT18), .B(G64gat), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n480_), .B(new_n481_), .Z(new_n482_));
  NAND3_X1  g281(.A1(new_n370_), .A2(new_n423_), .A3(new_n414_), .ZN(new_n483_));
  OAI211_X1 g282(.A(KEYINPUT20), .B(new_n483_), .C1(new_n475_), .C2(new_n370_), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n484_), .A2(KEYINPUT98), .A3(new_n456_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT98), .B1(new_n484_), .B2(new_n456_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n478_), .B(new_n482_), .C1(new_n485_), .C2(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n484_), .A2(new_n456_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n472_), .ZN(new_n489_));
  AOI211_X1 g288(.A(new_n465_), .B(new_n489_), .C1(new_n372_), .C2(new_n374_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT20), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT102), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT102), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n372_), .A2(new_n374_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(new_n472_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n493_), .B(KEYINPUT20), .C1(new_n495_), .C2(new_n465_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n492_), .A2(new_n496_), .A3(new_n477_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n488_), .B1(new_n497_), .B2(new_n456_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n482_), .B(KEYINPUT103), .ZN(new_n499_));
  OAI211_X1 g298(.A(KEYINPUT27), .B(new_n487_), .C1(new_n498_), .C2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT27), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n484_), .A2(new_n456_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT98), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n484_), .A2(KEYINPUT98), .A3(new_n456_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n482_), .B1(new_n506_), .B2(new_n478_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n487_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n501_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n500_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n354_), .A2(new_n443_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT99), .B1(new_n354_), .B2(new_n443_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G225gat), .A2(G233gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  OR2_X1    g316(.A1(new_n517_), .A2(KEYINPUT101), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(KEYINPUT101), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n512_), .A2(KEYINPUT4), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n520_), .B1(new_n515_), .B2(KEYINPUT4), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n516_), .B(KEYINPUT100), .Z(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n518_), .A2(new_n519_), .A3(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G1gat), .B(G29gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(new_n214_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT0), .B(G57gat), .ZN(new_n527_));
  XOR2_X1   g326(.A(new_n526_), .B(new_n527_), .Z(new_n528_));
  NAND2_X1  g327(.A1(new_n524_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n528_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n518_), .A2(new_n523_), .A3(new_n530_), .A4(new_n519_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n454_), .A2(new_n511_), .A3(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n507_), .A2(new_n508_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n521_), .A2(new_n516_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n515_), .A2(new_n522_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n536_), .A2(new_n528_), .A3(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n531_), .B(KEYINPUT33), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n535_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n482_), .A2(KEYINPUT32), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n506_), .A2(new_n478_), .A3(new_n541_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n532_), .B(new_n542_), .C1(new_n498_), .C2(new_n541_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n544_), .A2(new_n451_), .A3(new_n393_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n337_), .B1(new_n534_), .B2(new_n545_), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n246_), .A2(KEYINPUT12), .A3(new_n317_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT12), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n328_), .A2(KEYINPUT69), .A3(new_n329_), .ZN(new_n549_));
  AOI21_X1  g348(.A(KEYINPUT69), .B1(new_n328_), .B2(new_n329_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n246_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n547_), .B1(new_n548_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G230gat), .A2(G233gat), .ZN(new_n553_));
  XOR2_X1   g352(.A(new_n553_), .B(KEYINPUT64), .Z(new_n554_));
  OAI21_X1  g353(.A(new_n554_), .B1(new_n331_), .B2(new_n246_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n552_), .A2(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n245_), .A2(new_n241_), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n217_), .A2(new_n225_), .A3(new_n233_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  AOI22_X1  g359(.A1(new_n560_), .A2(new_n243_), .B1(new_n327_), .B2(new_n330_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT70), .B1(new_n331_), .B2(new_n246_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT70), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n258_), .A2(new_n563_), .A3(new_n330_), .A4(new_n327_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n561_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n557_), .B1(new_n565_), .B2(new_n554_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT71), .B(G204gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT5), .B(G176gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G120gat), .B(G148gat), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n569_), .B(new_n570_), .Z(new_n571_));
  NAND2_X1  g370(.A1(new_n566_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n571_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n557_), .B(new_n573_), .C1(new_n554_), .C2(new_n565_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT13), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n290_), .B(new_n249_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G229gat), .A2(G233gat), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n249_), .B(KEYINPUT15), .Z(new_n582_));
  OR2_X1    g381(.A1(new_n582_), .A2(new_n290_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n290_), .A2(new_n249_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n583_), .A2(new_n584_), .A3(new_n579_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n581_), .A2(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(G113gat), .B(G141gat), .Z(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(G197gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(KEYINPUT81), .B(G169gat), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n588_), .B(new_n589_), .Z(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n586_), .A2(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n581_), .A2(new_n585_), .A3(new_n590_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n577_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n546_), .A2(new_n596_), .ZN(new_n597_));
  NOR3_X1   g396(.A1(new_n597_), .A2(new_n533_), .A3(new_n286_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n598_), .A2(KEYINPUT38), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(KEYINPUT38), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n279_), .A2(new_n281_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT104), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n279_), .A2(KEYINPUT104), .A3(new_n281_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n606_), .B1(new_n534_), .B2(new_n545_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n607_), .A2(new_n335_), .A3(new_n596_), .ZN(new_n608_));
  OAI21_X1  g407(.A(G1gat), .B1(new_n608_), .B2(new_n533_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n599_), .A2(new_n600_), .A3(new_n609_), .ZN(G1324gat));
  NOR2_X1   g409(.A1(new_n511_), .A2(G8gat), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n546_), .A2(new_n596_), .A3(new_n611_), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n608_), .A2(new_n511_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(G8gat), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n614_), .A2(KEYINPUT39), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(KEYINPUT39), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n612_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT40), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  OAI211_X1 g418(.A(KEYINPUT40), .B(new_n612_), .C1(new_n615_), .C2(new_n616_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(G1325gat));
  OAI21_X1  g420(.A(G15gat), .B1(new_n608_), .B2(new_n451_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT41), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n597_), .A2(G15gat), .A3(new_n451_), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1326gat));
  OR3_X1    g424(.A1(new_n597_), .A2(G22gat), .A3(new_n393_), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n608_), .A2(new_n393_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n627_), .A2(G22gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n628_), .A2(new_n629_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n626_), .B1(new_n630_), .B2(new_n631_), .ZN(G1327gat));
  AOI21_X1  g431(.A(new_n605_), .B1(new_n534_), .B2(new_n545_), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n577_), .A2(new_n335_), .A3(new_n595_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(G29gat), .B1(new_n636_), .B2(new_n532_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n284_), .B1(new_n534_), .B2(new_n545_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT43), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  AOI211_X1 g439(.A(KEYINPUT43), .B(new_n284_), .C1(new_n534_), .C2(new_n545_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n634_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT44), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  OAI211_X1 g443(.A(KEYINPUT44), .B(new_n634_), .C1(new_n640_), .C2(new_n641_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n532_), .A2(G29gat), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n637_), .B1(new_n646_), .B2(new_n647_), .ZN(G1328gat));
  NAND3_X1  g447(.A1(new_n644_), .A2(new_n510_), .A3(new_n645_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(G36gat), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT106), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n500_), .A2(new_n509_), .A3(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n651_), .B1(new_n500_), .B2(new_n509_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n635_), .A2(G36gat), .A3(new_n656_), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n657_), .B(KEYINPUT45), .Z(new_n658_));
  NAND2_X1  g457(.A1(new_n650_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT46), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n650_), .A2(new_n658_), .A3(KEYINPUT46), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1329gat));
  NAND4_X1  g462(.A1(new_n644_), .A2(G43gat), .A3(new_n450_), .A4(new_n645_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n635_), .A2(new_n451_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n664_), .B1(G43gat), .B2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g466(.A1(new_n644_), .A2(new_n394_), .A3(new_n645_), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n668_), .A2(KEYINPUT107), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(KEYINPUT107), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(G50gat), .A3(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n636_), .A2(new_n356_), .A3(new_n394_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1331gat));
  NOR2_X1   g472(.A1(new_n576_), .A2(new_n594_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n607_), .A2(new_n335_), .A3(new_n674_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n675_), .A2(new_n293_), .A3(new_n533_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n546_), .A2(new_n674_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n293_), .B1(new_n677_), .B2(new_n533_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n679_), .A2(KEYINPUT108), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(KEYINPUT108), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n676_), .B1(new_n680_), .B2(new_n681_), .ZN(G1332gat));
  OR2_X1    g481(.A1(new_n675_), .A2(new_n656_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n683_), .A2(G64gat), .A3(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n683_), .B2(G64gat), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n655_), .A2(new_n294_), .ZN(new_n687_));
  OAI22_X1  g486(.A1(new_n685_), .A2(new_n686_), .B1(new_n677_), .B2(new_n687_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT110), .ZN(G1333gat));
  OAI21_X1  g488(.A(G71gat), .B1(new_n675_), .B2(new_n451_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT49), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n450_), .A2(new_n300_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT111), .Z(new_n693_));
  OAI21_X1  g492(.A(new_n691_), .B1(new_n677_), .B2(new_n693_), .ZN(G1334gat));
  OAI21_X1  g493(.A(G78gat), .B1(new_n675_), .B2(new_n393_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT50), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n394_), .A2(new_n302_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n696_), .B1(new_n677_), .B2(new_n697_), .ZN(G1335gat));
  NOR3_X1   g497(.A1(new_n576_), .A2(new_n335_), .A3(new_n594_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n633_), .A2(new_n699_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT112), .Z(new_n701_));
  AOI21_X1  g500(.A(G85gat), .B1(new_n701_), .B2(new_n532_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n699_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT113), .Z(new_n704_));
  OAI21_X1  g503(.A(new_n209_), .B1(new_n533_), .B2(new_n218_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n702_), .B1(new_n704_), .B2(new_n705_), .ZN(G1336gat));
  AOI21_X1  g505(.A(G92gat), .B1(new_n701_), .B2(new_n510_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n655_), .A2(G92gat), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT114), .Z(new_n709_));
  AOI21_X1  g508(.A(new_n707_), .B1(new_n704_), .B2(new_n709_), .ZN(G1337gat));
  NAND3_X1  g509(.A1(new_n701_), .A2(new_n231_), .A3(new_n450_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G99gat), .B1(new_n703_), .B2(new_n451_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n713_), .B(new_n715_), .ZN(G1338gat));
  NAND3_X1  g515(.A1(new_n701_), .A2(new_n232_), .A3(new_n394_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n394_), .B(new_n699_), .C1(new_n640_), .C2(new_n641_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT52), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n718_), .A2(new_n719_), .A3(G106gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n718_), .B2(G106gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g522(.A(G113gat), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n335_), .A2(new_n595_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT116), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n726_), .A2(new_n284_), .A3(new_n576_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT54), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n594_), .A2(new_n574_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT55), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n246_), .A2(new_n317_), .A3(KEYINPUT12), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n731_), .B1(new_n561_), .B2(KEYINPUT12), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n730_), .B1(new_n732_), .B2(new_n555_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n552_), .A2(KEYINPUT55), .A3(new_n556_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n562_), .A2(new_n564_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n554_), .B1(new_n552_), .B2(new_n736_), .ZN(new_n737_));
  OAI211_X1 g536(.A(KEYINPUT56), .B(new_n571_), .C1(new_n735_), .C2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  AOI221_X4 g538(.A(new_n547_), .B1(new_n551_), .B2(new_n548_), .C1(new_n562_), .C2(new_n564_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n733_), .B(new_n734_), .C1(new_n740_), .C2(new_n554_), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT56), .B1(new_n741_), .B2(new_n571_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n729_), .B1(new_n739_), .B2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT117), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n578_), .A2(new_n579_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n583_), .A2(new_n584_), .A3(new_n580_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n746_), .A2(new_n747_), .A3(new_n591_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n748_), .A2(new_n593_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n575_), .A2(new_n749_), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n729_), .B(KEYINPUT117), .C1(new_n739_), .C2(new_n742_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n745_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n752_), .A2(KEYINPUT57), .A3(new_n605_), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n574_), .B(new_n749_), .C1(new_n739_), .C2(new_n742_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT58), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n754_), .A2(KEYINPUT118), .A3(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n754_), .B2(KEYINPUT118), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n756_), .A2(new_n757_), .A3(new_n284_), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT57), .B1(new_n752_), .B2(new_n605_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n753_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n728_), .B1(new_n760_), .B2(new_n335_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT59), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n510_), .A2(new_n453_), .A3(new_n533_), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n761_), .A2(new_n762_), .A3(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n761_), .A2(KEYINPUT119), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT119), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n728_), .B(new_n766_), .C1(new_n760_), .C2(new_n335_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n765_), .A2(new_n767_), .A3(new_n763_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n764_), .B1(new_n768_), .B2(KEYINPUT59), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n724_), .B1(new_n769_), .B2(new_n594_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n768_), .A2(G113gat), .A3(new_n595_), .ZN(new_n771_));
  OAI21_X1  g570(.A(KEYINPUT120), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT120), .ZN(new_n773_));
  INV_X1    g572(.A(new_n771_), .ZN(new_n774_));
  AOI211_X1 g573(.A(new_n595_), .B(new_n764_), .C1(new_n768_), .C2(KEYINPUT59), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n773_), .B(new_n774_), .C1(new_n775_), .C2(new_n724_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n772_), .A2(new_n776_), .ZN(G1340gat));
  INV_X1    g576(.A(G120gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT60), .B1(new_n577_), .B2(new_n778_), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n768_), .A2(new_n779_), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n780_), .A2(new_n577_), .A3(new_n769_), .ZN(new_n781_));
  OAI22_X1  g580(.A1(new_n781_), .A2(new_n778_), .B1(KEYINPUT60), .B2(new_n780_), .ZN(G1341gat));
  INV_X1    g581(.A(new_n768_), .ZN(new_n783_));
  AOI21_X1  g582(.A(G127gat), .B1(new_n783_), .B2(new_n335_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n335_), .A2(G127gat), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n769_), .B2(new_n785_), .ZN(G1342gat));
  AOI21_X1  g585(.A(G134gat), .B1(new_n783_), .B2(new_n606_), .ZN(new_n787_));
  INV_X1    g586(.A(G134gat), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n284_), .A2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n787_), .B1(new_n769_), .B2(new_n789_), .ZN(G1343gat));
  NAND2_X1  g589(.A1(new_n765_), .A2(new_n767_), .ZN(new_n791_));
  NOR4_X1   g590(.A1(new_n791_), .A2(new_n533_), .A3(new_n452_), .A4(new_n655_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(new_n594_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n577_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(KEYINPUT121), .B(G148gat), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n795_), .B(new_n797_), .ZN(G1345gat));
  NAND2_X1  g597(.A1(new_n792_), .A2(new_n335_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(KEYINPUT61), .B(G155gat), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n799_), .B(new_n800_), .ZN(G1346gat));
  AOI21_X1  g600(.A(G162gat), .B1(new_n792_), .B2(new_n606_), .ZN(new_n802_));
  OAI21_X1  g601(.A(G162gat), .B1(new_n282_), .B2(new_n283_), .ZN(new_n803_));
  XOR2_X1   g602(.A(new_n803_), .B(KEYINPUT122), .Z(new_n804_));
  AOI21_X1  g603(.A(new_n802_), .B1(new_n792_), .B2(new_n804_), .ZN(G1347gat));
  INV_X1    g604(.A(KEYINPUT127), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n753_), .A2(new_n759_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n758_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n335_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n727_), .B(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n655_), .A2(KEYINPUT123), .A3(new_n533_), .A4(new_n450_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n510_), .A2(KEYINPUT106), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n814_), .A2(new_n533_), .A3(new_n450_), .A4(new_n652_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT123), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n813_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n812_), .A2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n806_), .B1(new_n820_), .B2(new_n393_), .ZN(new_n821_));
  NOR4_X1   g620(.A1(new_n812_), .A2(new_n819_), .A3(KEYINPUT127), .A4(new_n394_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n823_), .A2(new_n470_), .A3(new_n594_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n394_), .A2(new_n595_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n818_), .B(new_n825_), .C1(new_n809_), .C2(new_n811_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT124), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT124), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n761_), .A2(new_n828_), .A3(new_n818_), .A4(new_n825_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n827_), .A2(G169gat), .A3(new_n829_), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n830_), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT126), .B1(new_n830_), .B2(KEYINPUT62), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT62), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n827_), .A2(new_n834_), .A3(G169gat), .A4(new_n829_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT125), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n835_), .B(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n824_), .B1(new_n833_), .B2(new_n837_), .ZN(G1348gat));
  AOI21_X1  g637(.A(G176gat), .B1(new_n823_), .B2(new_n577_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n791_), .A2(new_n394_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n819_), .A2(new_n420_), .A3(new_n576_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n839_), .B1(new_n840_), .B2(new_n841_), .ZN(G1349gat));
  AND2_X1   g641(.A1(new_n335_), .A2(new_n462_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n840_), .A2(new_n335_), .A3(new_n818_), .ZN(new_n844_));
  INV_X1    g643(.A(G183gat), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n823_), .A2(new_n843_), .B1(new_n844_), .B2(new_n845_), .ZN(G1350gat));
  NAND3_X1  g645(.A1(new_n823_), .A2(new_n606_), .A3(new_n403_), .ZN(new_n847_));
  INV_X1    g646(.A(G190gat), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n821_), .A2(new_n822_), .A3(new_n284_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n847_), .B1(new_n848_), .B2(new_n849_), .ZN(G1351gat));
  INV_X1    g649(.A(new_n452_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n656_), .A2(new_n532_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n765_), .A2(new_n851_), .A3(new_n767_), .A4(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n594_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n577_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g657(.A(KEYINPUT63), .B(G211gat), .C1(new_n854_), .C2(new_n335_), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n854_), .A2(new_n335_), .ZN(new_n860_));
  XOR2_X1   g659(.A(KEYINPUT63), .B(G211gat), .Z(new_n861_));
  AOI21_X1  g660(.A(new_n859_), .B1(new_n860_), .B2(new_n861_), .ZN(G1354gat));
  INV_X1    g661(.A(G218gat), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n853_), .A2(new_n863_), .A3(new_n284_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n854_), .A2(new_n606_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n863_), .B2(new_n865_), .ZN(G1355gat));
endmodule


