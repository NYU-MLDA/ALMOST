//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 1 1 1 0 1 1 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n782_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n897_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n928_, new_n929_,
    new_n930_, new_n932_, new_n933_, new_n934_, new_n935_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n942_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_, new_n952_,
    new_n953_;
  OAI21_X1  g000(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(G169gat), .ZN(new_n204_));
  INV_X1    g003(.A(G176gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n203_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT23), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(G183gat), .A3(G190gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  OR3_X1    g010(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n206_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT82), .B(G190gat), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n214_), .B1(new_n215_), .B2(KEYINPUT26), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT25), .B(G183gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT83), .B1(new_n216_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT83), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT26), .ZN(new_n221_));
  OR2_X1    g020(.A1(KEYINPUT82), .A2(G190gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(KEYINPUT82), .A2(G190gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n221_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n220_), .B(new_n217_), .C1(new_n224_), .C2(new_n214_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n213_), .B1(new_n219_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT84), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n210_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n208_), .A2(new_n210_), .A3(new_n227_), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n228_), .B(new_n229_), .C1(G183gat), .C2(new_n215_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(new_n204_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n230_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n226_), .A2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G71gat), .B(G99gat), .ZN(new_n237_));
  INV_X1    g036(.A(G43gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n236_), .B(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(G127gat), .B(G134gat), .Z(new_n241_));
  XOR2_X1   g040(.A(G113gat), .B(G120gat), .Z(new_n242_));
  XOR2_X1   g041(.A(new_n241_), .B(new_n242_), .Z(new_n243_));
  XNOR2_X1  g042(.A(new_n240_), .B(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G227gat), .A2(G233gat), .ZN(new_n245_));
  XOR2_X1   g044(.A(new_n245_), .B(G15gat), .Z(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT30), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT31), .ZN(new_n248_));
  XOR2_X1   g047(.A(new_n244_), .B(new_n248_), .Z(new_n249_));
  XNOR2_X1  g048(.A(G1gat), .B(G29gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(G85gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT0), .B(G57gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n251_), .B(new_n252_), .Z(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT88), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G155gat), .A2(G162gat), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(G155gat), .A2(G162gat), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT87), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G141gat), .A2(G148gat), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n260_), .B1(new_n261_), .B2(KEYINPUT85), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT2), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT85), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n264_), .B1(new_n263_), .B2(KEYINPUT87), .ZN(new_n265_));
  AOI22_X1  g064(.A1(new_n262_), .A2(new_n263_), .B1(new_n265_), .B2(new_n261_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(G141gat), .A2(G148gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT3), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n259_), .B1(new_n266_), .B2(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n256_), .A2(KEYINPUT1), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT1), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n272_), .B1(G155gat), .B2(G162gat), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n271_), .B1(new_n256_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT86), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n261_), .A2(KEYINPUT85), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n264_), .A2(G141gat), .A3(G148gat), .ZN(new_n277_));
  OR2_X1    g076(.A1(G141gat), .A2(G148gat), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n276_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  NOR3_X1   g078(.A1(new_n274_), .A2(new_n275_), .A3(new_n279_), .ZN(new_n280_));
  AND3_X1   g079(.A1(new_n276_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n272_), .A2(G155gat), .A3(G162gat), .ZN(new_n282_));
  INV_X1    g081(.A(G155gat), .ZN(new_n283_));
  INV_X1    g082(.A(G162gat), .ZN(new_n284_));
  AOI21_X1  g083(.A(KEYINPUT1), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n282_), .B1(new_n285_), .B2(new_n257_), .ZN(new_n286_));
  AOI21_X1  g085(.A(KEYINPUT86), .B1(new_n281_), .B2(new_n286_), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n255_), .B(new_n270_), .C1(new_n280_), .C2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n275_), .B1(new_n274_), .B2(new_n279_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n281_), .A2(new_n286_), .A3(KEYINPUT86), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n255_), .B1(new_n292_), .B2(new_n270_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n289_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT98), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT4), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n294_), .A2(new_n295_), .A3(new_n296_), .A4(new_n243_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n270_), .B1(new_n280_), .B2(new_n287_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT88), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n299_), .A2(new_n296_), .A3(new_n288_), .A4(new_n243_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT98), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n297_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT99), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n299_), .A2(new_n288_), .A3(new_n243_), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n298_), .A2(new_n243_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(KEYINPUT4), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G225gat), .A2(G233gat), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n307_), .B(KEYINPUT97), .Z(new_n308_));
  NAND4_X1  g107(.A1(new_n302_), .A2(new_n303_), .A3(new_n306_), .A4(new_n308_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n304_), .A2(new_n305_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(new_n307_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n306_), .A2(new_n308_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n303_), .B1(new_n314_), .B2(new_n302_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n254_), .B1(new_n312_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT102), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n300_), .B(new_n295_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT99), .B1(new_n318_), .B2(new_n313_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n319_), .A2(new_n253_), .A3(new_n309_), .A4(new_n311_), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n316_), .A2(new_n317_), .A3(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n317_), .B1(new_n316_), .B2(new_n320_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n249_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT89), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT28), .B1(new_n294_), .B2(KEYINPUT29), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n299_), .A2(new_n288_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT28), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT29), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G22gat), .B(G50gat), .ZN(new_n330_));
  AND3_X1   g129(.A1(new_n325_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n330_), .B1(new_n325_), .B2(new_n329_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n324_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  XOR2_X1   g132(.A(G211gat), .B(G218gat), .Z(new_n334_));
  OR2_X1    g133(.A1(G197gat), .A2(G204gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G197gat), .A2(G204gat), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n334_), .A2(KEYINPUT21), .A3(new_n335_), .A4(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n335_), .A2(KEYINPUT21), .A3(new_n336_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT21), .ZN(new_n339_));
  AND2_X1   g138(.A1(G197gat), .A2(G204gat), .ZN(new_n340_));
  NOR2_X1   g139(.A1(G197gat), .A2(G204gat), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n339_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G211gat), .B(G218gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n338_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(KEYINPUT91), .B1(new_n337_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n337_), .A2(new_n344_), .A3(KEYINPUT91), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G228gat), .A2(G233gat), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n349_), .B(KEYINPUT90), .Z(new_n350_));
  NOR2_X1   g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n351_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT93), .ZN(new_n353_));
  INV_X1    g152(.A(new_n349_), .ZN(new_n354_));
  XOR2_X1   g153(.A(KEYINPUT92), .B(KEYINPUT29), .Z(new_n355_));
  AND2_X1   g154(.A1(new_n298_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n337_), .A2(new_n344_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n353_), .B(new_n354_), .C1(new_n356_), .C2(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n358_), .B1(new_n298_), .B2(new_n355_), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT93), .B1(new_n360_), .B2(new_n349_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n352_), .A2(new_n359_), .A3(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G78gat), .B(G106gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT94), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n362_), .A2(new_n365_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n352_), .A2(new_n359_), .A3(new_n364_), .A4(new_n361_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n330_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n329_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n327_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n369_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n325_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(new_n373_), .A3(KEYINPUT89), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n333_), .A2(new_n368_), .A3(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n331_), .A2(new_n332_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n352_), .A2(new_n361_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n377_), .A2(KEYINPUT95), .A3(new_n364_), .A4(new_n359_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT95), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n367_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n362_), .A2(new_n363_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n376_), .A2(new_n378_), .A3(new_n380_), .A4(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n375_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT96), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT103), .ZN(new_n385_));
  XOR2_X1   g184(.A(G8gat), .B(G36gat), .Z(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT18), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G64gat), .B(G92gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n337_), .A2(new_n344_), .A3(KEYINPUT91), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n390_), .A2(new_n345_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n391_), .B1(new_n235_), .B2(new_n226_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G226gat), .A2(G233gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT19), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT20), .ZN(new_n396_));
  NOR2_X1   g195(.A1(G183gat), .A2(G190gat), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n397_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n232_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT26), .B(G190gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n217_), .A2(new_n400_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n401_), .A2(new_n206_), .A3(new_n212_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n228_), .A2(new_n229_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n399_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n396_), .B1(new_n405_), .B2(new_n358_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n392_), .A2(new_n395_), .A3(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT20), .B1(new_n405_), .B2(new_n358_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n408_), .B1(new_n348_), .B2(new_n236_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n389_), .B(new_n407_), .C1(new_n409_), .C2(new_n395_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT27), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT100), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n401_), .A2(new_n206_), .A3(new_n212_), .ZN(new_n413_));
  OAI22_X1  g212(.A1(new_n413_), .A2(new_n403_), .B1(new_n232_), .B2(new_n398_), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT20), .B1(new_n414_), .B2(new_n357_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n219_), .A2(new_n225_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n213_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(new_n234_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n415_), .B1(new_n419_), .B2(new_n391_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n412_), .B1(new_n420_), .B2(new_n395_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n395_), .B1(new_n392_), .B2(new_n406_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT100), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n348_), .A2(new_n418_), .A3(new_n234_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n396_), .B1(new_n414_), .B2(new_n357_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n421_), .B(new_n423_), .C1(new_n394_), .C2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n389_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n411_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n392_), .A2(new_n395_), .A3(new_n406_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n395_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n428_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(KEYINPUT27), .B1(new_n432_), .B2(new_n410_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n385_), .B1(new_n429_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n433_), .ZN(new_n435_));
  OAI22_X1  g234(.A1(new_n422_), .A2(KEYINPUT100), .B1(new_n426_), .B2(new_n394_), .ZN(new_n436_));
  NOR3_X1   g235(.A1(new_n420_), .A2(new_n412_), .A3(new_n395_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n438_), .A2(new_n389_), .ZN(new_n439_));
  OAI211_X1 g238(.A(KEYINPUT103), .B(new_n435_), .C1(new_n439_), .C2(new_n411_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n434_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT96), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n375_), .A2(new_n382_), .A3(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n384_), .A2(new_n441_), .A3(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n323_), .A2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n321_), .A2(new_n322_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n429_), .A2(new_n433_), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n375_), .A2(new_n382_), .A3(new_n442_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n442_), .B1(new_n375_), .B2(new_n382_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n447_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n316_), .A2(new_n320_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n389_), .A2(KEYINPUT32), .ZN(new_n452_));
  NOR3_X1   g251(.A1(new_n430_), .A2(new_n431_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n452_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT101), .B1(new_n438_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT101), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n427_), .A2(new_n456_), .A3(new_n452_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n453_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT33), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n254_), .A2(new_n459_), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n319_), .A2(new_n311_), .A3(new_n309_), .A4(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n432_), .A2(new_n410_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n302_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n253_), .B1(new_n310_), .B2(new_n308_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n462_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n461_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n320_), .A2(new_n459_), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n451_), .A2(new_n458_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n384_), .A2(new_n443_), .ZN(new_n469_));
  OAI22_X1  g268(.A1(new_n446_), .A2(new_n450_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n249_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n445_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G229gat), .A2(G233gat), .ZN(new_n473_));
  INV_X1    g272(.A(G1gat), .ZN(new_n474_));
  INV_X1    g273(.A(G8gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT14), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT72), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT72), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n478_), .B(KEYINPUT14), .C1(new_n474_), .C2(new_n475_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G15gat), .B(G22gat), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n477_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT73), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G1gat), .B(G8gat), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n482_), .A2(new_n483_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G29gat), .B(G36gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G43gat), .B(G50gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n486_), .A2(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n489_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n473_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(G113gat), .B(G141gat), .Z(new_n495_));
  XNOR2_X1  g294(.A(G169gat), .B(G197gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT80), .B(KEYINPUT81), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n497_), .B(new_n498_), .Z(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n500_), .A2(KEYINPUT79), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n482_), .B(new_n483_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n489_), .B(KEYINPUT15), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT77), .B1(new_n503_), .B2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT77), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n486_), .A2(new_n507_), .A3(new_n504_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n473_), .B(KEYINPUT78), .Z(new_n510_));
  NAND2_X1  g309(.A1(new_n492_), .A2(new_n510_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n494_), .B(new_n502_), .C1(new_n509_), .C2(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n511_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n501_), .B1(new_n513_), .B2(new_n493_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n472_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G99gat), .A2(G106gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT6), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G85gat), .A2(G92gat), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n520_), .A2(KEYINPUT9), .ZN(new_n521_));
  OR2_X1    g320(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n522_));
  INV_X1    g321(.A(G106gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n522_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(G85gat), .ZN(new_n526_));
  INV_X1    g325(.A(G92gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n528_), .A2(KEYINPUT9), .A3(new_n520_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n519_), .A2(new_n521_), .A3(new_n525_), .A4(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n528_), .A2(new_n520_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT6), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n518_), .B(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT7), .ZN(new_n535_));
  INV_X1    g334(.A(G99gat), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n535_), .A2(new_n536_), .A3(new_n523_), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n532_), .B1(new_n534_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT8), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n533_), .B1(G99gat), .B2(G106gat), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n518_), .A2(KEYINPUT6), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n538_), .B(new_n537_), .C1(new_n542_), .C2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT8), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(new_n545_), .A3(new_n532_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n531_), .B1(new_n541_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT66), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n544_), .A2(new_n545_), .A3(new_n532_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n545_), .B1(new_n544_), .B2(new_n532_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n530_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT66), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n549_), .A2(new_n553_), .A3(new_n504_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT70), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n555_), .B1(new_n547_), .B2(new_n489_), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n554_), .A2(KEYINPUT69), .A3(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G232gat), .A2(G233gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT35), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n554_), .A2(new_n556_), .ZN(new_n562_));
  AOI22_X1  g361(.A1(new_n557_), .A2(new_n560_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n560_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT69), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n564_), .B1(new_n562_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G190gat), .B(G218gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G134gat), .B(G162gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n570_), .A2(KEYINPUT36), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n567_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT37), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n570_), .B(KEYINPUT36), .Z(new_n574_));
  NAND3_X1  g373(.A1(new_n563_), .A2(new_n566_), .A3(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n572_), .A2(new_n573_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n571_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n577_), .B1(new_n563_), .B2(new_n566_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n563_), .A2(new_n566_), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n574_), .B(KEYINPUT71), .Z(new_n580_));
  AOI21_X1  g379(.A(new_n578_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n576_), .B1(new_n581_), .B2(new_n573_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT74), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n486_), .B(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(G71gat), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT64), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT64), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(G71gat), .ZN(new_n589_));
  INV_X1    g388(.A(G78gat), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n587_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n588_), .A2(G71gat), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n586_), .A2(KEYINPUT64), .ZN(new_n593_));
  OAI21_X1  g392(.A(G78gat), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(G64gat), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(G57gat), .ZN(new_n596_));
  INV_X1    g395(.A(G57gat), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(G64gat), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n596_), .A2(new_n598_), .A3(KEYINPUT11), .ZN(new_n599_));
  AOI21_X1  g398(.A(KEYINPUT11), .B1(new_n596_), .B2(new_n598_), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n591_), .B(new_n594_), .C1(new_n599_), .C2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n596_), .A2(new_n598_), .A3(KEYINPUT11), .ZN(new_n602_));
  INV_X1    g401(.A(new_n591_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n590_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n602_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n601_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n585_), .A2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n503_), .B(new_n584_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n601_), .A2(new_n605_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT17), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G127gat), .B(G155gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT16), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G183gat), .B(G211gat), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n613_), .B(new_n614_), .Z(new_n615_));
  NAND4_X1  g414(.A1(new_n607_), .A2(new_n610_), .A3(new_n611_), .A4(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(KEYINPUT75), .B1(new_n607_), .B2(new_n610_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n615_), .A2(new_n611_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n618_), .ZN(new_n620_));
  AOI211_X1 g419(.A(KEYINPUT75), .B(new_n620_), .C1(new_n607_), .C2(new_n610_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n616_), .B1(new_n619_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n582_), .A2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT76), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G230gat), .A2(G233gat), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n547_), .A2(new_n606_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n552_), .A2(new_n609_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n626_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n629_), .A2(KEYINPUT65), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(KEYINPUT65), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT12), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n606_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n549_), .A2(new_n553_), .A3(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n632_), .B1(new_n547_), .B2(new_n606_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT67), .ZN(new_n637_));
  AOI211_X1 g436(.A(new_n637_), .B(new_n626_), .C1(new_n547_), .C2(new_n606_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n541_), .A2(new_n546_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n639_), .A2(new_n606_), .A3(new_n530_), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT67), .B1(new_n640_), .B2(new_n625_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n638_), .A2(new_n641_), .ZN(new_n642_));
  OAI22_X1  g441(.A1(new_n630_), .A2(new_n631_), .B1(new_n636_), .B2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(G120gat), .B(G148gat), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT5), .ZN(new_n645_));
  XOR2_X1   g444(.A(G176gat), .B(G204gat), .Z(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n643_), .B(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n648_), .B1(KEYINPUT68), .B2(KEYINPUT13), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n643_), .A2(new_n647_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n643_), .A2(new_n647_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(KEYINPUT68), .B(KEYINPUT13), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n651_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n649_), .A2(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n624_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n517_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n451_), .A2(KEYINPUT102), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n316_), .A2(new_n317_), .A3(new_n320_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n657_), .A2(G1gat), .A3(new_n660_), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n661_), .A2(KEYINPUT38), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(KEYINPUT38), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n572_), .A2(new_n575_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n472_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n622_), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n655_), .A2(new_n667_), .A3(new_n516_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(G1gat), .B1(new_n669_), .B2(new_n660_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n662_), .A2(new_n663_), .A3(new_n670_), .ZN(G1324gat));
  INV_X1    g470(.A(new_n441_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n666_), .A2(new_n672_), .A3(new_n668_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT39), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(new_n674_), .A3(G8gat), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n674_), .B1(new_n673_), .B2(G8gat), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n672_), .A2(new_n475_), .ZN(new_n678_));
  OAI22_X1  g477(.A1(new_n676_), .A2(new_n677_), .B1(new_n657_), .B2(new_n678_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g479(.A(G15gat), .B1(new_n669_), .B2(new_n471_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT41), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n657_), .A2(G15gat), .A3(new_n471_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1326gat));
  NOR2_X1   g483(.A1(new_n448_), .A2(new_n449_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G22gat), .B1(new_n669_), .B2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT42), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n685_), .A2(G22gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n687_), .B1(new_n657_), .B2(new_n688_), .ZN(G1327gat));
  NAND2_X1  g488(.A1(new_n667_), .A2(new_n665_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n690_), .A2(new_n655_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n517_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(G29gat), .B1(new_n693_), .B2(new_n446_), .ZN(new_n694_));
  XOR2_X1   g493(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n695_));
  XOR2_X1   g494(.A(KEYINPUT105), .B(KEYINPUT43), .Z(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n697_), .B1(new_n472_), .B2(new_n582_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n582_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n660_), .A2(new_n469_), .A3(new_n447_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n451_), .A2(new_n458_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n466_), .A2(new_n467_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n685_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n249_), .B1(new_n701_), .B2(new_n704_), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n699_), .B(new_n700_), .C1(new_n705_), .C2(new_n445_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n698_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n649_), .A2(new_n654_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n708_), .A2(new_n667_), .A3(new_n515_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT104), .Z(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n695_), .B1(new_n707_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713_));
  AOI211_X1 g512(.A(new_n713_), .B(new_n710_), .C1(new_n698_), .C2(new_n706_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n712_), .A2(new_n714_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n446_), .A2(G29gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n694_), .B1(new_n715_), .B2(new_n716_), .ZN(G1328gat));
  NOR3_X1   g516(.A1(new_n692_), .A2(G36gat), .A3(new_n441_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT45), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n710_), .B1(new_n698_), .B2(new_n706_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT44), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n722_), .B1(new_n721_), .B2(new_n695_), .ZN(new_n723_));
  OAI21_X1  g522(.A(G36gat), .B1(new_n723_), .B2(new_n441_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n720_), .A2(new_n724_), .A3(KEYINPUT46), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT46), .ZN(new_n726_));
  INV_X1    g525(.A(G36gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n727_), .B1(new_n715_), .B2(new_n672_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n726_), .B1(new_n728_), .B2(new_n719_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n725_), .A2(new_n729_), .ZN(G1329gat));
  NAND3_X1  g529(.A1(new_n715_), .A2(G43gat), .A3(new_n249_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n238_), .B1(new_n692_), .B2(new_n471_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n731_), .A2(new_n732_), .A3(new_n734_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(G1330gat));
  NOR3_X1   g537(.A1(new_n692_), .A2(G50gat), .A3(new_n685_), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n722_), .B(new_n469_), .C1(new_n721_), .C2(new_n695_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n740_), .B2(G50gat), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT108), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  AOI211_X1 g542(.A(KEYINPUT108), .B(new_n739_), .C1(new_n740_), .C2(G50gat), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1331gat));
  NOR3_X1   g544(.A1(new_n708_), .A2(new_n667_), .A3(new_n515_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n666_), .A2(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G57gat), .B1(new_n747_), .B2(new_n660_), .ZN(new_n748_));
  NOR4_X1   g547(.A1(new_n472_), .A2(new_n624_), .A3(new_n515_), .A4(new_n708_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n749_), .A2(new_n597_), .A3(new_n446_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(G1332gat));
  OAI21_X1  g550(.A(G64gat), .B1(new_n747_), .B2(new_n441_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT48), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n749_), .A2(new_n595_), .A3(new_n672_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1333gat));
  NAND3_X1  g554(.A1(new_n666_), .A2(new_n249_), .A3(new_n746_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(G71gat), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT49), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n749_), .A2(new_n586_), .A3(new_n249_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT109), .ZN(G1334gat));
  OAI21_X1  g560(.A(G78gat), .B1(new_n747_), .B2(new_n685_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n762_), .B(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n685_), .A2(G78gat), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT111), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n749_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n764_), .A2(new_n767_), .ZN(G1335gat));
  OR4_X1    g567(.A1(new_n472_), .A2(new_n515_), .A3(new_n708_), .A4(new_n690_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n526_), .B1(new_n769_), .B2(new_n660_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT112), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n655_), .A2(new_n516_), .A3(new_n667_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT113), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n707_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT114), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n707_), .A2(new_n777_), .A3(new_n774_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n660_), .A2(new_n526_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n771_), .B1(new_n779_), .B2(new_n780_), .ZN(G1336gat));
  OAI21_X1  g580(.A(new_n527_), .B1(new_n769_), .B2(new_n441_), .ZN(new_n782_));
  XOR2_X1   g581(.A(new_n782_), .B(KEYINPUT115), .Z(new_n783_));
  NOR2_X1   g582(.A1(new_n441_), .A2(new_n527_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n779_), .B2(new_n784_), .ZN(G1337gat));
  NAND3_X1  g584(.A1(new_n249_), .A2(new_n522_), .A3(new_n524_), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n769_), .A2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n471_), .B1(new_n776_), .B2(new_n778_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n788_), .B2(new_n536_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT51), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n791_), .B(new_n787_), .C1(new_n788_), .C2(new_n536_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(G1338gat));
  AOI211_X1 g592(.A(new_n685_), .B(new_n773_), .C1(new_n698_), .C2(new_n706_), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT116), .B1(new_n794_), .B2(new_n523_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n707_), .A2(new_n469_), .A3(new_n774_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n797_), .A3(G106gat), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n795_), .A2(KEYINPUT52), .A3(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n800_));
  OAI211_X1 g599(.A(KEYINPUT116), .B(new_n800_), .C1(new_n794_), .C2(new_n523_), .ZN(new_n801_));
  OR3_X1    g600(.A1(new_n769_), .A2(G106gat), .A3(new_n685_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT53), .B1(new_n799_), .B2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n795_), .A2(KEYINPUT52), .A3(new_n798_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n805_), .A2(new_n806_), .A3(new_n801_), .A4(new_n802_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n804_), .A2(new_n807_), .ZN(G1339gat));
  NAND2_X1  g607(.A1(new_n622_), .A2(new_n516_), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n655_), .A2(new_n809_), .A3(new_n699_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n810_), .B(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n642_), .B2(new_n636_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n637_), .B1(new_n628_), .B2(new_n626_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n640_), .A2(KEYINPUT67), .A3(new_n625_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n817_), .A2(KEYINPUT55), .A3(new_n635_), .A4(new_n634_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n626_), .B1(new_n636_), .B2(new_n628_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n814_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n647_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n650_), .B1(new_n821_), .B2(KEYINPUT56), .ZN(new_n822_));
  INV_X1    g621(.A(new_n510_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n492_), .A2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n824_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n823_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n499_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n500_), .B1(new_n513_), .B2(new_n493_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT56), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n820_), .A2(new_n830_), .A3(new_n647_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n822_), .A2(KEYINPUT58), .A3(new_n829_), .A4(new_n831_), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n832_), .A2(KEYINPUT118), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n821_), .A2(KEYINPUT56), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n834_), .A2(new_n829_), .A3(new_n651_), .A4(new_n831_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT117), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT58), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT117), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n822_), .A2(new_n838_), .A3(new_n829_), .A4(new_n831_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n836_), .A2(new_n837_), .A3(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n582_), .B1(new_n832_), .B2(KEYINPUT118), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n833_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n834_), .A2(new_n515_), .A3(new_n651_), .A4(new_n831_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n648_), .A2(new_n829_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n664_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n845_), .A2(KEYINPUT57), .A3(new_n664_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n667_), .B1(new_n842_), .B2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n812_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n444_), .A2(new_n660_), .A3(new_n471_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n852_), .A2(new_n853_), .A3(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n854_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n842_), .B2(new_n850_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n833_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n859_), .A2(KEYINPUT119), .A3(new_n848_), .A4(new_n849_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n858_), .A2(new_n667_), .A3(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n856_), .B1(new_n861_), .B2(new_n812_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n855_), .B(new_n515_), .C1(new_n862_), .C2(new_n853_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(G113gat), .ZN(new_n864_));
  INV_X1    g663(.A(G113gat), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n862_), .A2(new_n865_), .A3(new_n515_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT120), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n864_), .A2(new_n869_), .A3(new_n866_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n870_), .ZN(G1340gat));
  INV_X1    g670(.A(new_n862_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(KEYINPUT59), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT121), .B(G120gat), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n655_), .A2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n862_), .B1(KEYINPUT60), .B2(new_n875_), .ZN(new_n876_));
  AND4_X1   g675(.A1(new_n655_), .A2(new_n873_), .A3(new_n855_), .A4(new_n876_), .ZN(new_n877_));
  OAI22_X1  g676(.A1(new_n877_), .A2(new_n874_), .B1(KEYINPUT60), .B2(new_n876_), .ZN(G1341gat));
  INV_X1    g677(.A(G127gat), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n879_), .B1(new_n872_), .B2(new_n667_), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n880_), .A2(KEYINPUT122), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(KEYINPUT122), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n873_), .A2(new_n855_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n667_), .A2(new_n879_), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n881_), .A2(new_n882_), .B1(new_n884_), .B2(new_n885_), .ZN(G1342gat));
  OAI21_X1  g685(.A(G134gat), .B1(new_n883_), .B2(new_n582_), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n664_), .A2(G134gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n872_), .B2(new_n888_), .ZN(G1343gat));
  NAND2_X1  g688(.A1(new_n861_), .A2(new_n812_), .ZN(new_n890_));
  NOR4_X1   g689(.A1(new_n660_), .A2(new_n685_), .A3(new_n672_), .A4(new_n249_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n515_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g694(.A1(new_n892_), .A2(new_n708_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(KEYINPUT123), .B(G148gat), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n896_), .B(new_n897_), .ZN(G1345gat));
  XNOR2_X1  g697(.A(KEYINPUT61), .B(G155gat), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(KEYINPUT124), .B1(new_n892_), .B2(new_n667_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n892_), .A2(KEYINPUT124), .A3(new_n667_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n900_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n903_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n905_), .A2(new_n901_), .A3(new_n899_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n906_), .ZN(G1346gat));
  OAI21_X1  g706(.A(G162gat), .B1(new_n892_), .B2(new_n582_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n665_), .A2(new_n284_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n892_), .B2(new_n909_), .ZN(G1347gat));
  INV_X1    g709(.A(KEYINPUT62), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n469_), .B1(new_n812_), .B2(new_n851_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n323_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n672_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n912_), .A2(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(new_n516_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT22), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n911_), .B1(new_n917_), .B2(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(G169gat), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n204_), .B1(new_n917_), .B2(new_n911_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n919_), .B2(new_n921_), .ZN(G1348gat));
  INV_X1    g721(.A(new_n916_), .ZN(new_n923_));
  AOI21_X1  g722(.A(G176gat), .B1(new_n923_), .B2(new_n655_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n469_), .B1(new_n861_), .B2(new_n812_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n914_), .A2(new_n205_), .A3(new_n708_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n924_), .B1(new_n925_), .B2(new_n926_), .ZN(G1349gat));
  NOR2_X1   g726(.A1(new_n914_), .A2(new_n667_), .ZN(new_n928_));
  AOI21_X1  g727(.A(G183gat), .B1(new_n925_), .B2(new_n928_), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n914_), .A2(new_n217_), .A3(new_n667_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n929_), .B1(new_n912_), .B2(new_n930_), .ZN(G1350gat));
  OAI21_X1  g730(.A(G190gat), .B1(new_n916_), .B2(new_n582_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n665_), .A2(new_n400_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n916_), .B2(new_n933_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT125), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n934_), .B(new_n935_), .ZN(G1351gat));
  NOR4_X1   g735(.A1(new_n446_), .A2(new_n685_), .A3(new_n249_), .A4(new_n441_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n890_), .A2(new_n937_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n938_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(new_n515_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g740(.A1(new_n938_), .A2(new_n708_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(KEYINPUT126), .B(G204gat), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n942_), .B(new_n943_), .ZN(G1353gat));
  NAND2_X1  g743(.A1(new_n939_), .A2(new_n622_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n946_));
  AND2_X1   g745(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n947_));
  NOR3_X1   g746(.A1(new_n945_), .A2(new_n946_), .A3(new_n947_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n948_), .B1(new_n945_), .B2(new_n946_), .ZN(G1354gat));
  AND3_X1   g748(.A1(new_n939_), .A2(G218gat), .A3(new_n699_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n938_), .A2(new_n664_), .ZN(new_n951_));
  OR2_X1    g750(.A1(new_n951_), .A2(KEYINPUT127), .ZN(new_n952_));
  AOI21_X1  g751(.A(G218gat), .B1(new_n951_), .B2(KEYINPUT127), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n950_), .B1(new_n952_), .B2(new_n953_), .ZN(G1355gat));
endmodule


