//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 1 0 0 0 0 1 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n794_, new_n795_, new_n797_,
    new_n798_, new_n799_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n959_,
    new_n960_, new_n961_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n978_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n986_, new_n987_, new_n988_;
  NAND3_X1  g000(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n202_));
  INV_X1    g001(.A(G92gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n203_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n202_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT6), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT10), .B(G99gat), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n214_), .A2(G106gat), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n209_), .A2(new_n212_), .A3(new_n213_), .A4(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT7), .ZN(new_n217_));
  INV_X1    g016(.A(G99gat), .ZN(new_n218_));
  INV_X1    g017(.A(G106gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n220_), .A2(new_n212_), .A3(new_n213_), .A4(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT8), .ZN(new_n223_));
  XOR2_X1   g022(.A(G85gat), .B(G92gat), .Z(new_n224_));
  AND3_X1   g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n223_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n216_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT66), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G29gat), .B(G36gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G43gat), .B(G50gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT15), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n216_), .B(new_n233_), .C1(new_n226_), .C2(new_n225_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n228_), .A2(new_n232_), .A3(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT70), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT70), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n228_), .A2(new_n237_), .A3(new_n232_), .A4(new_n234_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G232gat), .A2(G233gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT34), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT35), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n227_), .ZN(new_n246_));
  AOI22_X1  g045(.A1(new_n246_), .A2(new_n231_), .B1(new_n243_), .B2(new_n242_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n239_), .A2(new_n245_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n245_), .B1(new_n239_), .B2(new_n247_), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT71), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n250_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT71), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(new_n253_), .A3(new_n248_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G190gat), .B(G218gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G134gat), .B(G162gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n257_), .B(KEYINPUT36), .Z(new_n258_));
  NAND3_X1  g057(.A1(new_n251_), .A2(new_n254_), .A3(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n257_), .A2(KEYINPUT36), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n252_), .A2(new_n260_), .A3(new_n248_), .ZN(new_n261_));
  AOI21_X1  g060(.A(KEYINPUT37), .B1(new_n259_), .B2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n258_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n263_), .A2(new_n261_), .A3(KEYINPUT37), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G1gat), .B(G8gat), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n267_), .A2(KEYINPUT72), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(KEYINPUT72), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G15gat), .B(G22gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G1gat), .A2(G8gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT14), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n270_), .A2(new_n274_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n268_), .A2(new_n273_), .A3(new_n271_), .A4(new_n269_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G231gat), .A2(G233gat), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n277_), .B(new_n278_), .Z(new_n279_));
  XNOR2_X1  g078(.A(G57gat), .B(G64gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G71gat), .B(G78gat), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n280_), .A2(new_n281_), .A3(KEYINPUT11), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(KEYINPUT11), .ZN(new_n283_));
  INV_X1    g082(.A(new_n281_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n280_), .A2(KEYINPUT11), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n282_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT67), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n279_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT17), .ZN(new_n291_));
  XOR2_X1   g090(.A(G127gat), .B(G155gat), .Z(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT16), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G183gat), .B(G211gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  NOR3_X1   g094(.A1(new_n290_), .A2(new_n291_), .A3(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n279_), .A2(new_n289_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n295_), .B(new_n291_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n299_), .B1(new_n279_), .B2(new_n287_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n300_), .B1(new_n287_), .B2(new_n279_), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n266_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT69), .ZN(new_n304_));
  INV_X1    g103(.A(new_n287_), .ZN(new_n305_));
  AOI21_X1  g104(.A(KEYINPUT12), .B1(new_n227_), .B2(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n306_), .B1(new_n246_), .B2(new_n287_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G230gat), .A2(G233gat), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n289_), .A2(new_n228_), .A3(KEYINPUT12), .A4(new_n234_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT65), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n311_), .B1(new_n227_), .B2(new_n305_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n312_), .B1(new_n227_), .B2(new_n305_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n246_), .A2(new_n311_), .A3(new_n287_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n313_), .A2(G230gat), .A3(G233gat), .A4(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G120gat), .B(G148gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT5), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G176gat), .B(G204gat), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n317_), .B(new_n318_), .Z(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n310_), .A2(new_n315_), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT68), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n320_), .B1(new_n310_), .B2(new_n315_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n310_), .A2(new_n315_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(new_n319_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n326_), .A2(KEYINPUT68), .A3(new_n321_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n324_), .A2(new_n327_), .A3(KEYINPUT13), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(KEYINPUT13), .B1(new_n327_), .B2(new_n324_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n304_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n324_), .A2(new_n327_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT13), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n334_), .A2(KEYINPUT69), .A3(new_n328_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n331_), .A2(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n303_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(G169gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT22), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT22), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(G169gat), .ZN(new_n341_));
  INV_X1    g140(.A(G176gat), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n339_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT78), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT79), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G169gat), .A2(G176gat), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n339_), .A2(new_n341_), .A3(new_n347_), .A4(new_n342_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .A4(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G183gat), .A2(G190gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT77), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n352_), .A2(G183gat), .A3(G190gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT23), .ZN(new_n355_));
  INV_X1    g154(.A(G183gat), .ZN(new_n356_));
  INV_X1    g155(.A(G190gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n355_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n349_), .A2(new_n361_), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n343_), .A2(KEYINPUT78), .B1(G169gat), .B2(G176gat), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n345_), .B1(new_n363_), .B2(new_n348_), .ZN(new_n364_));
  AND3_X1   g163(.A1(new_n350_), .A2(KEYINPUT76), .A3(KEYINPUT23), .ZN(new_n365_));
  AOI21_X1  g164(.A(KEYINPUT76), .B1(new_n350_), .B2(KEYINPUT23), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT23), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n352_), .B1(G183gat), .B2(G190gat), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n350_), .A2(KEYINPUT77), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n368_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n367_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n356_), .A2(KEYINPUT25), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT25), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(G183gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n357_), .A2(KEYINPUT26), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT26), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(G190gat), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n373_), .A2(new_n375_), .A3(new_n376_), .A4(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n338_), .A2(new_n342_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n380_), .A2(KEYINPUT24), .A3(new_n346_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(KEYINPUT75), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n372_), .A2(new_n382_), .ZN(new_n383_));
  NOR3_X1   g182(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT25), .B(G183gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT26), .B(G190gat), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n386_), .A2(new_n387_), .B1(new_n389_), .B2(new_n346_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n385_), .B1(new_n390_), .B2(KEYINPUT75), .ZN(new_n391_));
  OAI22_X1  g190(.A1(new_n362_), .A2(new_n364_), .B1(new_n383_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G227gat), .A2(G233gat), .ZN(new_n393_));
  XOR2_X1   g192(.A(new_n393_), .B(G71gat), .Z(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(new_n218_), .ZN(new_n395_));
  OR2_X1    g194(.A1(new_n392_), .A2(new_n395_), .ZN(new_n396_));
  XOR2_X1   g195(.A(KEYINPUT82), .B(KEYINPUT31), .Z(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT83), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n392_), .A2(new_n395_), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n396_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n398_), .B1(new_n396_), .B2(new_n399_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G15gat), .B(G43gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT80), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT30), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G113gat), .B(G120gat), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(G134gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(G127gat), .ZN(new_n408_));
  INV_X1    g207(.A(G127gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(G134gat), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT81), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n408_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n411_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n406_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n409_), .A2(G134gat), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n407_), .A2(G127gat), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT81), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n408_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n417_), .A2(new_n418_), .A3(new_n405_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n414_), .A2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n404_), .B(new_n420_), .ZN(new_n421_));
  OR3_X1    g220(.A1(new_n400_), .A2(new_n401_), .A3(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n421_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(G211gat), .B(G218gat), .Z(new_n426_));
  INV_X1    g225(.A(KEYINPUT21), .ZN(new_n427_));
  INV_X1    g226(.A(G204gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(G197gat), .ZN(new_n429_));
  INV_X1    g228(.A(G197gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(G204gat), .ZN(new_n431_));
  AND2_X1   g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n426_), .B1(new_n427_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n429_), .A2(KEYINPUT87), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT87), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n435_), .A2(new_n428_), .A3(G197gat), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n434_), .A2(new_n436_), .A3(new_n431_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT21), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n432_), .A2(new_n427_), .ZN(new_n439_));
  AOI22_X1  g238(.A1(new_n433_), .A2(new_n438_), .B1(new_n439_), .B2(new_n426_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n392_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G226gat), .A2(G233gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT91), .ZN(new_n444_));
  XOR2_X1   g243(.A(KEYINPUT90), .B(KEYINPUT19), .Z(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n359_), .B1(new_n354_), .B2(KEYINPUT23), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT92), .B1(new_n447_), .B2(new_n385_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n368_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT92), .ZN(new_n450_));
  NOR4_X1   g249(.A1(new_n449_), .A2(new_n450_), .A3(new_n384_), .A4(new_n359_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n390_), .B1(new_n448_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n343_), .A2(new_n346_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n453_), .B1(new_n372_), .B2(new_n358_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n452_), .A2(new_n455_), .A3(new_n440_), .ZN(new_n456_));
  AND4_X1   g255(.A1(KEYINPUT20), .A2(new_n442_), .A3(new_n446_), .A4(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n379_), .A2(new_n381_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n355_), .A2(new_n385_), .A3(new_n360_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(new_n450_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n447_), .A2(KEYINPUT92), .A3(new_n385_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n458_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n441_), .B1(new_n462_), .B2(new_n454_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT93), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT75), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n458_), .A2(new_n465_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n466_), .A2(new_n385_), .A3(new_n382_), .A4(new_n372_), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n467_), .B(new_n440_), .C1(new_n364_), .C2(new_n362_), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n468_), .A2(KEYINPUT20), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n452_), .A2(new_n455_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT93), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(new_n471_), .A3(new_n441_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n464_), .A2(new_n469_), .A3(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n446_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n457_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  XOR2_X1   g274(.A(G8gat), .B(G36gat), .Z(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G64gat), .B(G92gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT95), .B1(new_n475_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT95), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n471_), .B1(new_n470_), .B2(new_n441_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n468_), .A2(KEYINPUT20), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n446_), .B1(new_n486_), .B2(new_n472_), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n483_), .B(new_n480_), .C1(new_n487_), .C2(new_n457_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n475_), .A2(new_n481_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n482_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT27), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(G155gat), .ZN(new_n493_));
  INV_X1    g292(.A(G162gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(new_n494_), .A3(KEYINPUT84), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT84), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n496_), .B1(G155gat), .B2(G162gat), .ZN(new_n497_));
  AOI22_X1  g296(.A1(new_n495_), .A2(new_n497_), .B1(G155gat), .B2(G162gat), .ZN(new_n498_));
  AOI21_X1  g297(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT85), .ZN(new_n500_));
  NOR2_X1   g299(.A1(G141gat), .A2(G148gat), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT3), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n498_), .B1(new_n500_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G155gat), .A2(G162gat), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT1), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n495_), .A2(new_n497_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  AND2_X1   g311(.A1(G141gat), .A2(G148gat), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n513_), .A2(new_n501_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n507_), .A2(new_n515_), .ZN(new_n516_));
  OR3_X1    g315(.A1(new_n516_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n517_));
  OAI21_X1  g316(.A(KEYINPUT28), .B1(new_n516_), .B2(KEYINPUT29), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G22gat), .B(G50gat), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n520_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G228gat), .A2(G233gat), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT86), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n516_), .A2(KEYINPUT29), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n525_), .B1(new_n526_), .B2(new_n441_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT29), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n528_), .B1(new_n507_), .B2(new_n515_), .ZN(new_n529_));
  NOR3_X1   g328(.A1(new_n529_), .A2(KEYINPUT86), .A3(new_n440_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n524_), .B1(new_n527_), .B2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n526_), .A2(new_n525_), .A3(new_n441_), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT86), .B1(new_n529_), .B2(new_n440_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n532_), .A2(new_n533_), .A3(G228gat), .A4(G233gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G78gat), .B(G106gat), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n535_), .B(KEYINPUT88), .Z(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n531_), .A2(new_n534_), .A3(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n537_), .B1(new_n531_), .B2(new_n534_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT89), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n538_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  AOI211_X1 g340(.A(KEYINPUT89), .B(new_n537_), .C1(new_n531_), .C2(new_n534_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n523_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n539_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n531_), .A2(new_n535_), .A3(new_n534_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n544_), .A2(new_n521_), .A3(new_n522_), .A4(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n511_), .A2(new_n508_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n506_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT85), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n499_), .B(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n548_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n514_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n553_), .B1(new_n511_), .B2(new_n510_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n420_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n507_), .A2(new_n515_), .A3(new_n419_), .A4(new_n414_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G225gat), .A2(G233gat), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n555_), .A2(new_n556_), .A3(KEYINPUT4), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT4), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n516_), .A2(new_n562_), .A3(new_n420_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n561_), .A2(new_n559_), .A3(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n560_), .B1(new_n564_), .B2(KEYINPUT96), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT96), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n561_), .A2(new_n566_), .A3(new_n559_), .A4(new_n563_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G1gat), .B(G29gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(G85gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT0), .B(G57gat), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n570_), .B(new_n571_), .Z(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n568_), .A2(new_n573_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n555_), .A2(new_n556_), .A3(KEYINPUT4), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n563_), .A2(new_n559_), .ZN(new_n576_));
  OAI21_X1  g375(.A(KEYINPUT96), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n560_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n577_), .A2(new_n572_), .A3(new_n578_), .A4(new_n567_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT97), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n565_), .A2(KEYINPUT97), .A3(new_n572_), .A4(new_n567_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n574_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n442_), .A2(KEYINPUT20), .A3(new_n456_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n474_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n586_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(new_n480_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n489_), .A2(new_n588_), .A3(KEYINPUT27), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n492_), .A2(new_n547_), .A3(new_n584_), .A4(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n573_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n563_), .A2(new_n558_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n591_), .B1(new_n592_), .B2(new_n561_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n579_), .A2(KEYINPUT33), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT33), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n565_), .A2(new_n595_), .A3(new_n572_), .A4(new_n567_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n593_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n597_), .A2(new_n482_), .A3(new_n488_), .A4(new_n489_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n481_), .A2(KEYINPUT32), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n586_), .B(new_n599_), .C1(new_n473_), .C2(new_n474_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n600_), .B1(new_n475_), .B2(new_n599_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(new_n583_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n547_), .B1(new_n598_), .B2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n590_), .B1(KEYINPUT98), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n598_), .A2(new_n602_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n547_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n605_), .A2(KEYINPUT98), .A3(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n425_), .B1(new_n604_), .B2(new_n607_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n492_), .A2(new_n589_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n425_), .A2(new_n583_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n609_), .A2(KEYINPUT99), .A3(new_n606_), .A4(new_n610_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n606_), .A2(new_n610_), .A3(new_n492_), .A4(new_n589_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT99), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n608_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n232_), .A2(new_n277_), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n275_), .A2(new_n231_), .A3(new_n276_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G229gat), .A2(G233gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT73), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n617_), .A2(new_n619_), .A3(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n231_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n623_));
  OAI211_X1 g422(.A(G229gat), .B(G233gat), .C1(new_n618_), .C2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G113gat), .B(G141gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G169gat), .B(G197gat), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n626_), .B(new_n627_), .Z(new_n628_));
  AND3_X1   g427(.A1(new_n625_), .A2(KEYINPUT74), .A3(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n628_), .B1(new_n625_), .B2(KEYINPUT74), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(KEYINPUT100), .B1(new_n616_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT100), .ZN(new_n633_));
  INV_X1    g432(.A(new_n631_), .ZN(new_n634_));
  AOI211_X1 g433(.A(new_n633_), .B(new_n634_), .C1(new_n608_), .C2(new_n615_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n337_), .B1(new_n632_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT101), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n637_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n584_), .A2(G1gat), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT38), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n640_), .A2(KEYINPUT38), .A3(new_n641_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n259_), .A2(new_n261_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n616_), .A2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT103), .ZN(new_n649_));
  OAI21_X1  g448(.A(KEYINPUT102), .B1(new_n336_), .B2(new_n634_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n331_), .A2(new_n335_), .A3(new_n651_), .A4(new_n631_), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n650_), .A2(new_n302_), .A3(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n649_), .A2(new_n583_), .A3(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(G1gat), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n644_), .A2(new_n645_), .A3(new_n655_), .ZN(G1324gat));
  NOR2_X1   g455(.A1(new_n609_), .A2(G8gat), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n638_), .A2(new_n639_), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n609_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n649_), .A2(new_n659_), .A3(new_n653_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT39), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n660_), .A2(new_n661_), .A3(G8gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n661_), .B1(new_n660_), .B2(G8gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n658_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT40), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  OAI211_X1 g465(.A(KEYINPUT40), .B(new_n658_), .C1(new_n662_), .C2(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1325gat));
  INV_X1    g467(.A(G15gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n640_), .A2(new_n669_), .A3(new_n424_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n649_), .A2(new_n424_), .A3(new_n653_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n671_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT41), .B1(new_n671_), .B2(G15gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n670_), .B1(new_n672_), .B2(new_n673_), .ZN(G1326gat));
  INV_X1    g473(.A(G22gat), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n640_), .A2(new_n675_), .A3(new_n547_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n649_), .A2(new_n547_), .A3(new_n653_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G22gat), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n678_), .A2(KEYINPUT42), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n678_), .A2(KEYINPUT42), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n676_), .B1(new_n679_), .B2(new_n680_), .ZN(G1327gat));
  NOR2_X1   g480(.A1(new_n647_), .A2(new_n302_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n683_), .A2(new_n336_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n605_), .A2(new_n606_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT98), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n603_), .A2(KEYINPUT98), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n688_), .A2(new_n689_), .A3(new_n590_), .ZN(new_n690_));
  AOI22_X1  g489(.A1(new_n690_), .A2(new_n425_), .B1(new_n614_), .B2(new_n611_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n633_), .B1(new_n691_), .B2(new_n634_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n616_), .A2(KEYINPUT100), .A3(new_n631_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n685_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(G29gat), .B1(new_n694_), .B2(new_n583_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n302_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n650_), .A2(new_n696_), .A3(new_n652_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(KEYINPUT43), .B1(new_n266_), .B2(KEYINPUT104), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n691_), .A2(new_n700_), .A3(new_n266_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n264_), .B1(new_n646_), .B2(KEYINPUT37), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n699_), .B1(new_n616_), .B2(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n698_), .B1(new_n701_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n706_), .A2(G29gat), .A3(new_n583_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n700_), .B1(new_n691_), .B2(new_n266_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n616_), .A2(new_n702_), .A3(new_n699_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n710_), .A2(KEYINPUT44), .A3(new_n698_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n695_), .B1(new_n707_), .B2(new_n711_), .ZN(G1328gat));
  XOR2_X1   g511(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n609_), .A2(G36gat), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n684_), .B(new_n715_), .C1(new_n632_), .C2(new_n635_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT106), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT106), .B1(new_n694_), .B2(new_n715_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n714_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n716_), .A2(new_n717_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n694_), .A2(KEYINPUT106), .A3(new_n715_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n722_), .A3(new_n713_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n720_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n725_));
  NOR2_X1   g524(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n706_), .A2(new_n659_), .A3(new_n711_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n727_), .B2(G36gat), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n724_), .A2(new_n725_), .A3(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n725_), .B1(new_n724_), .B2(new_n728_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1329gat));
  INV_X1    g530(.A(G43gat), .ZN(new_n732_));
  INV_X1    g531(.A(new_n694_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(new_n425_), .ZN(new_n734_));
  AOI21_X1  g533(.A(KEYINPUT44), .B1(new_n710_), .B2(new_n698_), .ZN(new_n735_));
  AOI211_X1 g534(.A(new_n705_), .B(new_n697_), .C1(new_n708_), .C2(new_n709_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n425_), .A2(new_n732_), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT108), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  AND4_X1   g538(.A1(KEYINPUT108), .A2(new_n706_), .A3(new_n711_), .A4(new_n738_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n734_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT47), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT47), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n743_), .B(new_n734_), .C1(new_n739_), .C2(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1330gat));
  NAND2_X1  g544(.A1(new_n737_), .A2(new_n547_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(G50gat), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n606_), .A2(G50gat), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT109), .Z(new_n749_));
  OAI21_X1  g548(.A(new_n747_), .B1(new_n733_), .B2(new_n749_), .ZN(G1331gat));
  NAND2_X1  g549(.A1(new_n302_), .A2(new_n634_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n649_), .A2(new_n336_), .A3(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(G57gat), .B1(new_n753_), .B2(new_n584_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n336_), .ZN(new_n755_));
  NOR4_X1   g554(.A1(new_n691_), .A2(new_n631_), .A3(new_n755_), .A4(new_n303_), .ZN(new_n756_));
  INV_X1    g555(.A(G57gat), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(new_n757_), .A3(new_n583_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n754_), .A2(new_n758_), .ZN(G1332gat));
  INV_X1    g558(.A(G64gat), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n756_), .A2(new_n760_), .A3(new_n659_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT48), .ZN(new_n762_));
  INV_X1    g561(.A(new_n753_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n659_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n762_), .B1(new_n764_), .B2(G64gat), .ZN(new_n765_));
  AOI211_X1 g564(.A(KEYINPUT48), .B(new_n760_), .C1(new_n763_), .C2(new_n659_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n761_), .B1(new_n765_), .B2(new_n766_), .ZN(G1333gat));
  NOR2_X1   g566(.A1(new_n425_), .A2(G71gat), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT110), .Z(new_n769_));
  NAND2_X1  g568(.A1(new_n756_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n763_), .A2(new_n424_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT49), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n771_), .A2(new_n772_), .A3(G71gat), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n771_), .B2(G71gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n770_), .B1(new_n773_), .B2(new_n774_), .ZN(G1334gat));
  INV_X1    g574(.A(G78gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n756_), .A2(new_n776_), .A3(new_n547_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT50), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n763_), .A2(new_n547_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(G78gat), .ZN(new_n780_));
  AOI211_X1 g579(.A(KEYINPUT50), .B(new_n776_), .C1(new_n763_), .C2(new_n547_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n777_), .B1(new_n780_), .B2(new_n781_), .ZN(G1335gat));
  NOR2_X1   g581(.A1(new_n691_), .A2(new_n631_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n683_), .A2(new_n755_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(G85gat), .B1(new_n786_), .B2(new_n583_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n755_), .A2(new_n631_), .A3(new_n302_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n710_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n204_), .A2(new_n205_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n583_), .A2(new_n790_), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT111), .Z(new_n792_));
  AOI21_X1  g591(.A(new_n787_), .B1(new_n789_), .B2(new_n792_), .ZN(G1336gat));
  NAND3_X1  g592(.A1(new_n786_), .A2(new_n203_), .A3(new_n659_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n789_), .A2(new_n659_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(new_n203_), .ZN(G1337gat));
  AND2_X1   g595(.A1(new_n789_), .A2(new_n424_), .ZN(new_n797_));
  OR2_X1    g596(.A1(new_n425_), .A2(new_n214_), .ZN(new_n798_));
  OAI22_X1  g597(.A1(new_n797_), .A2(new_n218_), .B1(new_n785_), .B2(new_n798_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n788_), .B(new_n547_), .C1(new_n701_), .C2(new_n703_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n802_), .A2(new_n803_), .A3(G106gat), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n803_), .B1(new_n802_), .B2(G106gat), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n801_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n802_), .A2(G106gat), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(KEYINPUT113), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n802_), .A2(new_n803_), .A3(G106gat), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(KEYINPUT52), .A3(new_n809_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n785_), .A2(G106gat), .A3(new_n606_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(KEYINPUT112), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n806_), .A2(new_n810_), .A3(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT53), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n806_), .A2(new_n810_), .A3(new_n815_), .A4(new_n812_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n816_), .ZN(G1339gat));
  NOR2_X1   g616(.A1(new_n329_), .A2(new_n330_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n818_), .A2(new_n751_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n819_), .A2(new_n820_), .A3(new_n266_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n820_), .B1(new_n819_), .B2(new_n266_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n308_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n310_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n307_), .A2(KEYINPUT55), .A3(new_n308_), .A4(new_n309_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n828_), .A2(KEYINPUT114), .A3(KEYINPUT56), .A4(new_n319_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n631_), .A2(new_n321_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT56), .B1(new_n828_), .B2(new_n319_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT56), .ZN(new_n833_));
  AOI211_X1 g632(.A(new_n833_), .B(new_n320_), .C1(new_n826_), .C2(new_n827_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n832_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT114), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n831_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n621_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n617_), .A2(new_n619_), .A3(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n621_), .B1(new_n618_), .B2(new_n623_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  MUX2_X1   g640(.A(new_n841_), .B(new_n625_), .S(new_n628_), .Z(new_n842_));
  NAND3_X1  g641(.A1(new_n327_), .A2(new_n324_), .A3(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n324_), .A2(new_n327_), .A3(KEYINPUT115), .A4(new_n842_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n647_), .B1(new_n837_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  XOR2_X1   g649(.A(KEYINPUT116), .B(KEYINPUT58), .Z(new_n851_));
  NAND2_X1  g650(.A1(new_n842_), .A2(new_n321_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n835_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n852_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n854_), .B(KEYINPUT58), .C1(new_n832_), .C2(new_n834_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT117), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n828_), .A2(new_n319_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n833_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n828_), .A2(KEYINPUT56), .A3(new_n319_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n860_), .A2(new_n861_), .A3(KEYINPUT58), .A4(new_n854_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n702_), .A2(new_n853_), .A3(new_n856_), .A4(new_n862_), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n832_), .A2(new_n834_), .A3(KEYINPUT114), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n845_), .B(new_n846_), .C1(new_n864_), .C2(new_n831_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n865_), .A2(KEYINPUT57), .A3(new_n647_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n850_), .A2(new_n863_), .A3(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n823_), .B1(new_n696_), .B2(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n659_), .A2(new_n547_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n425_), .A2(new_n584_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(KEYINPUT59), .B1(new_n868_), .B2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n862_), .A2(new_n856_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n852_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n851_), .ZN(new_n876_));
  OAI22_X1  g675(.A1(new_n875_), .A2(new_n876_), .B1(new_n262_), .B2(new_n265_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n874_), .A2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(KEYINPUT57), .B1(new_n865_), .B2(new_n647_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n873_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n850_), .A2(KEYINPUT118), .A3(new_n863_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n880_), .A2(new_n881_), .A3(new_n866_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n823_), .B1(new_n882_), .B2(new_n696_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n871_), .A2(KEYINPUT59), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n872_), .B1(new_n883_), .B2(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(G113gat), .B1(new_n886_), .B2(new_n634_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n868_), .A2(new_n871_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  OR2_X1    g688(.A1(new_n634_), .A2(G113gat), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n887_), .B1(new_n889_), .B2(new_n890_), .ZN(G1340gat));
  OAI21_X1  g690(.A(G120gat), .B1(new_n886_), .B2(new_n755_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT60), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(G120gat), .ZN(new_n894_));
  AOI21_X1  g693(.A(G120gat), .B1(new_n336_), .B2(new_n893_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(KEYINPUT119), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n896_), .B1(KEYINPUT119), .B2(new_n895_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n888_), .A2(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n892_), .A2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(KEYINPUT120), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n892_), .A2(new_n901_), .A3(new_n898_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n902_), .ZN(G1341gat));
  OAI21_X1  g702(.A(G127gat), .B1(new_n886_), .B2(new_n696_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n888_), .A2(new_n409_), .A3(new_n302_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1342gat));
  AOI21_X1  g705(.A(G134gat), .B1(new_n888_), .B2(new_n646_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n886_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT121), .B(G134gat), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n266_), .A2(new_n909_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n907_), .B1(new_n908_), .B2(new_n910_), .ZN(G1343gat));
  NOR2_X1   g710(.A1(new_n868_), .A2(new_n424_), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n659_), .A2(new_n606_), .A3(new_n584_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n914_), .A2(new_n634_), .ZN(new_n915_));
  XOR2_X1   g714(.A(KEYINPUT122), .B(G141gat), .Z(new_n916_));
  XNOR2_X1  g715(.A(new_n915_), .B(new_n916_), .ZN(G1344gat));
  NOR2_X1   g716(.A1(new_n914_), .A2(new_n755_), .ZN(new_n918_));
  XOR2_X1   g717(.A(new_n918_), .B(G148gat), .Z(G1345gat));
  OR3_X1    g718(.A1(new_n914_), .A2(KEYINPUT123), .A3(new_n696_), .ZN(new_n920_));
  OAI21_X1  g719(.A(KEYINPUT123), .B1(new_n914_), .B2(new_n696_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(KEYINPUT61), .B(G155gat), .ZN(new_n922_));
  AND3_X1   g721(.A1(new_n920_), .A2(new_n921_), .A3(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n922_), .B1(new_n920_), .B2(new_n921_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1346gat));
  OAI21_X1  g724(.A(G162gat), .B1(new_n914_), .B2(new_n266_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n646_), .A2(new_n494_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n914_), .B2(new_n927_), .ZN(G1347gat));
  NAND3_X1  g727(.A1(new_n659_), .A2(new_n424_), .A3(new_n584_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n929_), .A2(new_n547_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n882_), .A2(new_n696_), .ZN(new_n932_));
  INV_X1    g731(.A(new_n823_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n931_), .B1(new_n932_), .B2(new_n933_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n338_), .B1(new_n934_), .B2(new_n631_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n936_));
  OAI21_X1  g735(.A(KEYINPUT125), .B1(new_n935_), .B2(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(new_n866_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n850_), .A2(new_n863_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n938_), .B1(new_n939_), .B2(new_n873_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n302_), .B1(new_n940_), .B2(new_n881_), .ZN(new_n941_));
  OAI211_X1 g740(.A(new_n631_), .B(new_n930_), .C1(new_n941_), .C2(new_n823_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n942_), .A2(new_n936_), .A3(G169gat), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n943_), .A2(new_n944_), .ZN(new_n945_));
  NAND4_X1  g744(.A1(new_n942_), .A2(KEYINPUT124), .A3(new_n936_), .A4(G169gat), .ZN(new_n946_));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n947_));
  NOR3_X1   g746(.A1(new_n883_), .A2(new_n634_), .A3(new_n931_), .ZN(new_n948_));
  OAI211_X1 g747(.A(new_n947_), .B(KEYINPUT62), .C1(new_n948_), .C2(new_n338_), .ZN(new_n949_));
  NAND4_X1  g748(.A1(new_n937_), .A2(new_n945_), .A3(new_n946_), .A4(new_n949_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n948_), .A2(new_n339_), .A3(new_n341_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n950_), .A2(new_n951_), .ZN(G1348gat));
  AOI21_X1  g751(.A(G176gat), .B1(new_n934_), .B2(new_n336_), .ZN(new_n953_));
  INV_X1    g752(.A(new_n868_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n954_), .A2(new_n606_), .ZN(new_n955_));
  INV_X1    g754(.A(new_n955_), .ZN(new_n956_));
  NOR3_X1   g755(.A1(new_n755_), .A2(new_n929_), .A3(new_n342_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n953_), .B1(new_n956_), .B2(new_n957_), .ZN(G1349gat));
  OAI21_X1  g757(.A(new_n930_), .B1(new_n941_), .B2(new_n823_), .ZN(new_n959_));
  NOR3_X1   g758(.A1(new_n959_), .A2(new_n386_), .A3(new_n696_), .ZN(new_n960_));
  OR3_X1    g759(.A1(new_n955_), .A2(new_n696_), .A3(new_n929_), .ZN(new_n961_));
  AOI21_X1  g760(.A(new_n960_), .B1(new_n356_), .B2(new_n961_), .ZN(G1350gat));
  NOR2_X1   g761(.A1(new_n959_), .A2(new_n266_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n963_), .A2(new_n357_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n646_), .A2(new_n387_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n959_), .A2(new_n965_), .ZN(new_n966_));
  OAI21_X1  g765(.A(KEYINPUT126), .B1(new_n964_), .B2(new_n966_), .ZN(new_n967_));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n968_));
  OAI221_X1 g767(.A(new_n968_), .B1(new_n959_), .B2(new_n965_), .C1(new_n963_), .C2(new_n357_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n967_), .A2(new_n969_), .ZN(G1351gat));
  NOR3_X1   g769(.A1(new_n609_), .A2(new_n606_), .A3(new_n583_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n912_), .A2(new_n971_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n972_), .A2(KEYINPUT127), .ZN(new_n973_));
  INV_X1    g772(.A(KEYINPUT127), .ZN(new_n974_));
  NAND3_X1  g773(.A1(new_n912_), .A2(new_n974_), .A3(new_n971_), .ZN(new_n975_));
  AOI21_X1  g774(.A(new_n634_), .B1(new_n973_), .B2(new_n975_), .ZN(new_n976_));
  XNOR2_X1  g775(.A(new_n976_), .B(new_n430_), .ZN(G1352gat));
  AOI21_X1  g776(.A(new_n755_), .B1(new_n973_), .B2(new_n975_), .ZN(new_n978_));
  XNOR2_X1  g777(.A(new_n978_), .B(new_n428_), .ZN(G1353gat));
  XNOR2_X1  g778(.A(KEYINPUT63), .B(G211gat), .ZN(new_n980_));
  AOI211_X1 g779(.A(new_n696_), .B(new_n980_), .C1(new_n973_), .C2(new_n975_), .ZN(new_n981_));
  NAND2_X1  g780(.A1(new_n973_), .A2(new_n975_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n982_), .A2(new_n302_), .ZN(new_n983_));
  NOR2_X1   g782(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n984_));
  AOI21_X1  g783(.A(new_n981_), .B1(new_n983_), .B2(new_n984_), .ZN(G1354gat));
  INV_X1    g784(.A(G218gat), .ZN(new_n986_));
  NAND3_X1  g785(.A1(new_n982_), .A2(new_n986_), .A3(new_n646_), .ZN(new_n987_));
  AOI21_X1  g786(.A(new_n266_), .B1(new_n973_), .B2(new_n975_), .ZN(new_n988_));
  OAI21_X1  g787(.A(new_n987_), .B1(new_n988_), .B2(new_n986_), .ZN(G1355gat));
endmodule


